* NGSPICE file created from Feedback_Divider_mag_flat.ext - technology: gf180mcuC

.subckt pex_Feedback_Divider_mag VSS VDD RST Vdiv F2 F1 F0 CLK
X0 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t2 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD90.t403 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1 Vdiv mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 VDD.t149 VDD.t148 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2 VDD96 RST.t2 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD96.t294 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X3 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 VDD93.t65 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X4 CLK_div_90_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_90_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS.t237 VSS.t236 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X5 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 a_50263_5143# VSS.t2016 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X6 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 a_39120_n10028# VSS.t1944 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X7 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t2 VSS.t2419 VSS.t2418 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X8 CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.t3 VSS.t2422 VSS.t721 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X9 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 VDD90.t367 VDD90.t366 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X10 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD99.t381 VDD99.t380 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X11 a_49276_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VSS.t1635 VSS.t1634 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X12 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t3 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD93.t449 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X13 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 VDD100.t289 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X14 dec3x8_ibr_mag_0.and_3_ibr_5.nand3_mag_ibr_0.OUT F0.t0 VDD.t62 VDD.t61 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X15 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_53892_n2243# VSS.t230 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X16 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t3 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VSS.t1258 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X17 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 VDD93.t128 VDD93.t127 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X18 VSS VDD90.t471 a_30502_11196# VSS.t225 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X19 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD90.t121 VDD90.t120 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X20 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD110.t4 VDD110.t3 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X21 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VDD99.t36 VDD99.t35 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X22 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_100_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 VDD100.t390 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X23 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 VSS.t2229 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X24 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT VDD99.t184 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X25 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD99.t112 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X26 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t3 a_33204_6159# VSS.t1164 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X27 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 a_27381_n699# VSS.t2550 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X28 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 VDD100.t462 VDD100.t461 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X29 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 a_46081_5187# VSS.t2120 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X30 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT VDD100.t35 VDD100.t34 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X31 VDD108 VDD108.t40 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VDD108.t41 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X32 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VDD105.t34 VDD105.t33 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X33 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_28495_6115# VSS.t239 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X34 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t1 VDD110.t420 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X35 a_44075_6240# VDD105.t476 VSS.t1088 VSS.t1087 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X36 VSS CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_31451_n17626# VSS.t1515 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X37 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN VSS.t1519 VSS.t1518 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X38 a_45006_10154# RST.t3 a_44846_10154# VSS.t2082 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X39 a_54751_n16684# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT VSS.t2311 VSS.t2310 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X40 CLK_div_108_new_mag_0.JK_FF_mag_1.QB CLK_div_108_new_mag_0.JK_FF_mag_1.Q a_51957_n6821# VSS.t2317 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X41 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_51239_n5724# VSS.t2320 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X42 a_27144_10099# CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t2 a_26984_10099# VSS.t1178 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X43 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.t3 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD90.t235 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X44 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD90.t414 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X45 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 a_25472_5018# VSS.t2263 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X46 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN VDD110.t117 VDD110.t116 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X47 a_21277_n6009# CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t4 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB VSS.t2385 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X48 a_52225_n13362# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 VDD110.t63 VDD110.t62 pfet_03v3 ad=0.624p pd=2.92u as=1.06p ps=5.68u w=2.4u l=0.28u
X49 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD90.t128 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X50 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t3 VDD100.t248 VDD100.t247 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X51 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD110.t67 VDD110.t66 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X52 a_44779_n16724# RST.t4 a_44619_n16724# VSS.t2081 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X53 VSS CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_32071_11196# VSS.t484 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X54 a_29801_1733# CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 VDD96.t257 VDD96.t256 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X55 a_45251_n1102# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t1800 VSS.t1799 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X56 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_55315_n16684# VSS.t1806 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X57 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB VDD93.t64 VDD93.t63 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X58 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t3 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VDD90.t252 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X59 a_53780_n10161# CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT VSS.t656 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X60 a_24116_n1789# CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t662 VSS.t661 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X61 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_46246_n10116# VSS.t663 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X62 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD90.t134 VDD90.t133 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X63 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD110.t382 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X64 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.CLK CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VDD100.t313 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X65 a_31346_5018# VDD90.t472 VSS.t224 VSS.t223 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X66 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT VDD108.t132 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X67 a_23123_n7106# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VSS.t268 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X68 a_22405_n6009# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VSS.t905 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X69 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_54568_5187# VSS.t910 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X70 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VSS.t865 VSS.t864 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X71 a_50441_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_50281_n17599# VSS.t875 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X72 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 VDD100.t165 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X73 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD93.t259 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X74 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD108.t190 VDD108.t189 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X75 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 VDD90.t365 VDD90.t364 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X76 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 a_50903_n5# VSS.t1039 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X77 CLK_div_96_mag_0.JK_FF_mag_2.Q CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD96.t315 VDD96.t314 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X78 a_45541_n18696# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t2163 VSS.t2162 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X79 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t3 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT VDD93.t452 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X80 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K VDD99.t400 VDD99.t399 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X81 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 VDD93.t422 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X82 a_33180_n17626# CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.t3 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB VSS.t852 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X83 a_51165_n17599# RST.t5 a_51005_n17599# VSS.t2080 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X84 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 VDD99.t440 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X85 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK VSS.t703 VSS.t702 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X86 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB VDD100.t164 VDD100.t163 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X87 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD93.t227 VDD93.t226 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X88 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD93.t231 VDD93.t230 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X89 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD90.t286 VDD90.t285 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X90 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_46105_n18696# VSS.t1317 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X91 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_29680_398# VSS.t1330 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X92 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K VDD90.t468 VDD90.t467 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X93 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT Vdiv96.t2 a_36873_n1222# VSS.t537 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X94 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT VDD99.t402 VDD99.t401 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X95 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 a_43719_n120# VDD100.t108 pfet_03v3 ad=1.06p pd=5.68u as=0.624p ps=2.92u w=2.4u l=0.28u
X96 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD99.t225 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X97 a_27227_398# CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t1401 VSS.t1400 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X98 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 a_29087_8532# VDD90.t311 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X99 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB VDD99.t230 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X100 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD110.t130 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X101 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_44625_n15583# VSS.t837 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X102 a_48380_6284# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VSS.t840 VSS.t839 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X103 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t2 a_51646_1671# VSS.t532 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X104 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VDD100.t126 VDD100.t125 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X105 CLK_div_96_mag_0.JK_FF_mag_3.QB CLK_div_96_mag_0.JK_FF_mag_3.Q a_30589_n2952# VSS.t446 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X106 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 VSS.t455 VSS.t454 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X107 CLK_div_100_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_100_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VDD100.t122 VDD100.t121 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_44475_n5176# VSS.t463 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X109 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT VDD99.t187 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X110 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB VDD100.t432 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X111 a_44799_n7920# CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.t3 CLK_div_108_new_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN VSS.t502 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X112 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_44282_10154# VSS.t2329 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X113 VDD96 CLK_div_96_mag_0.JK_FF_mag_2.Q CLK_div_96_mag_0.JK_FF_mag_2.QB VDD96.t326 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X114 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 VDD99.t432 VDD99.t431 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X115 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_45815_n1102# VSS.t2248 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X116 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t2 VDD108.t89 VDD108.t88 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X117 a_26426_11196# RST.t6 a_26266_11196# VSS.t2079 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X118 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD90.t410 VDD90.t409 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X119 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN VDD110.t442 VDD110.t441 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X120 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB VDD100.t458 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X121 VDD93 VDD93.t106 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD93.t107 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X122 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_26196_5018# VSS.t1418 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X123 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t3 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT VDD105.t89 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X124 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 VDD105.t268 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X125 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT VSS.t919 VSS.t918 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X126 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VDD108.t163 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X127 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 a_50358_1671# VSS.t929 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X128 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD99.t92 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X129 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT a_50923_n10161# VSS.t939 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X130 dec3x8_ibr_mag_0.and_3_ibr_1.nand3_mag_ibr_0.OUT dec3x8_ibr_mag_0.and_3_ibr_3.IN1 VDD.t14 VDD.t13 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X131 a_27375_n17626# CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t282 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X132 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 VDD93.t119 VDD93.t118 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X133 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 a_51871_n5# VSS.t886 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X134 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD93.t124 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X135 VDD100 VDD100.t102 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT VDD100.t103 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X136 VDD99 VDD99.t52 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD99.t53 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X137 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t5 VDD93.t301 VDD93.t300 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X138 a_50263_5143# CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 a_50103_5143# VSS.t688 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X139 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K VDD110.t113 VDD110.t112 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X140 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN VSS.t693 VSS.t692 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X141 a_37237_n8887# CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t1046 VSS.t1045 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X142 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_108_new_mag_0.JK_FF_mag_0.QB a_53255_n5765# VSS.t1048 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X143 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD96.t105 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X144 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_53973_n6862# VSS.t1057 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X145 VDD100 dec3x8_ibr_mag_0.and_3_ibr_2.nand3_mag_ibr_0.OUT VSS.t1061 VSS.t648 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X146 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_48148_n17599# VSS.t1999 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X147 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD100.t147 VDD100.t146 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X148 a_40818_n8887# CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t634 VSS.t633 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X149 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VDD105.t129 VDD105.t128 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X150 VDD96 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD96.t73 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X151 a_47994_n18696# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VSS.t642 VSS.t641 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X152 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT VDD108.t123 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X153 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 a_46623_2768# VSS.t2323 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X154 VDD mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I1 VDD.t150 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X155 a_50922_1671# CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 VSS.t2185 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X156 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_49042_n16682# VSS.t2190 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X157 a_54866_n1102# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t2194 VSS.t2193 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X158 a_32009_n18723# CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t2 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VSS.t2304 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X159 a_43831_7266# CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT a_43671_7266# VDD105.t440 pfet_03v3 ad=0.624p pd=2.92u as=0.624p ps=2.92u w=2.4u l=0.28u
X160 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_48944_6284# VSS.t1131 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X161 a_25646_n17626# CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.t3 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS.t2374 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X162 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 a_30915_n13291# VSS.t1134 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X163 a_27381_n699# CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t1054 VSS.t1053 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X164 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 VDD105.t226 VDD105.t225 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X165 a_46081_5187# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t1143 VSS.t1142 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X166 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t4 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VDD100.t254 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X167 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT RST.t7 VDD99.t377 VDD99.t376 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X168 VSS VDD90.t473 a_24133_11196# VSS.t220 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X169 a_28495_6115# CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 a_28335_6115# VSS.t2262 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X170 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 VSS.t1972 VSS.t1971 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X171 a_38561_880# mux_8x1_ibr_0.mux_2x1_ibr_0.I1 VSS.t1976 VSS.t1975 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X172 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 a_25482_n16632# VSS.t1982 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X173 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN VDD93.t380 VDD93.t379 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X174 a_51641_n9064# CLK.t0 a_51481_n9064# VSS.t2467 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X175 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_53469_n15631# VSS.t1808 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X176 a_27180_n15491# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t1991 VSS.t1990 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X177 VDD90 VDD90.t79 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VDD90.t80 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X178 a_25472_5018# CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 a_25312_5018# VSS.t1633 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X179 VSS VDD100.t477 a_48635_2768# VSS.t2388 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X180 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 VDD96.t369 VDD96.t368 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X181 VSS CLK.t1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VSS.t2468 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X182 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD90.t470 VDD90.t469 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X183 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 VDD110.t179 VDD110.t178 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X184 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 VSS.t972 VSS.t971 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X185 a_43963_n1146# VDD100.t478 VSS.t2392 VSS.t2391 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X186 a_44681_n2243# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS.t1887 VSS.t1886 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X187 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_51729_n17599# VSS.t832 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X188 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK.t2 VDD99.t489 VDD99.t488 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X189 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 VDD110.t348 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X190 Vdiv100 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT VSS.t1896 VSS.t1895 nfet_03v3 ad=86.8f pd=0.92u as=86.8f ps=0.92u w=0.22u l=0.28u
X191 a_50917_n9020# CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t1900 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X192 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t3 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 VSS.t1221 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X193 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 VDD100.t338 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X194 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.t2 VDD108.t326 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X195 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_43757_n6273# VSS.t493 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X196 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 a_28617_n16634# VSS.t2354 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X197 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT VDD99.t417 VDD99.t416 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X198 a_51983_7381# CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 VSS.t2015 VSS.t2014 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X199 VDD96 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD96.t301 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X200 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t3 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VDD105.t441 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X201 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VDD100.t366 VDD100.t365 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X202 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t3 a_30244_398# VSS.t2201 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X203 VDD96 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD96.t238 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X204 a_24901_n6010# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VSS.t1701 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X205 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT a_51040_10154# VSS.t1702 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X206 a_25619_n7107# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VSS.t295 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X207 a_54509_2768# CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t5 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VSS.t1261 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X208 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB VDD110.t440 VDD110.t439 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X209 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t2 VDD93.t355 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X210 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN VDD99.t410 VDD99.t409 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X211 a_54568_5187# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS.t1718 VSS.t1717 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X212 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK VDD110.t77 VDD110.t76 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X213 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 VDD100.t135 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X214 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD93.t229 VDD93.t228 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X215 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN VDD110.t93 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X216 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_37801_n8887# VSS.t561 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X217 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN VDD93.t175 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X218 a_46735_10154# CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t4 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB VSS.t487 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X219 VDD110 CLK.t3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT VDD110.t460 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X220 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VDD108.t176 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X221 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD93.t44 VDD93.t43 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X222 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_44885_n6273# VSS.t146 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X223 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB VDD110.t201 VDD110.t200 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X224 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 a_22551_n16006# VSS.t1981 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X225 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD108.t56 VDD108.t55 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X226 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VDD100.t40 VDD100.t39 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X227 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD93.t50 VDD93.t49 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X228 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t3 VDD100.t223 VDD100.t222 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X229 a_40254_n8887# CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t159 VSS.t158 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X230 a_53458_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_53298_n17599# VSS.t1328 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X231 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD100.t45 VDD100.t44 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X232 dec3x8_ibr_mag_0.and_3_ibr_5.nand3_mag_ibr_0.OUT F0.t1 a_37328_6265# VSS.t278 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X233 a_54302_n1102# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t229 VSS.t228 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X234 VSS VDD108.t455 a_51647_n10161# VSS.t508 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X235 a_29087_8532# CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.t3 CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN VDD90.t219 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X236 a_53221_2768# CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t2006 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X237 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD96.t14 VDD96.t13 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X238 a_48558_n18696# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VSS.t1998 VSS.t1997 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X239 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t6 VDD100.t258 VDD100.t257 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X240 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 VDD110.t435 VDD110.t434 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X241 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.t0 VDD99.t253 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X242 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD93.t365 VDD93.t364 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X243 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 VDD99.t332 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X244 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD110.t115 VDD110.t114 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X245 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_54592_n18696# VSS.t109 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X246 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_108_new_mag_0.JK_FF_mag_1.Q a_50105_n6865# VSS.t2316 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X247 a_45081_n10160# CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.t3 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VSS.t2219 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X248 a_44436_9057# CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t331 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X249 a_51592_n16680# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT VSS.t1725 VSS.t1724 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X250 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VSS.t1727 VSS.t1726 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X251 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD90.t395 VDD90.t394 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X252 a_55067_297# CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT a_54907_297# VDD100.t292 pfet_03v3 ad=0.624p pd=2.92u as=0.624p ps=2.92u w=2.4u l=0.28u
X253 a_26206_n16632# RST.t8 a_26046_n16632# VSS.t2078 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X254 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN VDD110.t293 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X255 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VDD90.t155 VDD90.t154 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X256 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t5 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN VDD105.t92 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X257 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 a_55132_5187# VSS.t911 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X258 a_50353_n9020# CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t1952 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X259 a_43383_n9019# CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t3 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.t0 VSS.t991 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X260 CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.t4 VSS.t2376 VSS.t2375 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X261 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VDD105.t373 VDD105.t372 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X262 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_40408_n9984# VSS.t705 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X263 a_50358_1671# CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 VSS.t1964 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X264 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_23142_n2930# VSS.t1970 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X265 a_53463_n16728# CLK.t4 a_53303_n16728# VSS.t2471 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X266 a_23967_10099# CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t3 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS.t1178 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X267 a_44799_6284# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS.t1743 VSS.t1742 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X268 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t2 VDD99.t481 VDD99.t480 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X269 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VDD108.t306 VDD108.t305 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X270 a_37999_n1822# mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 VSS.t1750 VSS.t795 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X271 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 VDD100.t217 VDD100.t216 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X272 a_46974_n2243# VDD100.t479 VSS.t2394 VSS.t2393 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X273 VDD96 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_2.OUT CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT VDD96.t248 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X274 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I1 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 VDD.t140 VDD.t139 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X275 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD110.t309 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X276 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT VDD110.t379 VDD110.t378 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X277 VSS CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_29772_10099# VSS.t1788 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X278 VSS VDD105.t477 a_54781_10154# VSS.t1089 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X279 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I1 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 VDD.t144 VDD.t143 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X280 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 a_37955_n9984# VSS.t287 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X281 VSS CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_30881_n18723# VSS.t1793 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X282 a_27850_n9876# VDD93.t474 VSS.t274 VSS.t273 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X283 dec3x8_ibr_mag_0.and_3_ibr_1.nand3_mag_ibr_0.OUT dec3x8_ibr_mag_0.and_3_ibr_3.IN1 a_37328_6821# VSS.t278 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X284 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD99.t302 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X285 a_43671_7266# CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 Vdiv105.t2 VDD105.t348 pfet_03v3 ad=0.624p pd=2.92u as=1.06p ps=5.68u w=2.4u l=0.28u
X286 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_44977_n18696# VSS.t1827 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X287 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_53333_10154# VSS.t636 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X288 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t6 a_46867_7960# VSS.t488 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X289 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT VDD110.t99 VDD110.t98 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X290 a_28546_n743# CLK_div_96_mag_0.JK_FF_mag_3.Q a_28386_n743# VSS.t445 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X291 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT RST.t9 VDD105.t406 VDD105.t405 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X292 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_2.Q VSS.t2160 VSS.t2159 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X293 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t1 VDD100.t314 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X294 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_26052_n15491# VSS.t1855 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X295 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB VDD99.t327 VDD99.t326 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X296 VSS CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_2.OUT a_23145_810# VSS.t1753 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X297 a_22718_8532# CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.t4 CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VDD90.t439 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X298 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t3 VDD100.t128 VDD100.t127 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X299 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 VDD105.t359 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X300 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 a_48986_n2199# VSS.t885 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X301 VDD90 VDD90.t75 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD90.t76 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X302 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT a_50922_1671# VSS.t1916 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X303 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD100.t329 VDD100.t328 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X304 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT RST.t10 VDD99.t375 VDD99.t374 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X305 a_26790_n9831# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t807 VSS.t806 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X306 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t3 a_55156_n18696# VSS.t109 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X307 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN VDD93.t253 VDD93.t252 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X308 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_45363_6284# VSS.t813 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X309 a_52156_n16680# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 VSS.t1784 VSS.t1783 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X310 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 VSS.t1805 VSS.t913 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X311 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VDD110.t381 VDD110.t380 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X312 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 VDD105.t347 VDD105.t346 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X313 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT RST.t11 VDD100.t386 VDD100.t385 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X314 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VDD105.t177 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X315 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD108.t82 VDD108.t81 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X316 VSS CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_31661_10099# VSS.t818 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X317 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD105.t1 VDD105.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X318 a_26932_n2952# CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VSS.t2142 VSS.t1697 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X319 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_53487_9057# VSS.t1426 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X320 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t4 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT VDD99.t150 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X321 a_53819_n5721# CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS.t1050 VSS.t1049 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X322 a_22011_n287# CLK_div_96_mag_0.JK_FF_mag_5.QB CLK_div_96_mag_0.JK_FF_mag_5.Q.t0 VSS.t65 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X323 VDD105 RST.t12 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VDD105.t402 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X324 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VDD100.t14 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X325 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 a_30760_n20290# VDD99.t8 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X326 a_23403_10099# CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t112 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X327 CLK_div_96_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 a_28828_1497# VSS.t2549 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X328 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN VDD99.t39 VDD99.t38 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X329 VSS CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t4 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VSS.t1236 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X330 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 VDD105.t434 VDD105.t433 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X331 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t5 VDD99.t154 VDD99.t153 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X332 a_54051_9057# CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t635 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X333 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 VDD110.t224 VDD110.t223 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X334 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN VDD110.t53 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X335 a_31129_n6271# CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 VSS.t412 VSS.t411 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X336 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t4 VDD105.t445 VDD105.t444 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X337 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD99.t98 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X338 a_45753_n15583# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t482 VSS.t481 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X339 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_47430_n18696# VSS.t895 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X340 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD100.t54 VDD100.t53 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X341 a_47190_n16726# CLK.t5 a_47030_n16726# VSS.t2472 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X342 VSS CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN VSS.t896 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X343 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD110.t317 VDD110.t316 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X344 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t0 VDD110.t50 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X345 a_28267_n7033# CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t3 VSS.t996 VSS.t125 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X346 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_53850_6284# VSS.t1716 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X347 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT VDD100.t319 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X348 VSS VDD96.t370 a_23863_n287# VSS.t1482 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X349 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.t4 VDD108.t368 VDD108.t367 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X350 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 VDD105.t149 VDD105.t148 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X351 a_50928_2768# RST.t13 a_50768_2768# VSS.t2077 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X352 a_50287_n18696# VDD110.t494 VSS.t1008 VSS.t1007 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X353 a_35032_n17626# CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.t4 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VSS.t853 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X354 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t3 a_43993_n13477# VDD110.t454 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X355 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.t3 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD99.t452 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X356 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VDD100.t325 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X357 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t4 a_50310_n15627# VSS.t2361 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X358 VDD96 CLK_div_96_mag_0.JK_FF_mag_5.Q.t3 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD96.t110 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X359 a_48888_n15585# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t2091 VSS.t2090 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X360 a_24778_n9875# VDD93.t475 VSS.t272 VSS.t271 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X361 a_33359_11196# CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.t3 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VSS.t753 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X362 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 Vdiv110.t4 VDD.t39 VDD.t38 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X363 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD93.t414 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X364 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN VSS.t811 VSS.t810 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X365 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VDD105.t466 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X366 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t4 VDD105.t233 VDD105.t232 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X367 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t7 VDD100.t238 VDD100.t237 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X368 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK.t6 VDD100.t469 VDD100.t346 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X369 VDD mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_2x1_ibr_0.I0 VDD.t133 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X370 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD110.t299 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X371 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t3 CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 VDD93.t239 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X372 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t2 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VDD90.t161 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X373 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.t4 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VDD108.t106 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X374 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t8 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN VDD100.t239 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X375 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VDD110.t303 VDD110.t302 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X376 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD105.t338 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X377 VSS CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.IN1 a_22575_n287# VSS.t1870 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X378 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t4 VDD93.t270 VDD93.t269 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X379 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT RST.t14 VDD93.t410 VDD93.t409 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X380 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 a_22455_5018# VSS.t1632 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X381 a_36024_n15495# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 VSS.t2545 VSS.t2544 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X382 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD100.t99 VDD100.t101 VDD100.t100 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X383 VSS CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_25856_10099# VSS.t112 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X384 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD96.t133 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X385 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t2 VDD100.t332 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X386 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_26099_398# VSS.t178 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X387 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD99.t329 VDD99.t328 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X388 a_22620_n9884# RST.t15 a_22460_n9884# VSS.t2076 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X389 a_21902_n8787# CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t6 a_21742_n8787# VSS.t1162 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X390 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD110.t266 VDD110.t265 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X391 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB VDD108.t364 VDD108.t363 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X392 a_31352_6115# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K VSS.t2540 VSS.t2539 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X393 a_25800_n18723# CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t2 a_25640_n18723# VSS.t1117 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X394 a_55020_n2199# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t627 VSS.t626 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X395 a_36667_n10028# CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS.t289 VSS.t288 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X396 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t9 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 VDD100.t242 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X397 a_46867_7960# CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t5 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN VSS.t488 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X398 a_51652_2768# CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t10 a_51492_2768# VSS.t1151 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X399 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB VDD105.t122 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X400 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VDD99.t403 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X401 VDD93 CLK.t7 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VDD93.t461 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X402 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_51551_5187# VSS.t1840 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X403 a_28386_n743# VDD96.t371 VSS.t1481 VSS.t1480 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X404 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 VDD100.t412 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X405 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 VDD110.t363 VDD110.t362 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X406 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN VSS.t584 VSS.t583 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X407 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD99.t60 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X408 VSS CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_28490_11196# VSS.t587 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X409 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.t4 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VDD90.t220 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X410 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_96_mag_0.JK_FF_mag_3.QB VDD96.t80 VDD96.t79 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X411 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD96.t203 VDD96.t202 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X412 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 a_45603_n5176# VSS.t1618 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X413 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t6 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT VDD99.t155 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X414 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT RST.t16 VDD108.t357 VDD108.t356 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X415 a_23289_n6009# CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t5 a_23129_n6009# VSS.t997 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X416 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.t0 VDD90.t189 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X417 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD108.t50 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X418 VSS VDD99.t510 a_32175_n17626# VSS.t2423 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X419 a_45570_10154# CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VSS.t1824 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X420 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB VDD100.t411 VDD100.t410 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X421 a_55357_n20487# CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT a_55197_n20487# VDD110.t264 pfet_03v3 ad=0.624p pd=2.92u as=0.624p ps=2.92u w=2.4u l=0.28u
X422 a_24944_n8778# CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 a_24784_n8778# VSS.t453 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X423 a_44247_n17599# VDD110.t495 VSS.t1010 VSS.t1009 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X424 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t3 VDD99.t172 VDD99.t171 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X425 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD90.t326 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X426 VDD105 VDD105.t73 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VDD105.t74 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X427 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD105.t70 VDD105.t72 VDD105.t71 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X428 VSS CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT VSS.t717 nfet_03v3 ad=86.8f pd=0.92u as=86.8f ps=0.92u w=0.22u l=0.28u
X429 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t2 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT VDD105.t210 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X430 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t6 VDD93.t272 VDD93.t271 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X431 a_45363_6284# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t1456 VSS.t1455 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X432 a_22264_n1833# VDD96.t372 VSS.t1479 VSS.t1478 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X433 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t6 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN VDD105.t234 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X434 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD105.t174 VDD105.t173 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X435 a_54504_n10161# CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.t3 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT VSS.t1187 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X436 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT VDD100.t189 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X437 a_47332_n5176# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS.t1660 VSS.t1659 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X438 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t0 VDD93.t374 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X439 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD93.t223 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X440 Vdiv108 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD108.t304 VDD108.t303 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X441 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD93.t342 VDD93.t341 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X442 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS.t1 VSS.t0 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X443 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K VDD99.t390 VDD99.t389 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X444 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD110.t155 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X445 a_53487_9057# CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t1960 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X446 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_1.IN2 VDD.t120 VDD.t119 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X447 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 a_23510_n15620# VDD99.t205 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X448 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.t2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB VDD93.t37 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X449 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD105.t197 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X450 a_28552_354# CLK_div_96_mag_0.JK_FF_mag_3.Q a_28392_354# VSS.t444 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X451 a_45449_n6273# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t147 VSS.t146 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X452 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD110.t426 VDD110.t425 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X453 a_24307_5062# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t2256 VSS.t1624 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X454 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD105.t207 VDD105.t206 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X455 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT VDD93.t426 VDD93.t425 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X456 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD93.t340 VDD93.t339 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X457 VSS CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_25292_10099# VSS.t112 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X458 VDD110 RST.t17 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VDD110.t410 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X459 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 a_34890_n16636# VSS.t1583 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X460 a_29110_n743# CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS.t1585 VSS.t1584 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X461 a_36588_n15495# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 VSS.t1587 VSS.t1586 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X462 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD90.t72 VDD90.t74 VDD90.t73 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X463 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VDD105.t343 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X464 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 VDD105.t312 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X465 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 VDD110.t197 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X466 a_50868_n16724# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT VSS.t1362 VSS.t1361 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X467 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB VDD110.t336 VDD110.t335 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X468 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD93.t233 VDD93.t232 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X469 a_26770_n16588# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT VSS.t1854 VSS.t1853 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X470 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_54597_n15587# VSS.t1364 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X471 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.IN2 a_50232_n7685# VDD108.t246 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X472 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t7 a_47835_7960# VSS.t488 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X473 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD99.t211 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X474 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD93.t370 VDD93.t369 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X475 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD93.t316 VDD93.t315 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X476 a_23863_n287# CLK_div_96_mag_0.JK_FF_mag_4.Q.t3 a_23703_n287# VSS.t2282 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X477 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 a_35614_n16636# VSS.t2543 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X478 a_29751_n15493# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t2140 VSS.t2139 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X479 a_22121_11196# CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.t5 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K VSS.t2386 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X480 a_50768_2768# CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT VSS.t928 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X481 VSS CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN VSS.t75 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X482 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.JK_FF_mag_3.QB a_30435_n1855# VSS.t448 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X483 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT VDD105.t261 VDD105.t260 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X484 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT VDD100.t295 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X485 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_51393_n6821# VSS.t1390 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X486 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_50675_n5724# VSS.t1392 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X487 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.t4 VDD90.t170 VDD90.t169 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X488 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_47760_n15585# VSS.t1673 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X489 a_21431_n7106# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t1 VSS.t720 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X490 a_46755_574# CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t3 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN VSS.t1082 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X491 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK.t8 VDD99.t491 VDD99.t490 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X492 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K VDD110.t281 VDD110.t280 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X493 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT VDD108.t298 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X494 VDD96 VDD96.t182 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_2.OUT VDD96.t183 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X495 VSS CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_1.IN2 a_22011_n287# VSS.t1686 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X496 VDD96 CLK_div_96_mag_0.JK_FF_mag_0.Q CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VDD96.t230 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X497 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VDD108.t260 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X498 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT CLK.t9 VDD108.t438 VDD108.t437 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X499 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_48268_n1102# VSS.t2466 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X500 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT VDD110.t250 VDD110.t249 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X501 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VDD105.t32 VDD105.t31 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X502 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t4 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT VDD100.t415 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X503 a_29871_n1855# CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VSS.t1612 VSS.t1611 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X504 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t4 a_30164_n7017# VSS.t314 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X505 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 Vdiv105.t0 VSS.t1499 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X506 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD105.t384 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X507 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_51849_n1102# VSS.t169 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X508 a_23552_n1789# CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t1969 VSS.t1968 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X509 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD100.t336 VDD100.t335 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X510 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.t3 VDD108.t408 VDD108.t407 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X511 VSS CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN VSS.t1079 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X512 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD99.t248 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X513 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD93.t331 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X514 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_54051_9057# VSS.t1861 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X515 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VDD90.t337 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X516 a_22575_n287# CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_1.IN2 VSS.t1535 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X517 a_39124_280# mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 VSS.t1537 VSS.t1536 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X518 CLK_div_100_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT VDD100.t162 VDD100.t161 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X519 a_47863_10154# CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT VSS.t1541 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X520 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD105.t86 VDD105.t85 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X521 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT a_50928_2768# VSS.t1760 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X522 a_50874_n15583# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT VSS.t2087 VSS.t2086 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X523 a_54615_9057# CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VSS.t817 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X524 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD110.t388 VDD110.t387 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X525 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t3 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD99.t482 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X526 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VDD110.t107 VDD110.t106 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X527 VSS VDD96.t374 a_23869_810# VSS.t1475 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X528 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 VDD100.t353 VDD100.t352 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X529 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS.t1605 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X530 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_54414_6284# VSS.t909 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X531 a_51492_2768# CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t5 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT VSS.t2273 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X532 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 VDD110.t154 VDD110.t153 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X533 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t5 VDD105.t447 VDD105.t446 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X534 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t3 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VDD99.t121 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X535 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN VDD99.t428 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X536 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VDD99.t283 VDD99.t282 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X537 VSS CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.t5 a_30496_10099# VSS.t754 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X538 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 F0.t2 a_35184_880# VSS.t1163 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X539 CLK_div_96_mag_0.JK_FF_mag_5.Q CLK_div_96_mag_0.JK_FF_mag_5.QB VDD96.t10 VDD96.t9 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X540 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_23706_n2886# VSS.t1647 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X541 CLK_div_99_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.t5 VDD99.t78 VDD99.t77 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X542 CLK_div_96_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_96_mag_0.JK_FF_mag_3.Q VDD96.t72 VDD96.t71 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X543 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_45189_n15583# VSS.t1547 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X544 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t3 VDD105.t189 VDD105.t188 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X545 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 a_33358_5062# VSS.t1812 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X546 VSS CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 a_25686_1919# VSS.t1551 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X547 a_28577_n2996# VDD96.t375 VSS.t1474 VSS.t1473 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X548 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD96.t197 VDD96.t196 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X549 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD110.t127 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X550 VSS CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_34468_n17626# VSS.t1841 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X551 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.CLK VDD105.t308 VDD105.t307 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X552 VDD108 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD108.t206 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X553 VDD108 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD108.t285 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X554 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 VSS.t687 VSS.t686 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X555 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD99.t311 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X556 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD105.t301 VDD105.t300 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X557 a_50204_2768# CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 VSS.t1963 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X558 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_29623_6159# VSS.t299 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X559 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t6 VDD105.t449 VDD105.t448 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X560 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t7 VDD93.t274 VDD93.t273 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X561 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_44321_n6273# VSS.t146 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X562 a_48252_n9063# CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t2 a_48092_n9063# VSS.t2232 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X563 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t3 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VDD90.t164 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X564 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD105.t14 VDD105.t13 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X565 VDD96 VDD96.t178 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_0.OUT VDD96.t179 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X566 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 a_29341_n16634# VSS.t2138 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X567 a_26183_n7107# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VSS.t1453 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X568 a_25465_n6010# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VSS.t1708 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X569 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_51285_n1102# VSS.t1284 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X570 a_50199_n10117# CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t1951 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X571 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD93.t352 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X572 a_29298_n9832# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT VSS.t1568 VSS.t1567 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X573 a_47528_n9019# CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t927 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X574 a_28580_n8735# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT VSS.t651 VSS.t650 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X575 a_49945_n6865# VDD108.t456 VSS.t512 VSS.t511 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X576 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t2 VDD105.t315 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X577 VSS CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t0 VSS.t1381 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X578 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT VDD110.t283 VDD110.t282 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X579 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I1 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT a_36873_n1822# VSS.t537 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X580 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT VDD108.t139 VDD108.t138 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X581 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VDD108.t75 VDD108.t74 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X582 a_31731_n16632# CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t7 a_31571_n16632# VSS.t1165 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X583 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN VDD93.t201 VDD93.t200 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X584 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 VDD105.t125 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X585 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 a_52115_5187# VSS.t2013 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X586 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_35460_n15495# VSS.t1380 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X587 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD100.t96 VDD100.t98 VDD100.t97 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X588 a_33353_10099# CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VSS.t1670 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X589 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 VDD105.t117 VDD105.t116 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X590 VDD110 CLK.t10 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT VDD110.t463 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X591 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_44123_n1146# VSS.t2247 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X592 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD90.t149 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X593 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 VDD90.t334 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X594 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD110.t220 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X595 VDD96 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_1.IN2 VDD96.t267 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X596 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD90.t157 VDD90.t156 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X597 a_54182_n17599# RST.t18 a_54022_n17599# VSS.t2075 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X598 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD110.t386 VDD110.t385 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X599 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 F0.t3 VDD.t64 VDD.t63 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X600 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 VDD105.t437 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X601 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD105.t121 VDD105.t120 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X602 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_49122_n18696# VSS.t894 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X603 a_28823_n17626# CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t4 a_28663_n17626# VSS.t1118 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X604 VDD110 RST.t19 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT VDD110.t407 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X605 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.t2 a_54658_n9064# VSS.t2264 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X606 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD110.t373 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X607 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD99.t222 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X608 a_28743_n1899# CLK_div_96_mag_0.JK_FF_mag_2.Q a_28583_n1899# VSS.t2158 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X609 a_47858_n2243# RST.t20 a_47698_n2243# VSS.t2074 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X610 a_30209_7256# CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 VSS.t1339 VSS.t1338 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X611 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VDD105.t24 VDD105.t23 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X612 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.t4 VDD90.t239 VDD90.t238 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X613 a_28016_n8779# CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t5 a_27856_n8779# VSS.t2420 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X614 a_25529_n743# CLK_div_96_mag_0.JK_FF_mag_3.Q a_25369_n743# VSS.t443 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X615 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 a_40375_n7552# VDD93.t373 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X616 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 VDD100.t185 VDD100.t184 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X617 a_50151_n2243# CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 a_49991_n2243# VSS.t884 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X618 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_108_new_mag_0.JK_FF_mag_0.QB VDD108.t197 VDD108.t196 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X619 a_25055_n7107# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VSS.t1700 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X620 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD108.t203 VDD108.t202 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X621 VSS CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_29208_10099# VSS.t1435 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X622 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB VDD108.t295 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X623 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN VDD110.t165 VDD110.t164 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X624 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t3 a_51758_9057# VSS.t1068 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X625 a_47970_5143# RST.t21 a_47810_5143# VSS.t2073 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X626 VSS CLK.t11 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 VSS.t2473 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X627 VDD mux_8x1_ibr_0.mux_2x1_ibr_0.I0 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT VDD.t136 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X628 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 a_49752_10154# VSS.t1356 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X629 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT a_53940_n10161# VSS.t1656 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X630 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN VSS.t1043 VSS.t1042 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X631 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 VDD105.t279 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X632 a_36310_n1822# Vdiv99.t2 VSS.t2291 VSS.t2290 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X633 a_53008_n2243# VDD100.t480 VSS.t2396 VSS.t2395 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X634 a_23794_n17626# CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.t5 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K VSS.t2377 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X635 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT VDD110.t230 VDD110.t229 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X636 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_5.Q.t4 VDD96.t114 VDD96.t113 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X637 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_1.IN2 Vdiv93.t2 VDD.t161 VDD.t160 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X638 a_45787_574# CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t4 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN VSS.t1081 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X639 a_46774_n6273# CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t3 a_46614_n6273# VSS.t493 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X640 CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD105.t321 VDD105.t320 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X641 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 F1.t0 VDD.t89 VDD.t88 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X642 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 VDD110.t219 VDD110.t218 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X643 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD110.t339 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X644 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD108.t302 VDD108.t301 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X645 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 a_46777_1671# VSS.t2127 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X646 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 VDD93.t328 VDD93.t327 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X647 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 a_29213_n7028# VSS.t143 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X648 a_41124_n14596# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 VSS.t408 VSS.t407 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X649 a_30050_n13332# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 VSS.t1133 VSS.t1132 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X650 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD108.t266 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X651 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD96.t82 VDD96.t81 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X652 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK VDD108.t314 VDD108.t313 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X653 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT VDD110.t139 VDD110.t138 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X654 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 a_50470_9057# VSS.t1591 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X655 a_35026_n18723# CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VSS.t2347 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X656 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t8 VDD99.t159 VDD99.t158 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X657 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 VSS.t2261 VSS.t2260 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X658 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD99.t235 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X659 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD108.t54 VDD108.t53 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X660 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD105.t430 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X661 a_33358_5062# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t2300 VSS.t2299 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X662 a_47534_n10160# RST.t22 a_47374_n10160# VSS.t2072 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X663 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 VDD93.t434 VDD93.t433 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X664 a_25686_1919# CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 VSS.t336 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X665 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN VSS.t974 VSS.t973 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X666 a_26253_n743# RST.t23 a_26093_n743# VSS.t2071 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X667 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_29187_n15493# VSS.t1282 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X668 a_51034_9057# CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 VSS.t1387 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X669 VSS CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.t5 a_24127_10099# VSS.t1178 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X670 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT VDD110.t273 VDD110.t272 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X671 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 a_47134_n2243# VSS.t883 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X672 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t1 VDD99.t338 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X673 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD90.t108 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X674 VSS CLK.t12 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VSS.t2476 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X675 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS.t349 VSS.t348 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X676 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 VDD93.t388 VDD93.t387 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X677 a_28463_n15537# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t2 VSS.t2367 VSS.t2366 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X678 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_46400_n9019# VSS.t363 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X679 a_50875_n2243# RST.t24 a_50715_n2243# VSS.t2070 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X680 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_54746_n17599# VSS.t1936 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X681 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t4 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 VDD99.t173 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X682 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 a_53370_n9020# VSS.t653 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X683 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_50833_6284# VSS.t307 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X684 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_0.OUT CLK_div_96_mag_0.JK_FF_mag_4.Q.t4 VDD96.t337 VDD96.t336 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X685 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK.t13 VDD99.t493 VDD99.t492 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X686 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t4 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 VDD110.t186 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X687 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.IN2 F0.t4 VDD.t66 VDD.t65 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X688 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 VDD93.t438 VDD93.t437 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X689 a_33334_n18723# CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.t1 VSS.t2346 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X690 dec3x8_ibr_mag_0.and_3_ibr_4.nand3_mag_ibr_0.OUT F0.t5 VDD.t68 VDD.t67 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X691 VSS CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_32225_10099# VSS.t1531 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X692 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 VDD105.t147 VDD105.t146 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X693 VDD96 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_1.IN2 CLK_div_96_mag_0.JK_FF_mag_5.Q.t2 VDD96.t217 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X694 VDD99 RST.t25 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT VDD99.t371 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X695 a_54383_n5721# CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t1056 VSS.t1055 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X696 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 F2.t0 a_38561_880# VSS.t1198 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X697 a_32301_n15491# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT VSS.t1433 VSS.t1432 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X698 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.IN2 F0.t6 VSS.t2440 VSS.t2439 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X699 a_30502_11196# CLK.t14 a_30342_11196# VSS.t2479 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X700 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT VDD99.t268 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X701 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t6 VDD100.t419 VDD100.t418 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X702 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_1.IN2 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 VDD96.t189 VDD96.t188 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X703 a_45039_n5176# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS.t465 VSS.t464 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X704 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_96_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD96.t35 VDD96.t34 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X705 a_24358_n17626# CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t1639 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X706 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD99.t273 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X707 a_45907_n16680# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t2293 VSS.t2292 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X708 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t3 VDD108.t377 VDD108.t376 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X709 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_108_new_mag_0.JK_FF_mag_1.Q VDD108.t425 VDD108.t424 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X710 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB VDD110.t162 VDD110.t161 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X711 a_29778_11196# RST.t26 a_29618_11196# VSS.t2069 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X712 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_45405_n2199# VSS.t1764 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X713 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 VDD110.t332 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X714 a_44846_10154# CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VSS.t324 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X715 a_51239_n5724# CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t1395 VSS.t1394 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X716 VSS CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_0.OUT a_26250_1919# VSS.t325 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X717 a_43591_n5176# VDD108.t457 VSS.t514 VSS.t513 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X718 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.t3 VDD99.t116 VDD99.t115 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X719 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD110.t24 VDD110.t26 VDD110.t25 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X720 VDD96 CLK_div_96_mag_0.JK_FF_mag_0.Q CLK_div_96_mag_0.JK_FF_mag_0.QB VDD96.t227 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X721 VSS CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.t6 a_32169_n18723# VSS.t854 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X722 a_44977_n18696# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS.t149 VSS.t148 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X723 VDD96 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_4.IN2 VDD96.t253 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X724 a_51871_n5# CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 VSS.t1038 VSS.t1037 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X725 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD105.t352 VDD105.t351 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X726 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_0.OUT CLK.t15 VDD96.t354 VDD96.t353 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X727 a_53120_5143# VDD105.t479 VSS.t1093 VSS.t1092 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X728 VSS CLK_div_99_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 VSS.t1650 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X729 a_26814_1919# CLK_div_96_mag_0.JK_FF_mag_4.QB CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_0.OUT VSS.t421 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X730 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 VDD99.t287 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X731 a_50144_n16724# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K VSS.t1412 VSS.t1411 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X732 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t9 VDD99.t161 VDD99.t160 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X733 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD93.t121 VDD93.t120 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X734 Vdiv105 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT VSS.t2199 VSS.t2198 nfet_03v3 ad=86.8f pd=0.92u as=86.8f ps=0.92u w=0.22u l=0.28u
X735 a_48098_n10160# CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.t5 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VSS.t503 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X736 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 VDD96.t350 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X737 a_25369_n743# VDD96.t377 VSS.t1472 VSS.t1471 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X738 a_49640_2768# CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t7 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB VSS.t2274 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X739 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT VDD110.t329 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X740 VDD96 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 CLK_div_96_mag_0.JK_FF_mag_4.Q.t0 VDD96.t29 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X741 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 a_21896_n9884# VSS.t452 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X742 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD90.t42 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X743 a_44061_n15627# CLK.t16 a_43901_n15627# VSS.t2480 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X744 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 a_22711_n14504# VSS.t2353 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X745 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_43793_n10116# VSS.t1512 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X746 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 a_28734_n9876# VSS.t1232 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X747 a_51758_9057# CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t7 a_51598_9057# VSS.t2205 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X748 a_25122_1919# CLK_div_96_mag_0.JK_FF_mag_4.QB CLK_div_96_mag_0.JK_FF_mag_4.Q.t1 VSS.t420 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X749 a_54456_n2199# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS.t233 VSS.t232 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X750 VDD90 RST.t27 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VDD90.t440 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X751 a_25484_n2996# VDD96.t378 VSS.t1470 VSS.t1469 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X752 a_24153_6159# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t388 VSS.t387 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X753 a_53089_n6862# VDD108.t458 VSS.t516 VSS.t515 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X754 VDD108 VDD108.t36 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT VDD108.t37 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X755 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT VDD93.t103 VDD93.t105 VDD93.t104 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X756 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 VDD93.t310 VDD93.t309 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X757 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD90.t48 VDD90.t47 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X758 VSS CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT a_22421_810# VSS.t1757 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X759 VSS CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_26420_10099# VSS.t112 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X760 VDD105 VDD105.t66 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT VDD105.t67 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X761 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 a_49906_9057# VSS.t1594 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X762 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD105.t63 VDD105.t65 VDD105.t64 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X763 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 VDD108.t317 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X764 a_28329_5018# VDD90.t476 VSS.t219 VSS.t218 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X765 VDD96 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD96.t68 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X766 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN VDD110.t196 VDD110.t195 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X767 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD108.t85 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X768 VSS CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_31507_11196# VSS.t1303 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X769 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 a_23748_n9840# VSS.t451 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X770 CLK_div_100_mag_0.CLK_div_10_mag_1.CLK CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 a_55067_297# VDD100.t313 pfet_03v3 ad=1.06p pd=5.68u as=0.624p ps=2.92u w=2.4u l=0.28u
X771 a_44687_n1102# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS.t1874 VSS.t1873 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X772 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t6 a_24938_n9875# VSS.t2421 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X773 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB VDD105.t253 VDD105.t252 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X774 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_32076_6159# VSS.t472 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X775 VSS VDD96.t379 a_26974_1919# VSS.t1466 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X776 a_46777_1671# CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t2 VSS.t2327 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X777 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT VDD99.t218 VDD99.t217 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X778 a_43895_n16724# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K VSS.t1377 VSS.t1376 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X779 a_50470_9057# CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 VSS.t613 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X780 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD99.t95 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X781 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t1 VSS.t732 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X782 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 Vdiv100.t2 VSS.t1910 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X783 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_48056_n5176# VSS.t2249 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X784 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB VDD108.t140 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X785 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t5 CLK_div_99_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD99.t124 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X786 CLK_div_108_new_mag_0.JK_FF_mag_1.Q CLK_div_108_new_mag_0.JK_FF_mag_1.QB a_51803_n5724# VSS.t2319 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X787 a_22559_n7106# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VSS.t720 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X788 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD105.t107 VDD105.t106 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X789 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VDD108.t71 VDD108.t70 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X790 VSS CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_29054_11196# VSS.t1439 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X791 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD90.t303 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X792 VDD99 RST.t28 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT VDD99.t368 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X793 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t2 VDD93.t291 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X794 a_32640_6159# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t475 VSS.t474 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X795 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB VDD96.t349 VDD96.t348 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X796 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD90.t69 VDD90.t71 VDD90.t70 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X797 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD96.t307 VDD96.t306 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X798 CLK_div_96_mag_0.JK_FF_mag_2.QB CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD96.t242 VDD96.t241 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X799 a_53464_n18696# CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_53304_n18696# VSS.t689 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X800 a_32795_11196# RST.t29 a_32635_11196# VSS.t2068 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X801 dec3x8_ibr_mag_0.and_3_ibr_5.IN3 F2.t1 VDD.t72 VDD.t71 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X802 a_26093_n743# CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS.t962 VSS.t961 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X803 a_45815_n1102# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t374 VSS.t373 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X804 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD90.t66 VDD90.t68 VDD90.t67 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X805 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD110.t21 VDD110.t23 VDD110.t22 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X806 VSS VDD100.t481 a_48629_1671# VSS.t2397 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X807 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN VSS.t1136 VSS.t1135 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X808 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD93.t411 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X809 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 VDD93.t419 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X810 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD93.t58 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X811 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK.t17 VDD93.t465 VDD93.t464 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X812 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD90.t115 VDD90.t114 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X813 dec3x8_ibr_mag_0.and_3_ibr_0.nand3_mag_ibr_0.OUT dec3x8_ibr_mag_0.and_3_ibr_3.IN1 VDD.t12 VDD.t11 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X814 a_43993_n13477# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 VDD110.t177 VDD110.t176 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X815 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT RST.t30 VDD108.t355 VDD108.t354 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X816 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD93.t217 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X817 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN VDD93.t255 VDD93.t254 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X818 VDD96 dec3x8_ibr_mag_0.and_3_ibr_1.nand3_mag_ibr_0.OUT VSS.t280 VSS.t279 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X819 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t4 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VDD108.t378 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X820 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VDD99.t147 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X821 a_28093_n18723# CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t893 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X822 a_53255_n5765# CLK_div_108_new_mag_0.JK_FF_mag_1.Q a_53095_n5765# VSS.t2315 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X823 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t10 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT VDD99.t162 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X824 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD90.t31 VDD90.t30 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X825 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT VDD99.t291 VDD99.t290 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X826 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_45695_n17599# VSS.t545 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X827 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.VOUT CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VSS.t578 VSS.t577 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X828 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 a_47341_1671# VSS.t1720 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X829 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 VDD110.t49 VDD110.t48 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X830 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD93.t100 VDD93.t102 VDD93.t101 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X831 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_43718_10154# VSS.t2096 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X832 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT a_51034_9057# VSS.t1449 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X833 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 VDD99.t451 VDD99.t450 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X834 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_0.Q VDD96.t226 VDD96.t225 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X835 a_50669_n6865# CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS.t1939 VSS.t1938 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X836 a_24133_11196# CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t5 a_23973_11196# VSS.t1239 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X837 Vdiv96 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS.t425 VSS.t424 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X838 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_23184_n9840# VSS.t679 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X839 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 VDD108.t269 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X840 a_47905_1671# CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 VSS.t118 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X841 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 a_27334_n16588# VSS.t1980 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X842 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD93.t97 VDD93.t99 VDD93.t98 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X843 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t4 a_53286_6240# VSS.t858 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X844 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK.t18 VDD90.t451 VDD90.t450 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X845 a_31291_n17626# CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VSS.t1792 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X846 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD93.t363 VDD93.t362 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X847 VSS VDD93.t476 a_23283_n7106# VSS.t268 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X848 VSS CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_22565_n6009# VSS.t42 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X849 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN VDD93.t184 VDD93.t183 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X850 VSS CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN VSS.t565 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X851 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VDD90.t3 VDD90.t2 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X852 a_33245_7558# CLK_div_90_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 VDD90.t397 VDD90.t396 pfet_03v3 ad=0.624p pd=2.92u as=1.06p ps=5.68u w=2.4u l=0.28u
X853 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_36109_n8931# VSS.t560 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X854 CLK_div_108_new_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 a_47050_n7372# VSS.t497 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X855 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD105.t381 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X856 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_29905_n16590# VSS.t55 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X857 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VDD90.t7 VDD90.t6 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X858 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t4 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD108.t90 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X859 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.JK_FF_mag_1.Q VSS.t2314 VSS.t2313 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X860 a_26990_11196# CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.t6 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS.t1181 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X861 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VDD96.t234 VDD96.t233 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X862 a_50827_5143# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VSS.t106 VSS.t105 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X863 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 VDD100.t457 VDD100.t456 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X864 VDD108 CLK.t19 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 VDD108.t439 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X865 a_47424_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_47264_n17599# VSS.t1327 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X866 a_22258_n2930# VDD96.t380 VSS.t1465 VSS.t1464 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X867 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD90.t91 VDD90.t90 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X868 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB VDD105.t84 VDD105.t83 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X869 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t7 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD93.t302 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X870 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 a_30341_5062# VSS.t1337 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X871 VDD93 RST.t31 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD93.t406 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X872 a_37801_n8887# CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t2095 VSS.t2094 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X873 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t5 VDD108.t382 VDD108.t381 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X874 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN VDD110.t343 VDD110.t342 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X875 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t3 a_48466_n6273# VSS.t146 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X876 a_53897_10154# CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VSS.t1425 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X877 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t8 VDD105.t451 VDD105.t450 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X878 dec3x8_ibr_mag_0.and_3_ibr_4.nand3_mag_ibr_0.OUT F0.t7 a_36202_6265# VSS.t356 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X879 VDD93 RST.t32 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD93.t403 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X880 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD105.t408 VDD105.t407 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X881 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD96.t175 VDD96.t177 VDD96.t176 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X882 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t5 VSS.t495 VSS.t494 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X883 a_31733_n19822# CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.t7 CLK_div_99_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN VSS.t857 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X884 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_46810_n10116# VSS.t924 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X885 a_26036_5018# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VSS.t714 VSS.t713 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X886 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 a_52839_n5# VSS.t1036 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X887 a_32076_6159# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS.t2542 VSS.t2541 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X888 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN VDD99.t140 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X889 a_51005_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VSS.t1342 VSS.t1341 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X890 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 VSS.t313 VSS.t312 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X891 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_50987_5143# VSS.t625 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X892 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD93.t151 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X893 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_46259_n17599# VSS.t1326 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X894 a_28817_n18723# CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t6 a_28657_n18723# VSS.t1119 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X895 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB VDD90.t36 VDD90.t35 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X896 VSS CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_25138_11196# VSS.t345 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X897 a_50105_n6865# CLK_div_108_new_mag_0.JK_FF_mag_1.CLK a_49945_n6865# VSS.t1749 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X898 VDD F0.t8 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 VDD.t166 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X899 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT VDD99.t386 VDD99.t385 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X900 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 VDD90.t363 VDD90.t362 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X901 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 VDD99.t411 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X902 CLK_div_96_mag_0.JK_FF_mag_4.QB CLK_div_96_mag_0.JK_FF_mag_4.Q.t5 VDD96.t339 VDD96.t338 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X903 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_96_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS.t390 VSS.t389 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X904 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VDD90.t278 VDD90.t277 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X905 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 VDD.t113 VDD.t112 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X906 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.t3 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT VDD108.t399 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X907 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD90.t391 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X908 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT a_48023_10154# VSS.t1422 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X909 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t8 VDD100.t421 VDD100.t420 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X910 a_30025_n2952# CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VSS.t1615 VSS.t1614 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X911 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD90.t218 VDD90.t217 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X912 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 F1.t1 VDD.t91 VDD.t90 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X913 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD108.t84 VDD108.t83 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X914 a_51764_10154# CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t9 a_51604_10154# VSS.t2206 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X915 VSS VDD99.t511 a_35192_n17626# VSS.t2426 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X916 VDD108 Vdiv108.t3 CLK_div_108_new_mag_0.JK_FF_mag_0.QB VDD108.t209 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X917 VDD100 RST.t33 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VDD100.t382 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X918 a_40408_n9984# CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS.t162 VSS.t161 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X919 a_23142_n2930# RST.t34 a_22982_n2930# VSS.t2067 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X920 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 VDD108.t245 VDD108.t244 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X921 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.IN2 VSS.t802 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X922 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN VDD99.t76 VDD99.t75 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X923 VSS CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_26965_n18723# VSS.t729 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X924 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD108.t33 VDD108.t35 VDD108.t34 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X925 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_2.OUT CLK.t20 VDD96.t356 VDD96.t355 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X926 VSS CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS.t1941 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X927 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD100.t181 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X928 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 VSS.t966 VSS.t965 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X929 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 VSS.t2189 VSS.t2188 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X930 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD96.t199 VDD96.t198 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X931 VDD96 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD96.t245 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X932 a_50923_n10161# RST.t35 a_50763_n10161# VSS.t2066 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X933 dec3x8_ibr_mag_0.and_3_ibr_0.nand3_mag_ibr_0.OUT dec3x8_ibr_mag_0.and_3_ibr_3.IN1 a_36202_6821# VSS.t277 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X934 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_100_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 VSS.t2132 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X935 VDD108 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD108.t434 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X936 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_1.IN2 F0.t9 a_35184_n1822# VSS.t2441 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X937 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT VDD110.t453 VDD110.t452 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X938 VDD108 CLK_div_108_new_mag_0.JK_FF_mag_1.Q CLK_div_108_new_mag_0.JK_FF_mag_1.QB VDD108.t421 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X939 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_44841_n2243# VSS.t1798 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X940 a_51438_n15583# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 VSS.t830 VSS.t829 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X941 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_25488_n15535# VSS.t970 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X942 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN VDD99.t268 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X943 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 VDD100.t195 VDD100.t194 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X944 a_53333_10154# CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t1959 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X945 VDD F1.t2 dec3x8_ibr_mag_0.and_3_ibr_5.nand3_mag_ibr_0.OUT VDD.t92 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X946 a_32455_n16632# RST.t36 a_32295_n16632# VSS.t2065 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X947 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD100.t93 VDD100.t95 VDD100.t94 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X948 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_50157_n1146# VSS.t168 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X949 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB VDD110.t326 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X950 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD90.t197 VDD90.t196 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X951 a_49042_n16682# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t341 VSS.t340 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X952 a_33204_6159# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t1993 VSS.t1992 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X953 VDD96 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 VDD96.t94 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X954 VDD110 RST.t37 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD110.t404 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X955 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t5 a_52002_n15583# VSS.t2362 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X956 a_53286_6240# CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 a_53126_6240# VSS.t2119 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X957 VSS CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_30163_n17626# VSS.t127 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X958 a_49906_9057# CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t1 VSS.t1309 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X959 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD105.t356 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X960 a_25322_n16632# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K VSS.t184 VSS.t183 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X961 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_48712_n17599# VSS.t397 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X962 a_53309_n15631# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K VSS.t1683 VSS.t1682 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X963 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 VDD110.t158 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X964 a_30915_n13291# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 VSS.t2343 VSS.t2342 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X965 a_24491_n7107# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t0 VSS.t1452 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X966 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t6 VDD90.t256 VDD90.t255 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X967 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD90.t188 VDD90.t187 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X968 VDD93 dec3x8_ibr_mag_0.and_3_ibr_4.nand3_mag_ibr_0.OUT VDD.t6 VDD.t5 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X969 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t11 VSS.t1167 VSS.t1166 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X970 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t7 VDD90.t258 VDD90.t257 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X971 a_39124_880# mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 VSS.t2172 VSS.t1536 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X972 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD105.t16 VDD105.t15 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X973 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 VDD99.t267 VDD99.t266 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X974 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT VDD110.t248 VDD110.t247 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X975 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t0 VDD105.t17 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X976 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 Vdiv105.t1 VSS.t1821 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X977 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 a_43760_1671# VSS.t1905 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X978 a_28457_n16634# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t3 VSS.t2369 VSS.t2368 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X979 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD100.t466 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X980 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK.t21 VDD99.t495 VDD99.t494 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X981 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_22466_n8743# VSS.t551 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X982 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.t4 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VDD99.t117 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X983 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 VSS.t1631 VSS.t1630 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X984 a_25420_n13385# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 VDD99.t107 VDD99.t106 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X985 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD108.t396 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X986 a_52652_n10117# CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.t4 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB VSS.t1188 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X987 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD105.t143 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X988 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 VDD100.t180 VDD100.t179 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X989 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD90.t24 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X990 a_44253_n18696# VDD110.t496 VSS.t1012 VSS.t1011 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X991 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT a_47905_1671# VSS.t546 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X992 VDD100 RST.t38 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VDD100.t379 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X993 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD110.t135 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X994 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD100.t271 VDD100.t270 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X995 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_39690_n8887# VSS.t160 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X996 VDD96 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.JK_FF_mag_3.QB VDD96.t65 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X997 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD90.t18 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X998 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 VSS.t2464 VSS.t2463 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X999 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT RST.t39 VDD100.t378 VDD100.t377 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1000 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.t3 a_23594_n8743# VSS.t538 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1001 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t0 VDD90.t37 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1002 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VDD100.t453 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1003 a_35747_280# mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 VSS.t1275 VSS.t1274 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1004 a_47723_574# CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t5 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN VSS.t1082 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1005 a_51487_n10161# CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.t4 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT VSS.t2269 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1006 a_43719_n120# CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT a_43559_n120# VDD100.t337 pfet_03v3 ad=0.624p pd=2.92u as=0.624p ps=2.92u w=2.4u l=0.28u
X1007 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 VDD110.t47 VDD110.t45 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1008 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VDD90.t359 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1009 VDD Vdiv90.t4 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT VDD.t155 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1010 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD96.t172 VDD96.t174 VDD96.t173 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1011 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 Vdiv105.t4 VDD.t165 VDD.t164 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1012 a_51646_1671# CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t11 a_51486_1671# VSS.t1152 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1013 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t8 VDD93.t306 VDD93.t305 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1014 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t7 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VDD99.t127 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1015 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK.t22 a_48783_n13424# VSS.t2481 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1016 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 a_51028_n16724# VSS.t828 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1017 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 a_49789_n9020# VSS.t1953 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1018 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t6 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN VDD100.t224 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1019 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD93.t299 VDD93.t298 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1020 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t7 VDD100.t228 VDD100.t227 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1021 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.CLK CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VSS.t2002 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1022 a_28268_n6266# CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t8 VSS.t999 VSS.t998 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1023 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT VDD100.t437 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1024 CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD93.t188 VDD93.t187 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1025 a_47911_2768# RST.t40 a_47751_2768# VSS.t2064 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1026 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 a_53168_n2243# VSS.t1833 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1027 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB VDD110.t431 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1028 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD108.t30 VDD108.t32 VDD108.t31 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1029 VSS CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 a_28644_10099# VSS.t762 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1030 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VDD93.t236 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1031 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VDD93.t256 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1032 a_26196_5018# RST.t41 a_26036_5018# VSS.t2063 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1033 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD110.t370 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1034 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT a_53934_n9020# VSS.t645 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1035 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB VDD90.t356 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1036 a_26046_n16632# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT VSS.t243 VSS.t242 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1037 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_29777_5062# VSS.t298 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1038 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK.t23 VSS.t2483 VSS.t2482 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1039 VDD F1.t3 dec3x8_ibr_mag_0.and_3_ibr_1.nand3_mag_ibr_0.OUT VDD.t95 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1040 a_36742_n16592# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 VSS.t728 VSS.t727 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1041 dec3x8_ibr_mag_0.and_3_ibr_7.nand3_mag_ibr_0.OUT F0.t10 VDD.t170 VDD.t169 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1042 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD90.t214 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1043 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t9 VDD100.t423 VDD100.t422 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1044 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD108.t292 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1045 a_50103_5143# VDD105.t481 VSS.t1095 VSS.t1094 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1046 a_21742_n8787# VDD93.t477 VSS.t267 VSS.t266 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1047 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD96.t19 VDD96.t18 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1048 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_54751_n16684# VSS.t1363 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1049 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD99.t357 VDD99.t356 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1050 a_53216_n10117# CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t1354 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1051 a_52385_n13362# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT a_52225_n13362# VDD110.t118 pfet_03v3 ad=0.624p pd=2.92u as=0.624p ps=2.92u w=2.4u l=0.28u
X1052 dec3x8_ibr_mag_0.and_3_ibr_5.nand3_mag_ibr_0.OUT dec3x8_ibr_mag_0.and_3_ibr_5.IN3 VDD.t25 VDD.t24 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1053 a_46623_2768# CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t8 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB VSS.t1083 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1054 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN VDD93.t295 VDD93.t294 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X1055 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD90.t320 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1056 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VDD100.t17 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1057 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 VDD93.t134 VDD93.t133 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1058 VDD90 RST.t42 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD90.t272 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1059 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VDD108.t69 VDD108.t68 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1060 VDD96 CLK_div_96_mag_0.JK_FF_mag_2.Q CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD96.t323 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1061 a_45603_n5176# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t798 VSS.t797 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1062 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VSS.t1510 VSS.t1509 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1063 a_23129_n6009# CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t9 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VSS.t1172 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1064 a_25082_n17626# RST.t43 a_24922_n17626# VSS.t2062 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1065 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t4 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 VDD108.t224 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1066 a_28335_6115# VDD90.t477 VSS.t217 VSS.t216 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1067 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_25535_354# VSS.t2452 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1068 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_51439_n2199# VSS.t1283 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1069 a_26368_n2996# RST.t44 a_26208_n2996# VSS.t2061 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1070 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD96.t298 VDD96.t297 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1071 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t10 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 VDD100.t424 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1072 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_50441_n17599# VSS.t1894 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1073 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t7 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT VDD93.t439 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1074 a_25312_5018# VDD90.t478 VSS.t215 VSS.t214 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1075 a_48635_2768# CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t11 a_48475_2768# VSS.t2275 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1076 VDD96 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD96.t62 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1077 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_29834_n699# VSS.t1329 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1078 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD110.t8 VDD110.t7 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1079 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB VDD105.t254 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1080 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_48534_5187# VSS.t1775 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1081 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 F1.t4 a_37436_n1822# VSS.t1207 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1082 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_45541_n18696# VSS.t544 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1083 a_26052_n15491# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT VSS.t131 VSS.t130 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1084 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 VDD93.t172 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1085 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK VSS.t701 VSS.t700 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1086 a_24968_3016# CLK_div_96_mag_0.JK_FF_mag_4.Q.t6 CLK_div_96_mag_0.JK_FF_mag_4.QB VSS.t2283 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1087 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t12 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT VDD99.t165 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1088 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 CLK_div_93_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD93.t115 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1089 a_43760_1671# CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t4 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 VSS.t535 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1090 VDD F0.t11 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 VDD.t171 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1091 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.t2 VDD90.t179 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1092 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD100.t154 VDD100.t153 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1093 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_29116_398# VSS.t1298 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1094 a_22275_10099# CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t4 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.t2 VSS.t112 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1095 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD93.t48 VDD93.t47 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1096 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 VDD90.t384 VDD90.t383 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1097 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB VDD96.t365 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1098 a_33652_n13270# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 VDD99.t342 VDD99.t341 pfet_03v3 ad=0.624p pd=2.92u as=1.06p ps=5.68u w=2.4u l=0.28u
X1099 a_47196_n15629# CLK.t24 a_47036_n15629# VSS.t2484 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1100 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD90.t63 VDD90.t65 VDD90.t64 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1101 a_26980_3016# CLK.t25 a_26820_3016# VSS.t2485 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1102 VDD105 VDD105.t59 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT VDD105.t60 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1103 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K a_45612_1671# VSS.t69 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1104 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB VDD99.t439 VDD99.t438 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1105 VSS CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t8 a_25364_n19822# VSS.t1120 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1106 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN VSS.t410 VSS.t409 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1107 a_42521_n13474# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 VDD110.t325 VDD110.t324 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X1108 VSS VDD90.t479 a_33519_11196# VSS.t211 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1109 VSS CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN VSS.t45 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X1110 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS.t53 VSS.t52 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1111 a_41124_n16098# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 VSS.t406 VSS.t405 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1112 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN VDD99.t351 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1113 a_47270_n18696# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t5 VSS.t1247 VSS.t1246 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1114 a_50232_n7685# CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.t5 CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN VDD108.t409 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X1115 a_26811_n17626# CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.t4 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB VSS.t2355 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1116 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD100.t274 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1117 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD110.t315 VDD110.t314 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1118 a_37328_6265# F1.t5 a_37168_6265# VSS.t1208 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1119 a_43559_n120# CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 Vdiv100.t3 VDD100.t346 pfet_03v3 ad=0.624p pd=2.92u as=1.06p ps=5.68u w=2.4u l=0.28u
X1120 VDD108 VDD108.t26 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VDD108.t27 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1121 VDD96 RST.t45 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD96.t291 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1122 a_30435_n1855# CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VSS.t11 VSS.t10 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1123 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK.t26 VSS.t2487 VSS.t2486 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1124 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB VDD93.t171 VDD93.t170 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1125 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 a_51983_7381# VSS.t685 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1126 VSS CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN VSS.t12 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X1127 a_51486_1671# CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT VSS.t1838 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1128 a_46768_n5176# CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t6 a_46608_n5176# VSS.t496 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1129 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 VDD.t126 VDD.t52 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1130 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD93.t220 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1131 a_47030_n16726# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t2 VSS.t2306 VSS.t2305 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1132 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 VDD105.t292 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1133 VSS CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT a_25532_3016# VSS.t952 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1134 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 VDD100.t215 VDD100.t214 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1135 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_44324_1671# VSS.t1850 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1136 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_48478_n16682# VSS.t1766 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1137 a_45927_6284# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t815 VSS.t814 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1138 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD108.t281 VDD108.t280 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1139 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD110.t215 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1140 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t8 VDD93.t443 VDD93.t442 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1141 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VDD105.t108 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X1142 a_51849_n1102# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VSS.t1868 VSS.t1867 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1143 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 VDD93.t348 VDD93.t347 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1144 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT VDD100.t148 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1145 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB VDD93.t112 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1146 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN VDD93.t178 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X1147 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VDD93.t123 VDD93.t122 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1148 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD90.t132 VDD90.t131 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1149 dec3x8_ibr_mag_0.and_3_ibr_3.nand3_mag_ibr_0.OUT dec3x8_ibr_mag_0.and_3_ibr_3.IN1 VDD.t10 VDD.t9 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1150 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_50269_6240# VSS.t367 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1151 a_55132_5187# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t912 VSS.t911 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1152 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 a_46889_9057# VSS.t185 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1153 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t12 a_45787_574# VSS.t1081 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1154 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD100.t211 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1155 a_25806_n17626# CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t9 a_25646_n17626# VSS.t1123 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1156 a_26616_n15491# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t1858 VSS.t1857 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1157 a_29777_5062# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VSS.t195 VSS.t194 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1158 dec3x8_ibr_mag_0.and_3_ibr_1.nand3_mag_ibr_0.OUT dec3x8_ibr_mag_0.and_3_ibr_5.IN3 VDD.t23 VDD.t22 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1159 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.CLK VDD90.t17 VDD90.t16 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1160 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD90.t127 VDD90.t126 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1161 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t9 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT VDD100.t229 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1162 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD99.t240 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1163 VDD F1.t6 dec3x8_ibr_mag_0.and_3_ibr_7.nand3_mag_ibr_0.OUT VDD.t98 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1164 CLK_div_96_mag_0.JK_FF_mag_5.QB CLK_div_96_mag_0.JK_FF_mag_5.Q.t5 VDD96.t116 VDD96.t115 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1165 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD99.t316 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1166 VSS VDD105.t483 a_45730_10154# VSS.t1096 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1167 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_52811_1671# VSS.t1881 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1168 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD110.t81 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1169 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD90.t143 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1170 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD100.t7 VDD100.t6 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1171 a_39844_n10028# RST.t46 a_39684_n10028# VSS.t2060 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1172 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.CLK CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VDD105.t304 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1173 a_37328_6821# F1.t7 a_37168_6821# VSS.t1208 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1174 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT a_47911_2768# VSS.t672 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1175 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD93.t251 VDD93.t250 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1176 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_25478_6115# VSS.t135 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1177 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_96_mag_0.JK_FF_mag_0.QB a_22424_n1833# VSS.t416 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1178 a_22988_n1789# CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS.t23 VSS.t22 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1179 a_23706_n2886# CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS.t1741 VSS.t1740 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1180 a_22685_11196# CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t652 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1181 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.t5 VDD90.t224 VDD90.t223 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1182 a_30496_10099# CLK.t27 a_30336_10099# VSS.t2488 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1183 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_47492_n5176# VSS.t1030 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1184 a_45075_n9063# CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t4 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VSS.t992 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1185 a_21995_n7106# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VSS.t720 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1186 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD105.t28 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1187 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 F1.t8 a_37436_880# VSS.t1209 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1188 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT CLK.t28 VDD108.t443 VDD108.t442 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1189 a_48475_2768# CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t10 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT VSS.t1084 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1190 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD96.t169 VDD96.t171 VDD96.t170 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1191 a_21857_810# CLK_div_96_mag_0.JK_FF_mag_5.Q.t6 CLK_div_96_mag_0.JK_FF_mag_5.QB VSS.t1062 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1192 Vdiv93 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VDD93.t318 VDD93.t317 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1193 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD100.t8 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1194 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VDD96.t300 VDD96.t299 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1195 a_51040_10154# RST.t47 a_50880_10154# VSS.t2059 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1196 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_48832_n1102# VSS.t877 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1197 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD108.t199 VDD108.t198 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1198 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 VDD93.t150 VDD93.t149 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1199 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD108.t205 VDD108.t204 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1200 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K VDD100.t283 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1201 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K VDD99.t388 VDD99.t387 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1202 a_23019_5018# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS.t1033 VSS.t1032 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1203 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.t8 VDD99.t80 VDD99.t79 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1204 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 VDD93.t308 VDD93.t307 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1205 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB VDD100.t176 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1206 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD96.t166 VDD96.t168 VDD96.t167 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1207 VSS CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t3 a_35186_n18723# VSS.t2371 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1208 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.t5 VSS.t2221 VSS.t2220 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X1209 a_44321_n6273# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS.t2135 VSS.t146 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1210 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD108.t23 VDD108.t25 VDD108.t24 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1211 CLK_div_90_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_90_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VDD90.t84 VDD90.t83 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X1212 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB VDD90.t210 VDD90.t209 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1213 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD110.t212 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1214 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK VDD93.t216 VDD93.t215 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1215 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 VDD93.t372 VDD93.t371 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1216 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 VDD105.t142 VDD105.t141 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1217 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN VSS.t1350 VSS.t1349 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1218 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD110.t69 VDD110.t68 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1219 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN VSS.t920 VSS.t918 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X1220 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD96.t109 VDD96.t108 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1221 VDD110 dec3x8_ibr_mag_0.and_3_ibr_7.nand3_mag_ibr_0.OUT VDD.t58 VDD.t57 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1222 a_44517_n10160# RST.t48 a_44357_n10160# VSS.t2058 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1223 VDD96 CLK_div_96_mag_0.JK_FF_mag_0.QB CLK_div_96_mag_0.JK_FF_mag_0.Q VDD96.t38 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1224 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD93.t169 VDD93.t168 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1225 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_108_new_mag_0.JK_FF_mag_1.QB a_50111_n5768# VSS.t2318 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1226 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_3.Q VDD96.t61 VDD96.t60 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1227 a_33583_n16588# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 VSS.t1399 VSS.t1398 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1228 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t13 VSS.t1169 VSS.t1168 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1229 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD90.t202 VDD90.t201 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1230 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t9 VDD93.t445 VDD93.t444 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1231 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 VDD93.t148 VDD93.t147 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1232 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD105.t209 VDD105.t208 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1233 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t13 VDD100.t246 VDD100.t245 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1234 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_44894_2768# VSS.t26 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1235 a_34730_n16636# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K VSS.t2169 VSS.t2168 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1236 dec3x8_ibr_mag_0.and_3_ibr_7.nand3_mag_ibr_0.OUT F0.t12 a_39580_6265# VSS.t276 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1237 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_30025_n2952# VSS.t1829 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1238 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD110.t416 VDD110.t415 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1239 a_55019_7683# CLK_div_105_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 VDD105.t88 VDD105.t87 pfet_03v3 ad=0.624p pd=2.92u as=1.06p ps=5.68u w=2.4u l=0.28u
X1240 a_44123_n1146# CLK.t29 a_43963_n1146# VSS.t2489 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1241 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_36178_n16592# VSS.t1369 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1242 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT RST.t49 VDD90.t276 VDD90.t275 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1243 a_28828_1497# CLK_div_96_mag_0.JK_FF_mag_3.Q VSS.t442 VSS.t441 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1244 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_23179_5018# VSS.t950 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1245 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K VDD110.t279 VDD110.t278 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1246 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_43947_n9019# VSS.t1489 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1247 a_37168_6265# dec3x8_ibr_mag_0.and_3_ibr_5.IN3 VSS.t360 VSS.t358 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1248 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD100.t331 VDD100.t330 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1249 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD100.t310 VDD100.t309 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1250 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 a_26206_n16632# VSS.t1856 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1251 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD110.t226 VDD110.t225 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1252 a_30317_n18723# CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t4 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.t2 VSS.t2370 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1253 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 VDD108.t323 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1254 VSS VDD90.t480 a_27150_11196# VSS.t208 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1255 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD96.t101 VDD96.t100 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1256 a_33744_n17626# CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t1641 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1257 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB VDD110.t209 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1258 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VDD90.t198 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1259 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VDD99.t32 VDD99.t31 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1260 a_53850_6284# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS.t1549 VSS.t1548 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1261 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_50721_n1102# VSS.t92 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1262 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t0 VDD100.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1263 a_46980_n1146# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t4 VSS.t1175 VSS.t1174 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1264 a_47698_n2243# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VSS.t369 VSS.t368 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1265 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 VDD90.t87 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1266 VDD93 dec3x8_ibr_mag_0.and_3_ibr_4.nand3_mag_ibr_0.OUT VSS.t100 VSS.t99 nfet_03v3 ad=0.157p pd=1.68u as=0.152p ps=1.64u w=0.22u l=0.28u
X1267 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VDD100.t116 VDD100.t115 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1268 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD99.t508 VDD99.t507 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1269 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t1 VDD99.t425 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1270 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.t4 VDD108.t403 VDD108.t402 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1271 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD105.t183 VDD105.t182 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1272 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_54057_10154# VSS.t1442 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1273 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 F0.t13 a_36310_880# VSS.t2442 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1274 VDD108 CLK_div_108_new_mag_0.JK_FF_mag_1.Q CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD108.t418 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1275 a_29208_10099# CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t57 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1276 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t5 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VDD99.t466 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1277 VDD F1.t9 dec3x8_ibr_mag_0.and_3_ibr_3.nand3_mag_ibr_0.OUT VDD.t101 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1278 VDD F2.t2 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 VDD.t73 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1279 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t6 CLK_div_108_new_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN VDD108.t383 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1280 CLK_div_105_mag_0.CLK_div_10_mag_1.CLK CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 a_55179_7683# VDD105.t304 pfet_03v3 ad=1.06p pd=5.68u as=0.624p ps=2.92u w=2.4u l=0.28u
X1281 a_50269_6240# CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 a_50109_6240# VSS.t684 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1282 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.t6 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD99.t474 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1283 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD108.t154 VDD108.t153 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1284 a_32789_10099# CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t483 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1285 a_46889_9057# CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t2 VSS.t569 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1286 VDD100 VDD100.t89 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VDD100.t90 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1287 VDD110 RST.t50 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT VDD110.t401 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1288 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VDD105.t8 VDD105.t7 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1289 a_29862_n9832# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 VSS.t383 VSS.t382 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1290 a_22455_5018# CLK_div_90_mag_0.CLK_div_10_mag_0.CLK a_22295_5018# VSS.t96 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1291 a_37955_n9984# CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t381 VSS.t380 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1292 a_49752_10154# CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t8 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB VSS.t1226 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1293 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS.t604 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X1294 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD96.t143 VDD96.t142 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1295 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_43606_2768# VSS.t2 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1296 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 VDD90.t100 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1297 VDD mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT VDD.t54 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1298 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 VDD105.t77 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1299 dec3x8_ibr_mag_0.and_3_ibr_3.nand3_mag_ibr_0.OUT dec3x8_ibr_mag_0.and_3_ibr_3.IN1 a_39580_6821# VSS.t276 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1300 a_24512_n18723# CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t1638 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1301 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD108.t330 VDD108.t329 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1302 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_45927_6284# VSS.t2122 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1303 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB VDD100.t204 VDD100.t203 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1304 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD100.t301 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1305 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_96_mag_0.JK_FF_mag_3.Q a_28737_n2996# VSS.t440 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1306 a_46614_n6273# CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 VSS.t1617 VSS.t493 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1307 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB a_26636_n8734# VSS.t21 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1308 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t10 a_29214_n6271# VSS.t1665 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1309 VSS VDD105.t484 a_48741_9057# VSS.t1099 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1310 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD100.t145 VDD100.t144 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1311 a_45969_n2199# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t320 VSS.t319 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1312 a_37168_6821# dec3x8_ibr_mag_0.and_3_ibr_5.IN3 VSS.t359 VSS.t358 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1313 a_29213_n7028# CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 VSS.t144 VSS.t143 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1314 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD96.t12 VDD96.t11 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1315 a_49488_n13383# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 VSS.t404 VSS.t403 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1316 a_25478_6115# CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 a_25318_6115# VSS.t1629 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1317 a_51551_5187# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VSS.t306 VSS.t305 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1318 VSS VDD100.t483 a_45618_2768# VSS.t2400 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1319 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD100.t112 VDD100.t111 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1320 VSS CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN VSS.t34 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X1321 VSS VDD93.t478 a_26343_n7107# VSS.t263 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1322 VSS CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_25625_n6010# VSS.t1413 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1323 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_26778_n1855# VSS.t1698 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1324 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD110.t38 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1325 VDD100 VDD100.t85 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VDD100.t86 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1326 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT RST.t51 VDD100.t376 VDD100.t375 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1327 a_24127_10099# CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t8 a_23967_10099# VSS.t1178 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1328 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t10 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VSS.t2207 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1329 VDD100 CLK.t30 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD100.t470 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1330 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 VSS.t469 VSS.t468 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X1331 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT VDD105.t322 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1332 a_47134_n2243# CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 a_46974_n2243# VSS.t2462 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1333 a_34308_n17626# CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VSS.t1273 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1334 a_52293_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VSS.t1889 VSS.t1888 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1335 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_44055_n16724# VSS.t557 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1336 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VDD90.t125 VDD90.t124 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1337 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 a_47453_9057# VSS.t1538 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1338 a_46400_n9019# CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.t2 VSS.t738 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1339 a_50715_n2243# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VSS.t1752 VSS.t1751 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1340 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD100.t57 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1341 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD90.t13 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1342 a_29181_n16634# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT VSS.t2137 VSS.t2136 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1343 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD99.t272 VDD99.t271 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1344 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT Vdiv90.t5 a_35747_n1222# VSS.t759 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1345 a_31737_n15535# CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t14 a_31577_n15535# VSS.t1170 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1346 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_23030_n8743# VSS.t678 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1347 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 VDD90.t146 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1348 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t7 VDD105.t96 VDD105.t95 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1349 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_45753_n15583# VSS.t964 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1350 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT VDD110.t170 VDD110.t169 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X1351 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t7 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD108.t93 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1352 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 VDD108.t373 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1353 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD110.t236 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1354 a_32225_10099# CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t49 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1355 a_49991_n2243# VDD100.t485 VSS.t2404 VSS.t2403 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1356 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 a_30165_n6282# VSS.t450 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1357 a_54978_6284# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t1609 VSS.t1608 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1358 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 VDD100.t312 VDD100.t311 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1359 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD110.t18 VDD110.t20 VDD110.t19 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1360 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 VDD100.t141 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1361 a_24391_n20290# CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.t7 CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VDD99.t477 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X1362 a_30315_n15493# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t603 VSS.t602 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1363 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD99.t396 VDD99.t395 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1364 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t14 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 VSS.t1155 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1365 a_30342_11196# CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.t6 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VSS.t1077 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1366 VDD96 CLK_div_96_mag_0.JK_FF_mag_3.QB CLK_div_96_mag_0.JK_FF_mag_3.Q VDD96.t76 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1367 a_44894_2768# RST.t52 a_44734_2768# VSS.t2057 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1368 VDD108 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD108.t253 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1369 VDD108 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD108.t431 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1370 VSS CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t1 VSS.t170 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1371 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD110.t269 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1372 a_39580_6265# F1.t10 a_39420_6265# VSS.t1210 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1373 VSS CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_0.OUT a_23139_n287# VSS.t1277 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1374 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 VDD100.t452 VDD100.t451 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1375 a_26965_n18723# CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.t2 VSS.t1408 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1376 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB VDD105.t138 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1377 a_23179_5018# RST.t53 a_23019_5018# VSS.t2056 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1378 VDD108 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD108.t310 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1379 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS.t1771 VSS.t1770 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X1380 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VDD93.t359 VDD93.t358 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1381 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_26072_n8734# VSS.t457 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1382 a_29618_11196# CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VSS.t1434 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1383 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD96.t201 VDD96.t200 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1384 a_45405_n2199# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS.t1522 VSS.t1521 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1385 CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.t5 VSS.t1074 VSS.t1073 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X1386 VSS CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t6 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN VSS.t2363 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X1387 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_26760_5062# VSS.t111 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1388 a_25076_n18723# CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t990 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1389 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 a_52806_n9020# VSS.t799 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1390 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t9 VDD93.t276 VDD93.t275 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1391 a_47835_7960# CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t8 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN VSS.t488 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1392 a_23703_n287# CLK_div_96_mag_0.JK_FF_mag_5.QB CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_0.OUT VSS.t64 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1393 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K VDD100.t156 VDD100.t155 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1394 a_54022_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS.t618 VSS.t617 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1395 mux_8x1_ibr_0.mux_2x1_ibr_0.I0 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 VDD.t132 VDD.t131 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1396 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD90.t99 VDD90.t98 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1397 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_49276_n17599# VSS.t874 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1398 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT VDD110.t414 VDD110.t413 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1399 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD90.t184 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1400 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VDD99.t296 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1401 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 mux_8x1_ibr_0.mux_2x1_ibr_0.I1 VDD.t146 VDD.t145 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1402 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 VDD99.t350 VDD99.t349 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1403 a_55179_7683# CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT a_55019_7683# VDD105.t463 pfet_03v3 ad=0.624p pd=2.92u as=0.624p ps=2.92u w=2.4u l=0.28u
X1404 VSS CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.t5 a_25800_n18723# VSS.t2356 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1405 a_28734_n9876# RST.t54 a_28574_n9876# VSS.t2055 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1406 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 a_31506_5018# VSS.t1811 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1407 a_53174_n1146# CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 a_53014_n1146# VSS.t2461 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1408 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD108.t188 VDD108.t187 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1409 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VDD105.t265 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1410 VSS CLK_div_99_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 VSS.t739 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1411 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT CLK.t31 VDD108.t445 VDD108.t444 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1412 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD108.t44 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1413 a_22295_5018# VDD90.t481 VSS.t207 VSS.t206 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1414 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 VDD99.t68 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1415 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD93.t1 VDD93.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1416 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB VDD105.t227 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1417 a_26420_10099# CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t112 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1418 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VDD90.t139 VDD90.t138 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1419 VDD96 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD96.t212 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1420 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 VDD99.t449 VDD99.t448 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1421 VDD90 dec3x8_ibr_mag_0.and_3_ibr_0.nand3_mag_ibr_0.OUT VDD.t27 VDD.t26 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1422 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t5 VDD100.t250 VDD100.t249 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1423 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_2.Q VDD96.t322 VDD96.t321 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1424 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 VDD108.t334 VDD108.t333 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1425 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t1 VSS.t31 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1426 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t4 VDD105.t214 VDD105.t213 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1427 a_39580_6821# F1.t11 a_39420_6821# VSS.t1210 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1428 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 a_44779_n16724# VSS.t480 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1429 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD110.t256 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1430 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD108.t366 VDD108.t365 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1431 a_31507_11196# CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.t6 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB VSS.t757 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1432 a_23748_n9840# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t707 VSS.t706 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1433 a_44407_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.CLK a_44247_n17599# VSS.t543 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1434 a_31445_n18723# CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t1150 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1435 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t4 VDD90.t229 VDD90.t228 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1436 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_33019_n16588# VSS.t1397 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1437 a_53940_n10161# RST.t55 a_53780_n10161# VSS.t2054 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1438 a_54414_6284# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t1836 VSS.t1835 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1439 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_3.Q VSS.t439 VSS.t438 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1440 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.t6 VDD108.t110 VDD108.t109 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1441 a_51803_n5724# CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t1295 VSS.t1294 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1442 CLK_div_90_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT VSS.t385 VSS.t384 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X1443 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VDD105.t156 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1444 dec3x8_ibr_mag_0.and_3_ibr_4.nand3_mag_ibr_0.OUT dec3x8_ibr_mag_0.and_3_ibr_6.IN3 VDD.t51 VDD.t50 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1445 a_54664_n10161# CLK.t32 a_54504_n10161# VSS.t2490 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1446 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB VDD93.t235 VDD93.t234 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1447 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_27227_398# VSS.t2451 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1448 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VDD105.t274 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1449 VDD105 RST.t56 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD105.t399 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1450 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.CLK VDD100.t360 VDD100.t359 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1451 a_32635_11196# CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VSS.t1530 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1452 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 a_52003_n2199# VSS.t1035 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1453 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT VSS.t104 VSS.t103 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1454 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 VDD110.t361 VDD110.t360 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1455 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_29059_6159# VSS.t193 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1456 VDD96 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 VDD96.t193 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1457 VSS CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_33180_n17626# VSS.t1931 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1458 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_51165_n17599# VSS.t668 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1459 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VSS.t1504 VSS.t1503 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1460 a_22544_n13819# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 VSS.t2341 VSS.t2340 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1461 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT VDD93.t338 VDD93.t337 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1462 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT VDD93.t190 VDD93.t189 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1463 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t11 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD93.t446 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1464 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD110.t252 VDD110.t251 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1465 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD110.t78 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1466 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_32230_5018# VSS.t473 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1467 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VSS.t59 VSS.t58 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1468 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t11 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VDD105.t452 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1469 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD99.t214 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1470 a_29623_6159# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VSS.t198 VSS.t197 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1471 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT VDD105.t249 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1472 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD105.t4 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1473 a_41117_n13911# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 VSS.t402 VSS.t401 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1474 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK.t33 VDD90.t453 VDD90.t452 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1475 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VDD100.t364 VDD100.t363 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1476 a_35747_880# mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 VSS.t1645 VSS.t1274 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1477 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.t9 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VDD99.t81 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1478 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 a_43751_n5176# VSS.t1616 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1479 VDD99 RST.t57 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT VDD99.t365 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1480 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_29751_n15493# VSS.t54 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1481 VSS CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 a_21277_n6009# VSS.t2018 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1482 a_43718_10154# CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K VSS.t1820 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1483 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD96.t277 VDD96.t276 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1484 VDD110 CLK.t34 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT VDD110.t466 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1485 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VDD105.t371 VDD105.t370 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1486 a_52115_5187# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VSS.t580 VSS.t579 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1487 a_25662_n9875# RST.t58 a_25502_n9875# VSS.t2053 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1488 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 a_43872_9057# VSS.t332 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1489 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD90.t300 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1490 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 a_31177_7256# VSS.t1336 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1491 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t4 VDD96.t330 VDD96.t329 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1492 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD93.t297 VDD93.t296 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1493 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD96.t33 VDD96.t32 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1494 VSS CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_23948_n18723# VSS.t1817 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1495 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t6 VDD110.t190 VDD110.t189 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1496 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN VDD110.t57 VDD110.t56 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1497 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 VDD105.t429 VDD105.t428 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1498 a_26760_5062# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VSS.t1421 VSS.t1420 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1499 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 VDD108.t168 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1500 VSS CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN VSS.t5 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X1501 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VDD90.t1 VDD90.t0 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1502 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 a_48620_n5176# VSS.t311 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1503 VSS CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_27375_n17626# VSS.t890 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1504 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT RST.t59 VDD108.t353 VDD108.t352 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1505 a_50150_n15627# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K VSS.t1410 VSS.t1409 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1506 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT VDD100.t304 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1507 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD90.t407 VDD90.t406 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1508 a_48587_10154# CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t9 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT VSS.t491 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1509 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_96_mag_0.JK_FF_mag_2.Q a_25644_n2996# VSS.t2157 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1510 a_32865_n15491# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 VSS.t2101 VSS.t2100 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1511 a_36109_n8931# CLK_div_93_mag_0.CLK_div_3_mag_0.CLK a_35949_n8931# VSS.t699 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1512 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_2.OUT Vdiv108.t4 a_53249_n6862# VSS.t1184 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1513 a_52161_n19793# CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 VSS.t1893 VSS.t868 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1514 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD100.t28 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1515 a_47754_n16726# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT VSS.t766 VSS.t765 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1516 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 VDD108.t291 VDD108.t290 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1517 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t5 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VDD108.t179 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1518 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t12 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 VDD105.t455 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1519 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_22461_6115# VSS.t1020 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1520 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t10 VDD99.t131 VDD99.t130 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1521 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 VSS.t1979 VSS.t1978 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X1522 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 a_47246_5143# VSS.t683 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1523 a_42529_n14305# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 VSS.t1804 VSS.t399 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1524 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD105.t170 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1525 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD93.t324 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1526 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VDD93.t349 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1527 a_38966_n8931# CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 VSS.t286 VSS.t285 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1528 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD93.t94 VDD93.t96 VDD93.t95 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1529 VDD110 dec3x8_ibr_mag_0.and_3_ibr_7.nand3_mag_ibr_0.OUT VSS.t1021 VSS.t610 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1530 a_51575_n18696# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VSS.t667 VSS.t666 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1531 VSS CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_23409_11196# VSS.t614 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1532 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT VSS.t1653 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1533 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT VDD99.t72 VDD99.t71 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X1534 VSS CLK.t35 a_51205_n7921# VSS.t2491 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1535 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_27180_n15491# VSS.t969 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1536 a_47810_5143# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VSS.t980 VSS.t979 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1537 a_43901_n15627# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K VSS.t1375 VSS.t1374 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1538 a_42083_n15712# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 VDD110.t28 VDD110.t27 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X1539 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 VSS.t770 VSS.t769 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X1540 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD100.t448 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1541 VDD99 VDD99.t48 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VDD99.t49 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1542 VDD99 CLK.t36 CLK_div_99_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN VDD99.t496 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1543 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 VDD.t128 VDD.t127 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1544 a_43957_n2243# VDD100.t486 VSS.t2406 VSS.t2405 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1545 VSS CLK_div_90_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 VSS.t595 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1546 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB VDD105.t222 VDD105.t221 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1547 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 a_27324_5062# VSS.t132 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1548 dec3x8_ibr_mag_0.and_3_ibr_0.nand3_mag_ibr_0.OUT dec3x8_ibr_mag_0.and_3_ibr_5.IN3 VDD.t21 VDD.t20 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1549 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD99.t198 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1550 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 VDD105.t427 VDD105.t426 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1551 VDD96 RST.t60 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VDD96.t288 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1552 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT a_50316_10154# VSS.t1384 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1553 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t12 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN VDD100.t427 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1554 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t7 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VSS.t2233 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1555 a_26189_n6010# CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t10 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VSS.t1000 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1556 a_25138_11196# CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.t7 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB VSS.t1182 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1557 a_24270_n2886# CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t1649 VSS.t1648 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1558 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VDD99.t57 VDD99.t56 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X1559 a_49951_n5768# VDD108.t461 VSS.t518 VSS.t517 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1560 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT RST.t61 VDD105.t398 VDD105.t397 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1561 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD105.t187 VDD105.t186 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1562 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K VDD105.t3 VDD105.t2 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1563 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT a_50199_n10117# VSS.t1897 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1564 a_29059_6159# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VSS.t241 VSS.t240 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1565 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 VDD96.t28 VDD96.t27 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1566 a_34462_n18723# CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t1930 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1567 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VSS.t582 VSS.t581 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1568 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 VDD108.t116 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1569 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_47970_5143# VSS.t838 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1570 a_28099_n17626# RST.t62 a_27939_n17626# VSS.t2052 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1571 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD110.t101 VDD110.t100 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1572 VDD110 CLK.t37 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT VDD110.t469 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1573 VDD96 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_0.OUT CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.IN1 VDD96.t128 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1574 a_51604_10154# CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t9 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT VSS.t1227 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1575 CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t6 a_54866_n1102# VSS.t1176 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1576 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD108.t201 VDD108.t200 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1577 CLK_div_108_new_mag_0.JK_FF_mag_0.QB CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD108.t61 VDD108.t60 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1578 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD100.t107 VDD100.t106 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1579 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT VDD99.t239 VDD99.t238 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1580 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 a_53458_n17599# VSS.t2108 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1581 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 a_31731_n16632# VSS.t2339 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1582 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 VDD93.t346 VDD93.t345 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1583 VSS CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.VOUT CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN VSS.t138 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X1584 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_48558_n18696# VSS.t396 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1585 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t7 VDD110.t456 VDD110.t455 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1586 a_50833_6284# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VSS.t2085 VSS.t2084 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1587 VDD96 CLK_div_96_mag_0.JK_FF_mag_5.QB CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_0.OUT VDD96.t6 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1588 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_50829_n6865# VSS.t1393 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1589 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t5 CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 VDD105.t190 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1590 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT VDD99.t197 VDD99.t196 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1591 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 F0.t14 VSS.t2444 VSS.t2443 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1592 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 a_48023_n7840# VDD108.t67 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X1593 a_52839_n5# CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 VSS.t2460 VSS.t2459 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1594 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD108.t259 VDD108.t258 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1595 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN VDD99.t207 VDD99.t206 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1596 a_45241_n10160# CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t8 a_45081_n10160# VSS.t2236 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1597 VDD dec3x8_ibr_mag_0.and_3_ibr_5.IN3 dec3x8_ibr_mag_0.and_3_ibr_4.nand3_mag_ibr_0.OUT VDD.t17 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1598 VSS VDD99.t513 a_28823_n17626# VSS.t2429 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1599 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_51592_n16680# VSS.t1782 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1600 a_44841_n2243# RST.t63 a_44681_n2243# VSS.t2051 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1601 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD105.t285 VDD105.t284 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1602 VSS CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t0 VSS.t1956 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1603 a_43872_9057# CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t5 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 VSS.t1071 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1604 a_31177_7256# CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 VSS.t1628 VSS.t1627 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1605 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 VSS.t1325 VSS.t1324 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1606 a_35454_n16636# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT VSS.t63 VSS.t62 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1607 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD93.t144 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1608 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT RST.t64 VDD105.t396 VDD105.t395 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1609 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_53463_n16728# VSS.t1803 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1610 a_26042_6159# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VSS.t1269 VSS.t1268 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1611 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_96_mag_0.JK_FF_mag_0.Q a_22418_n2930# VSS.t1694 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1612 a_55161_n15587# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 VSS.t902 VSS.t901 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1613 VSS CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_25702_11196# VSS.t342 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1614 VDD96 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_0.OUT CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 VDD96.t22 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1615 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD100.t298 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1616 VDD mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 VDD.t114 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1617 a_26250_1919# CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 VSS.t951 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1618 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT VSS.t1360 VSS.t1359 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X1619 a_51193_n19793# CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 VSS.t873 VSS.t868 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1620 a_36042_6265# dec3x8_ibr_mag_0.and_3_ibr_6.IN3 VSS.t786 VSS.t356 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1621 a_48324_n15585# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t1676 VSS.t1675 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1622 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K a_45724_9057# VSS.t777 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1623 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN VDD93.t13 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X1624 VDD96 CLK_div_96_mag_0.JK_FF_mag_4.QB CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_0.OUT VDD96.t46 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1625 a_37391_n9984# CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS.t190 VSS.t189 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1626 a_36673_n8887# CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS.t51 VSS.t50 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1627 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 F1.t12 VSS.t1212 VSS.t1211 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1628 a_22461_6115# CLK_div_90_mag_0.CLK_div_10_mag_0.CLK a_22301_6115# VSS.t95 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1629 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 VDD108.t237 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1630 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_47338_n6273# VSS.t146 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1631 dec3x8_ibr_mag_0.and_3_ibr_5.IN3 F2.t3 VSS.t1200 VSS.t1199 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1632 a_40972_n9984# CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t1962 VSS.t1961 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1633 a_52769_10154# CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t13 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB VSS.t2210 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1634 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VSS.t395 VSS.t394 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1635 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD100.t445 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1636 VDD99 CLK.t38 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VDD99.t499 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1637 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD110.t357 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1638 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.JK_FF_mag_4.QB VDD96.t45 VDD96.t44 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1639 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD99.t252 VDD99.t251 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1640 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD100.t294 VDD100.t293 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1641 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD100.t56 VDD100.t55 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1642 VDD105 RST.t65 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD105.t392 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1643 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VSS.t986 VSS.t985 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1644 VDD96 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD96.t209 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1645 a_41284_n14596# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_41124_n14596# VSS.t1802 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1646 a_51598_9057# CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT VSS.t1308 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1647 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD110.t253 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1648 VDD108 CLK_div_108_new_mag_0.JK_FF_mag_1.QB CLK_div_108_new_mag_0.JK_FF_mag_1.Q VDD108.t428 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1649 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD96.t163 VDD96.t165 VDD96.t164 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1650 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_47534_n10160# VSS.t921 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1651 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_51397_6284# VSS.t1839 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1652 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD100.t173 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1653 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD100.t22 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1654 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD100.t82 VDD100.t84 VDD100.t83 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1655 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_47140_n1146# VSS.t876 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1656 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD90.t282 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1657 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD90.t385 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1658 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VDD99.t308 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1659 VDD96 VDD96.t159 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_0.OUT VDD96.t160 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1660 a_29461_n2996# RST.t66 a_29301_n2996# VSS.t2050 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1661 a_36103_n10028# CLK_div_93_mag_0.CLK_div_3_mag_0.CLK a_35943_n10028# VSS.t698 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1662 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 a_43383_n9019# VSS.t1913 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1663 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VSS.t235 VSS.t234 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1664 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_52156_n16680# VSS.t400 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1665 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN VSS.t199 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X1666 VDD Vdiv108.t5 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT VDD.t28 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1667 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 VSS.t882 VSS.t881 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1668 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD105.t12 VDD105.t11 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1669 a_51961_6284# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VSS.t180 VSS.t179 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1670 VDD108 dec3x8_ibr_mag_0.and_3_ibr_3.nand3_mag_ibr_0.OUT VDD.t34 VDD.t33 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1671 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 VDD108.t289 VDD108.t288 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1672 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 VDD99.t265 VDD99.t264 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1673 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 VDD99.t424 VDD99.t423 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1674 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT VDD105.t150 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1675 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_93_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD93.t249 VDD93.t248 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1676 a_36042_6821# dec3x8_ibr_mag_0.and_3_ibr_5.IN3 VSS.t357 VSS.t277 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1677 CLK_div_96_mag_0.JK_FF_mag_2.Q CLK_div_96_mag_0.JK_FF_mag_2.QB a_27342_n1855# VSS.t2333 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1678 VSS CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_33334_n18723# VSS.t1642 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1679 VDD mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I1 VDD.t188 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1680 Vdiv108 CLK_div_108_new_mag_0.JK_FF_mag_0.QB a_54947_n5721# VSS.t1047 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1681 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 VDD105.t380 VDD105.t379 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1682 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 VSS.t2118 VSS.t2117 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1683 a_54187_n16728# RST.t67 a_54027_n16728# VSS.t2049 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1684 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT VDD110.t232 VDD110.t231 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1685 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_26606_6159# VSS.t110 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1686 VDD96 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_4.IN2 CLK_div_96_mag_0.JK_FF_mag_5.QB VDD96.t41 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1687 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD99.t506 VDD99.t505 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1688 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD110.t345 VDD110.t344 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1689 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.t7 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VDD90.t171 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1690 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_32301_n15491# VSS.t2104 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1691 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VSS.t2303 VSS.t2302 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1692 a_28644_10099# CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t4 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.t0 VSS.t742 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1693 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_23743_5062# VSS.t2255 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1694 a_48629_1671# CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t13 a_48469_1671# VSS.t2276 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1695 VDD dec3x8_ibr_mag_0.and_3_ibr_6.IN3 dec3x8_ibr_mag_0.and_3_ibr_0.nand3_mag_ibr_0.OUT VDD.t47 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1696 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_108_new_mag_0.JK_FF_mag_1.QB VDD108.t427 VDD108.t426 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1697 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_47190_n16726# VSS.t2187 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1698 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t0 VDD108.t64 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1699 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 VDD99.t446 VDD99.t445 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1700 dec3x8_ibr_mag_0.and_3_ibr_6.nand3_mag_ibr_0.OUT F0.t15 VDD.t175 VDD.t174 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1701 a_50447_n18696# CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_50287_n18696# VSS.t872 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1702 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t11 VDD99.t133 VDD99.t132 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1703 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 a_47914_n16726# VSS.t1674 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1704 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_5.Q.t7 VSS.t1064 VSS.t1063 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1705 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_48888_n15585# VSS.t2192 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1706 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK.t39 VSS.t2495 VSS.t2494 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1707 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 VDD105.t257 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1708 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 a_30398_n699# VSS.t2153 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1709 a_30469_n16590# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t1885 VSS.t1884 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1710 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN VSS.t151 VSS.t150 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1711 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 VDD99.t139 VDD99.t138 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1712 a_43229_n10116# CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.t6 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K VSS.t2222 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1713 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_51011_n18696# VSS.t1575 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1714 a_25328_n15535# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K VSS.t182 VSS.t181 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1715 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t5 a_31512_6115# VSS.t1159 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1716 a_30210_n13332# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 a_30050_n13332# VSS.t1582 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1717 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t12 a_26790_n9831# VSS.t1005 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1718 a_47341_1671# CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 VSS.t943 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1719 VSS CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_4.IN2 a_21857_810# VSS.t417 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1720 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 VDD110.t90 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1721 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT VDD105.t309 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1722 a_50304_n16724# CLK.t40 a_50144_n16724# VSS.t2496 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1723 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_54033_n15587# VSS.t2309 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1724 a_48258_n10160# CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t9 a_48098_n10160# VSS.t2237 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1725 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT VDD100.t41 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1726 a_25490_n1899# VDD96.t382 VSS.t1463 VSS.t1462 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1727 a_51439_n2199# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VSS.t91 VSS.t90 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1728 a_26208_n2996# CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VSS.t30 VSS.t29 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1729 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VDD93.t266 VDD93.t265 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1730 a_44953_5143# RST.t68 a_44793_5143# VSS.t2048 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1731 a_53129_n19793# CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 VSS.t1323 VSS.t1322 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1732 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.t3 a_28010_n9876# VSS.t126 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1733 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VSS.t353 VSS.t352 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1734 a_37436_n1822# mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I1 VSS.t1780 VSS.t1779 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1735 a_52002_n15583# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 VSS.t467 VSS.t466 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1736 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD110.t103 VDD110.t102 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1737 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD93.t418 VDD93.t417 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1738 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 F2.t4 VSS.t1202 VSS.t1201 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1739 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB VDD99.t443 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1740 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.t8 VDD99.t479 VDD99.t478 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1741 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB VDD110.t150 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1742 a_21896_n9884# CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t10 a_21736_n9884# VSS.t1173 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1743 CLK_div_93_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_3_mag_0.CLK VDD93.t214 VDD93.t213 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1744 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 Vdiv99.t3 VDD.t163 VDD.t162 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1745 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t11 VDD93.t278 VDD93.t277 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1746 a_36827_n10028# RST.t69 a_36667_n10028# VSS.t2047 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1747 a_53892_n2243# RST.t70 a_53732_n2243# VSS.t2046 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1748 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN VDD99.t144 VDD99.t143 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1749 a_49635_n10117# CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.t6 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K VSS.t2270 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1750 VSS CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_33898_n18723# VSS.t1270 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1751 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD110.t147 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1752 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.t4 a_28267_n7033# VSS.t125 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1753 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT VDD105.t325 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1754 VDD96 CLK_div_96_mag_0.JK_FF_mag_5.Q.t8 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_2.OUT VDD96.t117 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1755 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VDD99.t435 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1756 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_26042_6159# VSS.t1419 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1757 a_30341_5062# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VSS.t2251 VSS.t2250 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1758 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_96_mag_0.JK_FF_mag_3.Q VDD96.t59 VDD96.t58 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1759 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_105_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 VDD105.t111 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X1760 Vdiv110 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 a_55357_n20487# VDD110.t419 pfet_03v3 ad=1.06p pd=5.68u as=0.624p ps=2.92u w=2.4u l=0.28u
X1761 a_24938_n9875# CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 a_24778_n9875# VSS.t449 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1762 a_33519_11196# CLK.t41 a_33359_11196# VSS.t2497 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1763 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD99.t394 VDD99.t393 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1764 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t10 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT VDD105.t237 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1765 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t5 a_28552_354# VSS.t2202 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1766 a_36202_6265# dec3x8_ibr_mag_0.and_3_ibr_5.IN3 a_36042_6265# VSS.t356 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1767 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.VOUT CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VDD93.t182 VDD93.t181 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1768 a_32071_11196# CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t48 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1769 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD110.t73 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1770 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN VDD99.t109 VDD99.t108 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1771 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD105.t164 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1772 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 VDD.t35 VDD.t31 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1773 a_45131_n17599# RST.t71 a_44971_n17599# VSS.t2045 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1774 a_29054_11196# CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t56 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1775 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_48422_n2199# VSS.t2465 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1776 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VDD96.t208 VDD96.t207 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1777 a_27529_n18723# CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t281 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1778 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD93.t210 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1779 a_46608_n5176# VDD108.t462 VSS.t520 VSS.t519 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1780 VDD93 VDD93.t90 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VDD93.t91 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1781 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VDD93.t18 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1782 a_37999_280# mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 VSS.t1502 VSS.t24 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1783 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD93.t55 VDD93.t54 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1784 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t15 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT VDD99.t168 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1785 a_23709_810# CLK_div_96_mag_0.JK_FF_mag_5.Q.t9 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_2.OUT VSS.t1065 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1786 VSS CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN VSS.t2285 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X1787 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD105.t350 VDD105.t349 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1788 a_48623_n13424# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 VSS.t1735 VSS.t1734 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1789 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT a_35747_n1822# VSS.t759 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1790 dec3x8_ibr_mag_0.and_3_ibr_2.nand3_mag_ibr_0.OUT dec3x8_ibr_mag_0.and_3_ibr_3.IN1 VDD.t8 VDD.t7 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1791 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD93.t87 VDD93.t89 VDD93.t88 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1792 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 VDD93.t111 VDD93.t110 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1793 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t11 a_46755_574# VSS.t1082 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1794 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD110.t111 VDD110.t110 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1795 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_36588_n15495# VSS.t1860 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1796 VDD96 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_2.OUT CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT VDD96.t89 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1797 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK.t42 VDD105.t469 VDD105.t348 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1798 a_48469_1671# CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT VSS.t2326 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1799 VSS CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN VSS.t1346 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X1800 a_51028_n16724# RST.t72 a_50868_n16724# VSS.t2044 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1801 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD110.t126 VDD110.t125 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1802 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_26770_n16588# VSS.t1524 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1803 a_30727_n17626# CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t329 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1804 a_55310_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t1293 VSS.t1292 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1805 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VDD99.t279 VDD99.t278 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1806 a_36873_n1222# mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 VSS.t576 VSS.t575 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1807 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK.t43 VSS.t2499 VSS.t2498 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1808 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD96.t102 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1809 VSS VDD93.t480 a_23289_n6009# VSS.t260 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1810 VDD96 CLK_div_96_mag_0.JK_FF_mag_4.Q.t7 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_2.OUT VDD96.t340 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1811 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD110.t30 VDD110.t29 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1812 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t8 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 VDD110.t457 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1813 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD90.t388 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1814 a_30589_n2952# CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VSS.t429 VSS.t428 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1815 a_45730_10154# CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t14 a_45570_10154# VSS.t2211 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1816 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD90.t46 VDD90.t45 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1817 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_2x1_ibr_0.I0 a_39124_280# VSS.t1355 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1818 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.t10 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VDD99.t84 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1819 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 VDD108.t135 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1820 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_47252_6240# VSS.t1130 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1821 a_44475_n5176# RST.t73 a_44315_n5176# VSS.t2043 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1822 a_36202_6821# dec3x8_ibr_mag_0.and_3_ibr_6.IN3 a_36042_6821# VSS.t277 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1823 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD108.t274 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1824 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 a_44229_5143# VSS.t2116 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1825 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT VDD108.t316 VDD108.t315 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1826 a_44282_10154# CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t330 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1827 VDD96 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 CLK_div_96_mag_0.JK_FF_mag_4.QB VDD96.t97 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1828 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 VSS.t2352 VSS.t2351 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X1829 a_22424_n1833# CLK_div_96_mag_0.JK_FF_mag_5.Q.t10 a_22264_n1833# VSS.t1066 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1830 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD100.t79 VDD100.t81 VDD100.t80 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1831 a_26266_11196# CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS.t1875 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1832 a_30336_10099# CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t5 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VSS.t743 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1833 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_44888_1671# VSS.t72 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1834 Vdiv110 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 VSS.t1773 VSS.t1772 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X1835 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_47424_n17599# VSS.t871 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1836 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD93.t165 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1837 a_47050_n7372# CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t8 VSS.t498 VSS.t497 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1838 a_44793_5143# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS.t847 VSS.t846 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1839 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 VDD96.t26 VDD96.t25 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1840 a_53126_6240# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K VSS.t61 VSS.t60 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1841 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t2 VDD100.t354 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1842 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.t5 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT VDD108.t214 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1843 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD105.t119 VDD105.t118 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1844 a_50281_n17599# VDD110.t497 VSS.t1014 VSS.t1013 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1845 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_50874_n15583# VSS.t1723 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1846 a_48832_n1102# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VSS.t1496 VSS.t1495 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1847 CLK_div_105_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_105_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VDD105.t196 VDD105.t195 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X1848 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB VDD105.t436 VDD105.t435 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1849 VDD96 VDD96.t155 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_2.OUT VDD96.t156 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1850 a_24922_n17626# CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS.t1816 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1851 VDD93 RST.t74 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT VDD93.t400 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1852 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD93.t51 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1853 a_36873_280# mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 VSS.t622 VSS.t621 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1854 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_54537_n6818# VSS.t1562 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1855 a_22551_n14504# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 VSS.t2338 VSS.t2337 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1856 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD93.t207 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1857 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.t4 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 VDD93.t160 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1858 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD110.t354 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1859 VSS CLK.t44 a_31733_n19822# VSS.t2500 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1860 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT VSS.t724 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1861 RST CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN VSS.t1729 VSS.t1728 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1862 CLK_div_96_mag_0.JK_FF_mag_0.Q CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD96.t86 VDD96.t85 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1863 Vdiv99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT VDD99.t344 VDD99.t343 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1864 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD110.t109 VDD110.t108 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1865 a_50111_n5768# CLK_div_108_new_mag_0.JK_FF_mag_1.CLK a_49951_n5768# VSS.t1748 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1866 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD105.t56 VDD105.t58 VDD105.t57 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1867 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 VDD100.t31 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1868 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.VOUT CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN VDD93.t40 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X1869 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD90.t317 VDD90.t316 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1870 dec3x8_ibr_mag_0.and_3_ibr_6.nand3_mag_ibr_0.OUT F0.t16 a_38454_6265# VSS.t275 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1871 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_44953_5143# VSS.t1454 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1872 VSS CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t4 a_28817_n18723# VSS.t2380 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1873 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t4 VDD99.t463 VDD99.t462 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1874 a_51481_n9064# CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.t5 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT VSS.t2267 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1875 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t0 VDD108.t143 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1876 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD90.t290 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1877 VSS CLK.t45 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VSS.t2503 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1878 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_29871_n1855# VSS.t1828 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1879 a_47036_n15629# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t3 VSS.t2308 VSS.t2307 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1880 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT VDD100.t286 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1881 VDD100 RST.t75 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD100.t372 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1882 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT VSS.t2298 VSS.t2297 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1883 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 VDD108.t332 VDD108.t331 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1884 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t6 VDD108.t183 VDD108.t182 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1885 a_43757_n6273# CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t9 a_43597_n6273# VSS.t493 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1886 a_27150_11196# CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t9 a_26990_11196# VSS.t1240 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1887 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.t2 VDD90.t340 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1888 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 VDD105.t80 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1889 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_105_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 VSS.t607 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X1890 a_50721_n1102# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VSS.t947 VSS.t946 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1891 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB VDD93.t323 VDD93.t322 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1892 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t6 VDD90.t231 VDD90.t230 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1893 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.IN2 VDD.t147 VDD.t112 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1894 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD99.t91 VDD99.t90 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1895 a_48023_10154# RST.t76 a_47863_10154# VSS.t2042 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1896 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 a_37999_n1222# VSS.t1345 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1897 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t4 a_39126_n8931# VSS.t747 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1898 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT a_47187_2768# VSS.t115 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1899 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD99.t64 VDD99.t63 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1900 a_33429_n15491# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 VSS.t1334 VSS.t1333 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1901 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.t5 VSS.t124 VSS.t123 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X1902 VDD108 CLK.t46 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 VDD108.t446 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1903 a_44885_n6273# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t462 VSS.t146 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1904 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_3.Q VDD96.t57 VDD96.t56 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1905 VSS CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.CLK VSS.t1730 nfet_03v3 ad=86.8f pd=0.92u as=86.8f ps=0.92u w=0.22u l=0.28u
X1906 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT RST.t77 VDD96.t287 VDD96.t286 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1907 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD110.t233 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1908 CLK_div_108_new_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.t7 VDD108.t112 VDD108.t111 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1909 a_47751_2768# CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT VSS.t1719 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1910 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 a_44117_n2243# VSS.t2458 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1911 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 VDD110.t418 VDD110.t417 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1912 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_51438_n15583# VSS.t1781 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1913 a_23025_6159# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS.t976 VSS.t975 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1914 VDD F1.t13 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 VDD.t104 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1915 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_54182_n17599# VSS.t1935 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1916 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 a_32455_n16632# VSS.t2099 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1917 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 VDD90.t32 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1918 a_54004_5143# RST.t78 a_53844_5143# VSS.t2041 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1919 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD110.t35 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1920 VDD90 CLK.t47 CLK_div_90_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN VDD90.t454 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1921 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD90.t418 VDD90.t417 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1922 dec3x8_ibr_mag_0.and_3_ibr_2.nand3_mag_ibr_0.OUT dec3x8_ibr_mag_0.and_3_ibr_3.IN1 a_38454_6821# VSS.t275 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1923 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD99.t293 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1924 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VDD90.t123 VDD90.t122 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1925 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K VDD110.t246 VDD110.t245 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1926 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.t8 a_45235_n9063# VSS.t504 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1927 VSS CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 a_24337_n6010# VSS.t669 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1928 a_52139_n18696# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VSS.t834 VSS.t833 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1929 VDD93 RST.t79 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD93.t397 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1930 a_25482_n16632# CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t16 a_25322_n16632# VSS.t1171 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1931 a_53469_n15631# CLK.t48 a_53309_n15631# VSS.t2506 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1932 a_28737_n2996# CLK_div_96_mag_0.JK_FF_mag_2.Q a_28577_n2996# VSS.t2156 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1933 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t10 VSS.t500 VSS.t499 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1934 a_26636_n8734# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t41 VSS.t40 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1935 a_29214_n6271# CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 VSS.t1666 VSS.t1665 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1936 VDD110 CLK.t49 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT VDD110.t472 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1937 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.t6 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD90.t445 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1938 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN VDD93.t2 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X1939 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_44511_n9019# VSS.t1485 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1940 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT VDD99.t17 VDD99.t16 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1941 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT VDD105.t299 VDD105.t298 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1942 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_30187_6159# VSS.t238 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1943 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_96_mag_0.JK_FF_mag_2.Q VDD96.t320 VDD96.t319 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1944 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.t6 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD93.t34 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1945 a_44888_1671# CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t19 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1946 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VDD90.t376 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1947 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_47704_n1102# VSS.t156 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1948 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.JK_FF_mag_1.Q VDD108.t417 VDD108.t416 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1949 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_2.OUT Vdiv108.t6 VDD108.t213 VDD108.t212 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1950 a_45343_n16680# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT VSS.t836 VSS.t835 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1951 a_26343_n7107# CLK.t50 a_26183_n7107# VSS.t2507 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1952 a_25625_n6010# RST.t80 a_25465_n6010# VSS.t2040 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1953 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS.t2552 VSS.t2551 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1954 a_52951_7381# CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 VSS.t2115 VSS.t2114 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1955 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB VDD100.t318 VDD100.t317 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1956 CLK_div_100_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_100_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS.t459 VSS.t458 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X1957 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD100.t267 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1958 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t5 a_25420_n13385# VDD99.t176 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X1959 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 a_52652_n10117# VSS.t1024 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1960 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT a_28580_n8735# VSS.t1566 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1961 VDD105 dec3x8_ibr_mag_0.and_3_ibr_6.nand3_mag_ibr_0.OUT VDD.t37 VDD.t36 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1962 VSS CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_23794_n17626# VSS.t244 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1963 a_44413_n18696# CLK_div_110_mag_0.CLK_div_10_mag_0.CLK a_44253_n18696# VSS.t542 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1964 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t11 VDD105.t241 VDD105.t240 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1965 a_48534_5187# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VSS.t68 VSS.t67 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1966 a_29834_n699# CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS.t1297 VSS.t1296 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1967 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K VDD110.t242 VDD110.t241 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1968 a_29772_10099# CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t1438 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1969 a_54781_10154# CLK_div_105_mag_0.CLK_div_10_mag_1.CLK a_54621_10154# VSS.t1560 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1970 a_30244_398# CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t1332 VSS.t1331 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1971 a_35747_n1222# mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.IN2 VSS.t2021 VSS.t1343 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1972 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_47902_n6273# VSS.t146 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1973 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t6 VDD90.t168 VDD90.t167 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1974 CLK_div_105_mag_0.CLK_div_10_mag_1.CLK CLK_div_105_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 VSS.t431 VSS.t430 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X1975 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD108.t20 VDD108.t22 VDD108.t21 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1976 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD90.t249 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1977 a_34736_n15539# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K VSS.t2167 VSS.t2166 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1978 VSS CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_2.OUT a_26256_3016# VSS.t823 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1979 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t0 VDD90.t373 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1980 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t12 VDD99.t135 VDD99.t134 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1981 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 VDD100.t193 VDD100.t192 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1982 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD96.t273 VDD96.t272 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1983 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK.t51 VSS.t2509 VSS.t2508 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1984 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD90.t353 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1985 VSS CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t12 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 VSS.t1001 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X1986 a_26663_398# CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t175 VSS.t174 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1987 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD96.t1 VDD96.t0 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1988 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT VDD110.t84 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1989 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD90.t308 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1990 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_47858_n2243# VSS.t843 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X1991 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t12 VDD105.t243 VDD105.t242 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X1992 a_26820_3016# CLK_div_96_mag_0.JK_FF_mag_4.Q.t8 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_2.OUT VSS.t2284 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X1993 a_54592_n18696# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t1934 VSS.t109 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X1994 a_45612_1671# CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t15 a_45452_1671# VSS.t1158 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1995 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD110.t296 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1996 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t13 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD93.t285 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1997 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 VDD110.t46 VDD110.t45 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1998 a_28623_n15537# CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t17 a_28463_n15537# VSS.t1248 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1999 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD108.t17 VDD108.t19 VDD108.t18 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2000 VDD99 VDD99.t44 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VDD99.t45 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2001 a_52806_n9020# CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.t1 VSS.t644 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2002 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 VDD110.t44 VDD110.t43 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2003 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN VSS.t2246 VSS.t2245 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2004 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t11 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD93.t458 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2005 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t0 VDD90.t380 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2006 VSS CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 a_24968_3016# VSS.t955 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2007 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t14 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 VSS.t2277 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2008 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.t0 VDD99.t65 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2009 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD93.t69 VDD93.t68 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2010 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS.t142 VSS.t141 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2011 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 VDD100.t172 VDD100.t171 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2012 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD99.t322 VDD99.t321 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2013 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.IN2 VDD108.t158 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2014 a_31661_10099# CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.t1 VSS.t1669 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2015 a_47187_2768# CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 VSS.t942 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2016 VDD108 RST.t81 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD108.t349 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2017 a_25532_3016# CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 VSS.t335 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2018 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 VDD105.t224 VDD105.t223 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2019 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 a_36742_n16592# VSS.t1581 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2020 a_44324_1671# CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t427 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2021 a_53934_n9020# CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t660 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2022 a_46964_n9019# CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t362 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2023 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t5 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD90.t400 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2024 VDD F0.t17 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_1.IN2 VDD.t176 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2025 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT VDD110.t290 VDD110.t289 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2026 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD108.t257 VDD108.t256 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2027 Vdiv90 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 VSS.t1810 VSS.t1809 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X2028 VSS VDD96.t384 a_26980_3016# VSS.t1459 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2029 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT a_53216_n10117# VSS.t657 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2030 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t5 a_46774_n6273# VSS.t493 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2031 a_30881_n18723# CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t328 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2032 VSS CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_24358_n17626# VSS.t987 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2033 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD90.t12 VDD90.t11 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2034 VDD90 RST.t82 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD90.t203 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2035 CLK_div_108_new_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t11 VDD108.t97 VDD108.t96 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2036 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT RST.t83 VDD108.t348 VDD108.t347 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2037 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t6 VDD96.t332 VDD96.t331 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2038 CLK_div_90_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.t8 VDD90.t175 VDD90.t174 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2039 VDD100 RST.t84 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD100.t369 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2040 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_26226_n9831# VSS.t456 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2041 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_25508_n8734# VSS.t1926 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2042 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t0 VDD99.t13 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2043 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD110.t144 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2044 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 a_49098_5187# VSS.t682 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2045 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD93.t141 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2046 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD96.t244 VDD96.t243 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2047 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT RST.t85 VDD96.t285 VDD96.t284 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2048 VSS CLK_div_96_mag_0.JK_FF_mag_4.Q.t9 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 VSS.t1217 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2049 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.IN1 a_32750_n7675# VDD93.t381 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X2050 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VDD90.t323 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2051 dec3x8_ibr_mag_0.and_3_ibr_7.nand3_mag_ibr_0.OUT F2.t5 VDD.t77 VDD.t76 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2052 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD96.t152 VDD96.t154 VDD96.t153 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2053 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD110.t261 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2054 a_52811_1671# CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t0 VSS.t984 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2055 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN VDD99.t19 VDD99.t18 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2056 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK.t52 VDD110.t476 VDD110.t475 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2057 a_30187_6159# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VSS.t301 VSS.t300 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2058 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_50875_n2243# VSS.t434 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2059 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t18 VDD99.t178 VDD99.t177 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2060 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD90.t333 VDD90.t332 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2061 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_44061_n15627# VSS.t963 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2062 a_55156_n18696# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t1937 VSS.t109 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2063 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_23025_6159# VSS.t794 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2064 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD90.t411 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2065 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN VSS.t805 VSS.t767 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X2066 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_54004_5143# VSS.t1834 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2067 a_33812_n13270# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT a_33652_n13270# VDD99.t37 pfet_03v3 ad=0.624p pd=2.92u as=0.624p ps=2.92u w=2.4u l=0.28u
X2068 a_23145_810# RST.t86 a_22985_810# VSS.t2039 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2069 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_54383_n5721# VSS.t1561 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2070 VSS VDD100.t487 a_54663_1671# VSS.t2407 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2071 a_25856_10099# CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t112 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2072 a_30760_n20290# CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.t6 CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN VDD99.t120 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X2073 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_47196_n15629# VSS.t2191 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2074 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN VDD99.t244 VDD99.t243 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2075 a_22460_n9884# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS.t192 VSS.t191 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2076 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN VDD93.t430 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X2077 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t12 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD108.t98 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2078 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.CLK VSS.t94 VSS.t93 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2079 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 a_42521_n13474# VDD110.t168 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X2080 VDD96 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD96.t261 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2081 CLK_div_105_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_105_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS.t863 VSS.t862 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X2082 a_44055_n16724# CLK.t53 a_43895_n16724# VSS.t1376 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2083 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_41124_n16098# VSS.t556 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2084 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD99.t208 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2085 a_26256_3016# RST.t87 a_26096_3016# VSS.t2038 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2086 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 VDD105.t153 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2087 VSS CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_29778_11196# VSS.t590 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2088 VSS CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_26811_n17626# VSS.t1404 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2089 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD105.t423 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2090 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD110.t313 VDD110.t312 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2091 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD90.t434 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2092 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_29213_5018# VSS.t196 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2093 a_43751_n5176# CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t13 a_43591_n5176# VSS.t501 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2094 a_51957_n6821# CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t1389 VSS.t1388 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2095 a_26984_10099# CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS.t1178 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2096 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_3.Q VSS.t437 VSS.t436 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2097 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 a_52951_7381# VSS.t2012 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2098 VDD96 RST.t88 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VDD96.t280 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2099 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 VDD110.t208 VDD110.t207 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2100 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT VDD108.t320 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2101 a_28490_11196# CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.t7 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K VSS.t1078 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2102 VSS CLK.t54 a_30060_9000# VSS.t758 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2103 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_53375_1671# VSS.t599 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2104 CLK_div_100_mag_0.CLK_div_10_mag_1.CLK CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 VSS.t1832 VSS.t1831 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X2105 VDD99 CLK.t55 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VDD99.t502 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2106 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t7 a_53464_n18696# VSS.t689 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2107 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT VDD105.t101 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2108 VDD96 RST.t89 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD96.t278 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2109 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD108.t80 VDD108.t79 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2110 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t5 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VDD100.t129 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2111 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN VSS.t2253 VSS.t2252 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2112 a_25502_n9875# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS.t1307 VSS.t1306 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2113 a_24784_n8778# VDD93.t481 VSS.t259 VSS.t258 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2114 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD90.t193 VDD90.t192 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2115 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_90_mag_0.CLK_div_10_mag_0.CLK VDD90.t103 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2116 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD96.t139 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2117 VDD93 RST.t90 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD93.t394 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2118 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 VDD.t53 VDD.t52 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2119 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VDD108.t73 VDD108.t72 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2120 a_48620_n5176# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t736 VSS.t735 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2121 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD90.t438 VDD90.t437 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2122 VDD110 RST.t91 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD110.t398 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2123 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t12 VSS.t2450 VSS.t2449 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2124 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD90.t287 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2125 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_54456_n2199# VSS.t98 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2126 VSS CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_28093_n18723# VSS.t932 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2127 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 VDD93.t386 VDD93.t385 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2128 a_48017_9057# CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 VSS.t1545 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2129 a_25644_n2996# CLK_div_96_mag_0.JK_FF_mag_0.Q a_25484_n2996# VSS.t1693 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2130 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 VDD90.t352 VDD90.t351 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2131 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K VSS.t1677 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2132 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 VDD99.t105 VDD99.t104 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2133 a_39120_n10028# CLK_div_93_mag_0.CLK_div_3_mag_0.CLK a_38960_n10028# VSS.t697 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2134 a_53249_n6862# CLK_div_108_new_mag_0.JK_FF_mag_1.Q a_53089_n6862# VSS.t2312 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2135 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_44235_6240# VSS.t2121 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2136 VSS VDD99.t515 a_25806_n17626# VSS.t2432 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2137 VDD99 RST.t92 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT VDD99.t362 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2138 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_26616_n15491# VSS.t1523 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2139 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN VSS.t392 VSS.t391 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2140 Vdiv90 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 a_33405_7558# VDD90.t379 pfet_03v3 ad=1.06p pd=5.68u as=0.624p ps=2.92u w=2.4u l=0.28u
X2141 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 VDD100.t345 VDD100.t344 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2142 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t13 a_31128_n7028# VSS.t1507 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2143 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD93.t130 VDD93.t129 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2144 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 VDD93.t132 VDD93.t131 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2145 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_47816_6284# VSS.t66 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2146 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK.t56 VDD110.t478 VDD110.t477 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2147 a_25292_10099# CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.t1 VSS.t112 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2148 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VDD100.t263 VDD100.t262 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2149 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K VDD99.t23 VDD99.t22 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2150 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_45006_10154# VSS.t887 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2151 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_44687_n1102# VSS.t1520 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2152 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD90.t183 VDD90.t182 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2153 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 VDD93.t10 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2154 dec3x8_ibr_mag_0.and_3_ibr_3.nand3_mag_ibr_0.OUT F2.t6 VDD.t79 VDD.t78 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2155 a_50109_6240# VDD105.t485 VSS.t1103 VSS.t1102 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2156 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_39844_n10028# VSS.t157 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2157 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t14 VDD108.t102 VDD108.t101 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2158 a_23409_11196# RST.t93 a_23249_11196# VSS.t2037 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2159 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD100.t208 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2160 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD110.t194 VDD110.t193 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2161 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN VDD93.t21 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X2162 a_51205_n7921# CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.t6 CLK_div_108_new_mag_0.CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN VSS.t1189 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2163 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t16 VDD100.t404 VDD100.t403 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2164 a_31451_n17626# RST.t94 a_31291_n17626# VSS.t2036 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2165 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t13 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 VDD105.t244 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2166 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 a_29241_7256# VSS.t1335 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2167 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT RST.t95 VDD99.t361 VDD99.t360 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2168 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT VSS.t1920 VSS.t1919 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2169 VSS CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT a_22559_n7106# VSS.t720 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2170 VSS CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_21841_n6009# VSS.t906 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2171 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD96.t84 VDD96.t83 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2172 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t5 VDD99.t465 VDD99.t464 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2173 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 VSS.t9 VSS.t8 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X2174 a_26099_398# CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS.t355 VSS.t354 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2175 VDD96 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD96.t235 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2176 a_51393_n6821# CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS.t1391 VSS.t1390 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2177 a_50675_n5724# CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS.t982 VSS.t981 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2178 VSS CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_32795_11196# VSS.t958 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2179 a_43606_2768# CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K VSS.t1909 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2180 VSS CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t13 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VSS.t1124 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2181 a_44619_n16724# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT VSS.t571 VSS.t570 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2182 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD93.t330 VDD93.t329 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2183 a_32175_n17626# CLK.t57 a_32015_n17626# VSS.t2512 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2184 VDD F1.t14 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 VDD.t107 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2185 a_55315_n16684# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 VSS.t827 VSS.t826 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2186 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN VDD93.t5 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X2187 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD100.t308 VDD100.t307 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2188 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VDD96.t149 VDD96.t151 VDD96.t150 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2189 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD100.t63 VDD100.t62 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2190 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD96.t5 VDD96.t4 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2191 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD108.t393 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2192 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.t6 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT VDD108.t404 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2193 a_50316_10154# CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 VSS.t612 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2194 a_48741_9057# CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t14 a_48581_9057# VSS.t1228 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2195 a_48268_n1102# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VSS.t842 VSS.t841 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2196 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_34896_n15539# VSS.t1859 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2197 a_46246_n10116# CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.t9 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB VSS.t507 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2198 a_30164_n7017# CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 VSS.t315 VSS.t314 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2199 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_54028_n18696# VSS.t109 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2200 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.t7 VDD93.t33 VDD93.t32 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2201 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t5 VDD93.t243 VDD93.t242 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2202 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK VDD93.t206 VDD93.t205 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2203 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t7 CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 VDD100.t251 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2204 CLK_div_105_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT VDD105.t319 VDD105.t318 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X2205 a_25318_6115# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t7 VSS.t1161 VSS.t1160 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2206 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD90.t195 VDD90.t194 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2207 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VDD100.t3 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2208 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t17 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VDD100.t405 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2209 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 VDD110.t143 VDD110.t142 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2210 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t14 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD93.t455 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2211 a_33019_n16588# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT VSS.t2103 VSS.t2102 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2212 a_45618_2768# CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t18 a_45458_2768# VSS.t2200 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2213 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD93.t197 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2214 a_53973_n6862# RST.t96 a_53813_n6862# VSS.t2035 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2215 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_26817_n699# VSS.t1052 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2216 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 VDD110.t173 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2217 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VDD108.t167 VDD108.t166 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2218 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_45517_5187# VSS.t812 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2219 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN VSS.t716 VSS.t715 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2220 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD110.t15 VDD110.t17 VDD110.t16 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2221 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_44517_n10160# VSS.t119 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2222 a_54663_1671# CLK_div_100_mag_0.CLK_div_10_mag_1.CLK a_54503_1671# VSS.t2001 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2223 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD99.t59 VDD99.t58 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2224 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD100.t322 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2225 a_44971_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS.t376 VSS.t375 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2226 VDD90 VDD90.t59 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VDD90.t60 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2227 a_46105_n18696# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t1352 VSS.t1351 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2228 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.t0 VDD90.t269 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2229 a_47453_9057# CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 VSS.t1138 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2230 CLK_div_108_new_mag_0.JK_FF_mag_0.QB Vdiv108.t7 a_55101_n6818# VSS.t1185 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2231 a_34890_n16636# CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t19 a_34730_n16636# VSS.t1249 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2232 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD100.t158 VDD100.t157 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2233 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.t6 VDD99.t456 VDD99.t455 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2234 a_44625_n15583# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT VSS.t968 VSS.t967 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2235 a_50829_n6865# RST.t97 a_50669_n6865# VSS.t2034 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2236 VDD110 CLK.t58 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT VDD110.t479 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2237 VDD105 VDD105.t52 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT VDD105.t53 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2238 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD90.t56 VDD90.t58 VDD90.t57 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2239 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD110.t124 VDD110.t123 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2240 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD93.t138 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2241 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD105.t49 VDD105.t51 VDD105.t50 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2242 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_29307_n1855# VSS.t1613 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2243 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_44170_2768# VSS.t16 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2244 VDD mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT Vdiv.t1 VDD.t123 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2245 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD93.t157 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2246 VSS CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 a_30317_n18723# VSS.t1563 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2247 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB VDD100.t393 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2248 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_22988_n1789# VSS.t1739 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2249 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 VDD100.t444 VDD100.t443 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2250 VSS CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_33744_n17626# VSS.t1927 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2251 a_30060_9000# CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.t9 CLK_div_90_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN VSS.t758 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2252 a_53375_1671# CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t2005 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2253 VSS VDD105.t487 a_48747_10154# VSS.t1104 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2254 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK.t59 VDD110.t483 VDD110.t482 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2255 a_43947_n9019# CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t351 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2256 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 VDD90.t135 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2257 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB VDD108.t184 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2258 VSS CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_21995_n7106# VSS.t720 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2259 a_47760_n15585# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT VSS.t1710 VSS.t1709 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2260 a_37999_880# mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 VSS.t25 VSS.t24 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2261 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t6 VDD108.t228 VDD108.t227 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2262 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT a_47299_10154# VSS.t1542 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2263 a_44734_2768# CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VSS.t1849 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2264 VDD90 dec3x8_ibr_mag_0.and_3_ibr_0.nand3_mag_ibr_0.OUT VSS.t386 VSS.t99 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2265 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT VDD99.t25 VDD99.t24 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2266 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.t10 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VDD108.t113 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2267 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 VDD93.t46 VDD93.t45 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2268 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 VDD90.t206 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2269 a_39420_6265# F2.t7 VSS.t1204 VSS.t1203 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2270 a_23139_n287# CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.IN1 VSS.t1756 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2271 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD105.t342 VDD105.t341 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2272 a_22418_n2930# CLK_div_96_mag_0.JK_FF_mag_5.Q.t11 a_22258_n2930# VSS.t1067 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2273 a_25702_11196# CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t393 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2274 VDD100 VDD100.t75 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VDD100.t76 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2275 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD100.t273 VDD100.t272 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2276 VDD93 VDD93.t83 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD93.t84 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2277 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VDD93.t319 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2278 a_48092_n9063# CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VSS.t737 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2279 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t14 VDD99.t137 VDD99.t136 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2280 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT VDD99.t315 VDD99.t314 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2281 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VDD105.t25 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2282 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB a_29708_n8735# VSS.t203 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2283 VDD105 dec3x8_ibr_mag_0.and_3_ibr_6.nand3_mag_ibr_0.OUT VSS.t649 VSS.t648 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2284 CLK_div_100_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT VSS.t867 VSS.t866 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X2285 a_51285_n1102# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VSS.t433 VSS.t432 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2286 Vdiv93 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS.t1373 VSS.t1372 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2287 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_52657_2768# VSS.t2146 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2288 a_48148_n17599# RST.t98 a_47988_n17599# VSS.t2033 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2289 a_23948_n18723# CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t5 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.t2 VSS.t2383 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2290 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT RST.t99 VDD105.t391 VDD105.t390 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2291 a_36873_n1822# mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 VSS.t1778 VSS.t575 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2292 CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t6 a_54978_6284# VSS.t859 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2293 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 a_29801_1733# VDD96.t313 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X2294 a_47338_n6273# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS.t2083 VSS.t146 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2295 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD105.t465 VDD105.t464 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2296 VSS CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT Vdiv90.t3 VSS.t2177 nfet_03v3 ad=86.8f pd=0.92u as=86.8f ps=0.92u w=0.22u l=0.28u
X2297 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 VSS.t1580 VSS.t1579 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X2298 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS.t8 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X2299 VSS CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_24512_n18723# VSS.t1813 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2300 Vdiv mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT a_39124_880# VSS.t1355 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2301 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD90.t211 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2302 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD110.t369 VDD110.t368 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2303 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 a_23948_n13382# VDD99.t292 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X2304 VDD mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.OUT VDD.t54 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2305 a_31506_5018# CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 a_31346_5018# VSS.t1626 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2306 VSS VDD100.t489 a_54669_2768# VSS.t2410 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2307 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VDD100.t341 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2308 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD96.t275 VDD96.t274 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2309 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT a_50917_n9020# VSS.t1492 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2310 VSS VDD93.t483 a_26349_n6010# VSS.t255 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2311 CLK_div_108_new_mag_0.JK_FF_mag_1.Q CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD108.t241 VDD108.t240 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2312 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT a_48017_9057# VSS.t774 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2313 a_51729_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VSS.t1574 VSS.t1573 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2314 a_54658_n9064# CLK.t60 a_54498_n9064# VSS.t2513 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2315 VSS CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_24901_n6010# VSS.t292 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2316 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t10 VDD105.t98 VDD105.t97 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2317 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.CLK CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VSS.t1557 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2318 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT RST.t100 VDD100.t368 VDD100.t367 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2319 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD110.t134 VDD110.t133 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2320 a_45189_n15583# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t479 VSS.t478 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2321 a_47140_n1146# CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 a_46980_n1146# VSS.t2457 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2322 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT RST.t101 VDD90.t444 VDD90.t443 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2323 a_39420_6821# F2.t8 VSS.t1205 VSS.t1203 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2324 a_28583_n1899# VDD96.t385 VSS.t1458 VSS.t1457 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2325 a_29301_n2996# CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VSS.t761 VSS.t760 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2326 a_28617_n16634# CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t20 a_28457_n16634# VSS.t1250 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2327 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD90.t27 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2328 VSS VDD105.t488 a_51764_10154# VSS.t1107 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2329 a_48581_9057# CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT VSS.t568 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2330 a_51015_7381# CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 VSS.t681 VSS.t680 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2331 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 F0.t18 VSS.t2446 VSS.t2445 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2332 a_34468_n17626# RST.t102 a_34308_n17626# VSS.t2032 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2333 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t6 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VDD99.t471 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2334 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD100.t152 VDD100.t151 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2335 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.t0 VDD108.t76 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2336 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD90.t348 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2337 VDD110 CLK.t61 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT VDD110.t484 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2338 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 VDD108.t129 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2339 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 VDD100.t11 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2340 CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD100.t402 VDD100.t401 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2341 a_27856_n8779# VDD93.t484 VSS.t254 VSS.t253 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2342 a_40375_n7552# CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 VDD93.t247 VDD93.t246 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X2343 a_36873_880# mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 VSS.t1791 VSS.t621 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2344 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VDD100.t114 VDD100.t113 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2345 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT Vdiv100.t4 a_35747_280# VSS.t1276 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2346 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_53738_n1102# VSS.t231 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2347 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t15 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD108.t103 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2348 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t15 a_47723_574# VSS.t1082 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2349 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD100.t36 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2350 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t6 a_31737_n15535# VSS.t1193 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2351 a_45458_2768# CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VSS.t1908 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2352 VDD96 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT VDD96.t264 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2353 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 a_37999_280# VSS.t15 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2354 a_49997_n1146# VDD100.t490 VSS.t2414 VSS.t2413 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2355 a_27342_n1855# CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VSS.t2155 VSS.t2154 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2356 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 VDD110.t42 VDD110.t41 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2357 CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.t7 VSS.t2272 VSS.t2271 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X2358 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t15 VDD105.t459 VDD105.t458 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2359 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB VDD100.t205 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2360 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 a_29144_n8735# VSS.t2131 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2361 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VDD100.t200 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2362 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD110.t70 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2363 a_22551_n16006# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 VSS.t2336 VSS.t2335 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2364 a_53945_2768# RST.t103 a_53785_2768# VSS.t2031 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2365 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_30315_n15493# VSS.t2349 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2366 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t21 VSS.t1252 VSS.t1251 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2367 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD99.t3 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2368 a_23030_n8743# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t710 VSS.t709 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2369 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t6 VDD90.t399 VDD90.t398 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2370 a_53298_n17599# VDD110.t498 VSS.t1016 VSS.t1015 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2371 a_31571_n16632# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K VSS.t2126 VSS.t2125 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2372 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t22 VDD99.t180 VDD99.t179 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2373 a_32230_5018# RST.t104 a_32070_5018# VSS.t473 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2374 VDD108 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD108.t307 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2375 a_35460_n15495# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT VSS.t2171 VSS.t2170 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2376 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD108.t147 VDD108.t146 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2377 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB VDD90.t295 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2378 a_25375_354# CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t7 VSS.t2204 VSS.t2203 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2379 a_51647_n10161# CLK.t62 a_51487_n10161# VSS.t2514 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2380 a_27939_n17626# CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS.t938 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2381 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t4 VDD110.t446 VDD110.t445 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2382 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 a_45969_n2199# VSS.t2456 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2383 VDD90 VDD90.t52 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD90.t53 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2384 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t7 VDD99.t470 VDD99.t469 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2385 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VDD105.t185 VDD105.t184 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2386 a_44170_2768# CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t426 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2387 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VDD90.t368 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2388 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VDD99.t281 VDD99.t280 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2389 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t19 VDD100.t409 VDD100.t408 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2390 VSS CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 a_24491_n7107# VSS.t1711 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2391 a_22985_810# CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT VSS.t1869 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2392 a_28663_n17626# CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.t7 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS.t2359 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2393 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 F0.t19 VDD.t180 VDD.t179 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2394 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t10 CLK_div_90_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD90.t259 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2395 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 F1.t15 VSS.t1214 VSS.t1213 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2396 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 VSS.t870 VSS.t869 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2397 CLK_div_96_mag_0.JK_FF_mag_2.QB CLK_div_96_mag_0.JK_FF_mag_2.Q a_27496_n2952# VSS.t1697 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2398 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD99.t379 VDD99.t378 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2399 a_48986_n2199# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VSS.t632 VSS.t631 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2400 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD110.t367 VDD110.t366 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2401 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t13 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 VDD93.t279 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2402 VSS CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS.t1985 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X2403 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 a_43831_7266# VDD105.t286 pfet_03v3 ad=1.06p pd=5.68u as=0.624p ps=2.92u w=2.4u l=0.28u
X2404 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT Vdiv108.t8 a_36873_280# VSS.t1186 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2405 mux_8x1_ibr_0.mux_2x1_ibr_0.I0 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.OUT a_37999_n1822# VSS.t1345 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2406 VSS CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t11 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VSS.t1241 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2407 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 VDD90.t433 VDD90.t432 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2408 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS.t1637 VSS.t1636 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2409 a_53303_n16728# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K VSS.t1681 VSS.t1680 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2410 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 VDD105.t295 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2411 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.CLK VDD100.t358 VDD100.t357 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2412 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD110.t268 VDD110.t267 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2413 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN VSS.t85 VSS.t84 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X2414 a_53370_n9020# CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t1353 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2415 VSS CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t7 a_33513_10099# VSS.t744 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2416 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD100.t120 VDD100.t119 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2417 a_52657_2768# CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t20 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB VSS.t2435 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2418 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 F1.t16 VDD.t111 VDD.t110 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2419 a_21736_n9884# VDD93.t485 VSS.t252 VSS.t251 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2420 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT VDD105.t289 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2421 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB VDD105.t176 VDD105.t175 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2422 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 VDD99.t101 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2423 VDD108 CLK.t63 CLK_div_108_new_mag_0.CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN VDD108.t449 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2424 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_52385_n13362# VDD110.t89 pfet_03v3 ad=1.06p pd=5.68u as=0.624p ps=2.92u w=2.4u l=0.28u
X2425 VSS CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT VSS.t377 nfet_03v3 ad=86.8f pd=0.92u as=86.8f ps=0.92u w=0.22u l=0.28u
X2426 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD100.t52 VDD100.t51 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2427 a_53014_n1146# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K VSS.t849 VSS.t848 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2428 a_53732_n2243# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS.t945 VSS.t944 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2429 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VDD99.t277 VDD99.t276 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2430 CLK_div_93_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 a_39402_n7788# VSS.t284 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2431 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_96_mag_0.JK_FF_mag_0.QB VDD96.t37 VDD96.t36 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2432 VSS CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t7 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN VSS.t1194 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X2433 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD105.t335 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2434 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 VDD100.t259 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2435 a_47246_5143# CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 a_47086_5143# VSS.t2113 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2436 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_44407_n17599# VSS.t1321 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2437 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD105.t163 VDD105.t162 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2438 VSS CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_31445_n18723# VSS.t2195 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2439 a_54669_2768# CLK_div_100_mag_0.CLK_div_10_mag_1.CLK a_54509_2768# VSS.t2000 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2440 VDD96 CLK_div_96_mag_0.JK_FF_mag_2.Q CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD96.t316 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2441 VSS CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_25082_n17626# VSS.t675 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2442 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD108.t6 VDD108.t5 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2443 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN VDD110.t172 VDD110.t171 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X2444 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.t7 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VDD108.t369 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2445 VDD105 VDD105.t45 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VDD105.t46 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2446 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB VDD93.t389 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2447 VDD100 dec3x8_ibr_mag_0.and_3_ibr_2.nand3_mag_ibr_0.OUT VDD.t60 VDD.t59 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2448 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD105.t10 VDD105.t9 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2449 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VDD100.t138 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2450 CLK_div_96_mag_0.JK_FF_mag_0.QB CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD96.t216 VDD96.t215 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2451 a_47374_n10160# CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VSS.t1291 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2452 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t15 a_28268_n6266# VSS.t998 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2453 VSS CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_22839_10099# VSS.t112 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2454 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT VDD105.t262 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2455 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VDD99.t193 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2456 a_29187_n15493# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT VSS.t2322 VSS.t2321 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2457 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 a_22544_n13819# VSS.t1977 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2458 VDD90 CLK.t64 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VDD90.t457 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2459 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VDD105.t420 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2460 a_27324_5062# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VSS.t133 VSS.t132 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2461 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT VSS.t1767 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2462 VDD96 CLK_div_96_mag_0.JK_FF_mag_4.Q.t10 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 VDD96.t123 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2463 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_26214_n1855# VSS.t2141 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2464 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_26932_n2952# VSS.t1697 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2465 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VDD105.t159 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2466 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS.t2176 VSS.t2175 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2467 a_48422_n2199# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VSS.t155 VSS.t154 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2468 VDD105 CLK.t65 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD105.t470 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2469 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN VSS.t900 VSS.t899 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2470 a_52003_n2199# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VSS.t167 VSS.t166 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2471 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_53221_2768# VSS.t1265 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2472 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD110.t377 VDD110.t376 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2473 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t6 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT VDD100.t132 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2474 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K VDD99.t398 VDD99.t397 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2475 a_35943_n10028# VDD93.t486 VSS.t250 VSS.t249 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2476 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_41117_n13911# VSS.t555 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2477 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t6 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VDD105.t215 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2478 a_35747_n1822# mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_1.IN2 VSS.t1344 VSS.t1343 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2479 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_44436_9057# VSS.t321 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2480 a_53785_2768# CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VSS.t598 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2481 CLK_div_105_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT VSS.t1598 VSS.t1597 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X2482 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD99.t320 VDD99.t319 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2483 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 a_43826_n7684# VDD108.t57 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X2484 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VDD100.t234 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2485 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t8 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 VDD90.t232 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2486 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB VDD105.t417 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2487 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT VDD96.t252 VDD96.t251 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2488 a_32070_5018# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS.t773 VSS.t473 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2489 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 VDD110.t321 VDD110.t320 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2490 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT VSS.t1498 VSS.t1497 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2491 a_47430_n18696# CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_47270_n18696# VSS.t1320 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2492 a_54027_n16728# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT VSS.t1685 VSS.t1684 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2493 a_45000_9057# CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t2328 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2494 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 VDD90.t8 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2495 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 a_51015_7381# VSS.t2011 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2496 Vdiv110 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 VSS.t2107 VSS.t2106 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X2497 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VDD108.t277 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2498 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 VDD100.t186 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2499 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD99.t111 VDD99.t110 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2500 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD100.t61 VDD100.t60 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2501 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_96_mag_0.JK_FF_mag_2.QB a_25650_n1899# VSS.t2332 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2502 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_26368_n2996# VSS.t2145 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2503 VSS CLK.t66 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 VSS.t2515 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2504 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_44799_6284# VSS.t789 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2505 VDD96 CLK.t67 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 VDD96.t357 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2506 a_50310_n15627# CLK.t68 a_50150_n15627# VSS.t2518 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2507 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD110.t167 VDD110.t166 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2508 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 VDD108.t243 VDD108.t242 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2509 a_44315_n5176# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS.t822 VSS.t821 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2510 a_48056_n5176# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS.t1506 VSS.t1505 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2511 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD108.t359 VDD108.t358 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2512 VSS CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_90_mag_0.CLK_div_10_mag_0.CLK VSS.t316 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2513 CLK_div_90_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.t8 VDD90.t241 VDD90.t240 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2514 a_32169_n18723# CLK.t69 a_32009_n18723# VSS.t2519 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2515 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t8 VDD110.t192 VDD110.t191 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2516 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT VDD100.t400 VDD100.t399 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2517 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD110.t277 VDD110.t276 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2518 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_53945_2768# VSS.t1144 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2519 a_47914_n16726# RST.t105 a_47754_n16726# VSS.t2030 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2520 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t11 VDD105.t100 VDD105.t99 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2521 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD93.t25 VDD93.t24 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2522 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD105.t203 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2523 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD93.t57 VDD93.t56 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2524 VSS CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_22275_10099# VSS.t112 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2525 a_51011_n18696# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VSS.t414 VSS.t413 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2526 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t14 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD93.t282 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2527 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.t8 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD99.t457 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2528 a_35949_n8931# CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t6 VSS.t749 VSS.t748 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2529 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VDD108.t234 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2530 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD93.t378 VDD93.t377 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2531 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 a_28546_n743# VSS.t2152 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2532 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.t5 a_21902_n8787# VSS.t539 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2533 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_42529_n14305# VSS.t399 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2534 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT VDD96.t93 VDD96.t92 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2535 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD110.t444 VDD110.t443 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2536 a_43793_n10116# CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t350 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2537 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 a_55020_n2199# VSS.t1830 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2538 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_4.IN2 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 VDD96.t187 VDD96.t186 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2539 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 VDD.t130 VDD.t129 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2540 a_54033_n15587# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT VSS.t1989 VSS.t1988 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2541 a_53095_n5765# VDD108.t463 VSS.t522 VSS.t521 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2542 VDD108 dec3x8_ibr_mag_0.and_3_ibr_3.nand3_mag_ibr_0.OUT VSS.t611 VSS.t610 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2543 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD96.t136 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2544 a_54537_n6818# CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS.t1060 VSS.t1059 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2545 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_26663_398# VSS.t1051 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2546 a_25640_n18723# CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t6 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS.t2384 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2547 VSS CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t7 a_27144_10099# VSS.t1178 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2548 a_45724_9057# CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t16 a_45564_9057# VSS.t2212 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2549 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 a_22718_8532# VDD90.t158 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X2550 Vdiv90 CLK_div_90_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 VSS.t2010 VSS.t2009 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X2551 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD96.t145 VDD96.t144 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2552 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT VDD108.t171 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2553 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 VDD100.t48 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2554 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t0 VDD108.t2 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2555 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD105.t181 VDD105.t180 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2556 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 VDD105.t369 VDD105.t368 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2557 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD99.t146 VDD99.t145 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2558 a_45899_7960# CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t12 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN VSS.t492 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2559 a_22301_6115# VDD90.t484 VSS.t205 VSS.t204 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2560 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD90.t95 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2561 a_47086_5143# VDD105.t490 VSS.t1111 VSS.t1110 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2562 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_45251_n1102# VSS.t1763 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2563 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB a_24944_n8778# VSS.t20 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2564 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t1 VDD105.t409 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2565 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.CLK VDD105.t303 VDD105.t302 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2566 CLK_div_96_mag_0.JK_FF_mag_0.Q CLK_div_96_mag_0.JK_FF_mag_0.QB a_24116_n1789# VSS.t415 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2567 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 a_46768_n5176# VSS.t308 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2568 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 VDD110.t88 VDD110.t87 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2569 a_23184_n9840# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS.t550 VSS.t549 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2570 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB VDD100.t47 VDD100.t46 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2571 a_33898_n18723# CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t1640 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2572 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD105.t278 VDD105.t277 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2573 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.t10 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VDD90.t176 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2574 CLK_div_99_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.t9 VDD99.t461 VDD99.t460 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2575 VSS CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN VSS.t913 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X2576 a_22565_n6009# RST.t106 a_22405_n6009# VSS.t2029 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2577 CLK_div_105_mag_0.CLK_div_10_mag_1.CLK CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 VSS.t1950 VSS.t1949 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X2578 a_22421_810# CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_4.IN2 VSS.t1534 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2579 a_55197_n20487# CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 VDD110.t305 VDD110.t304 pfet_03v3 ad=0.624p pd=2.92u as=1.06p ps=5.68u w=2.4u l=0.28u
X2580 a_23283_n7106# CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t15 a_23123_n7106# VSS.t268 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2581 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT VDD99.t392 VDD99.t391 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2582 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t23 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT VDD99.t181 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2583 VDD96 CLK_div_96_mag_0.JK_FF_mag_2.QB CLK_div_96_mag_0.JK_FF_mag_2.Q VDD96.t345 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2584 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB VDD99.t335 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2585 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t2 VDD105.t271 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2586 VDD108 CLK_div_108_new_mag_0.JK_FF_mag_0.QB Vdiv108.t0 VDD108.t193 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2587 a_51397_6284# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VSS.t624 VSS.t623 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2588 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t7 VDD105.t194 VDD105.t193 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2589 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_29270_n743# VSS.t1880 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2590 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD100.t199 VDD100.t198 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2591 a_43597_n6273# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t7 VSS.t1235 VSS.t493 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2592 VSS CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t12 a_23691_9000# VSS.t1183 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2593 VSS CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_28099_n17626# VSS.t1846 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2594 VDD105 VDD105.t41 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VDD105.t42 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2595 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 VDD90.t298 VDD90.t297 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2596 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD105.t38 VDD105.t40 VDD105.t39 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2597 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD99.t382 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2598 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD110.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2599 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.t0 VDD93.t135 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2600 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS.t423 VSS.t422 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X2601 a_23510_n15620# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 VDD99.t74 VDD99.t73 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X2602 a_39126_n8931# CLK_div_93_mag_0.CLK_div_3_mag_0.CLK a_38966_n8931# VSS.t696 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2603 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD90.t344 VDD90.t343 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2604 VDD96 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD96.t53 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2605 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD93.t62 VDD93.t61 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2606 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 a_33583_n16588# VSS.t2334 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2607 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VDD108.t150 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2608 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 VDD105.t218 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2609 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN VSS.t1302 VSS.t1301 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2610 a_48466_n6273# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t1031 VSS.t146 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2611 VDD F0.t20 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 VDD.t181 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2612 VSS VDD108.t464 a_45241_n10160# VSS.t523 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2613 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD110.t34 VDD110.t33 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2614 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 VDD110.t436 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2615 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD105.t231 VDD105.t230 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2616 a_44117_n2243# CLK.t70 a_43957_n2243# VSS.t2520 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2617 a_45695_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS.t1826 VSS.t1825 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2618 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD93.t312 VDD93.t311 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2619 a_52923_9057# CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t1 VSS.t816 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2620 a_26606_6159# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VSS.t1417 VSS.t1416 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2621 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD110.t228 VDD110.t227 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2622 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t10 a_44799_n7920# VSS.t2238 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2623 VDD100 VDD100.t71 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT VDD100.t72 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2624 a_38960_n10028# VDD93.t487 VSS.t248 VSS.t247 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2625 a_48023_n7840# CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 VDD108.t1 VDD108.t0 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X2626 a_54597_n15587# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 VSS.t1787 VSS.t1786 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2627 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK.t71 VDD90.t461 VDD90.t460 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2628 a_23743_5062# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS.t793 VSS.t792 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2629 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t14 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB VDD93.t288 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2630 a_35614_n16636# RST.t107 a_35454_n16636# VSS.t2028 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2631 VSS CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_22685_11196# VSS.t1310 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2632 VSS CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_26426_11196# VSS.t1864 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2633 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t1 VDD90.t140 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2634 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 VDD100.t351 VDD100.t350 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2635 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.t0 VDD99.t305 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2636 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD99.t87 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2637 VDD F2.t9 dec3x8_ibr_mag_0.and_3_ibr_6.nand3_mag_ibr_0.OUT VDD.t80 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2638 a_45235_n9063# CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t11 a_45075_n9063# VSS.t2241 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2639 a_24337_n6010# CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t16 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB VSS.t1004 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2640 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD110.t449 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2641 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD93.t314 VDD93.t313 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2642 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD93.t80 VDD93.t82 VDD93.t81 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2643 VDD108 VDD108.t13 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT VDD108.t14 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2644 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD93.t268 VDD93.t267 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2645 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_51961_6284# VSS.t366 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2646 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD100.t264 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2647 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN VSS.t586 VSS.t585 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X2648 VSS VDD105.t492 a_54775_9057# VSS.t1112 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2649 a_30398_n699# CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t1555 VSS.t1554 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2650 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 VDD105.t115 VDD105.t114 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2651 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t8 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 VDD96.t333 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2652 a_44511_n9019# CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t1511 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2653 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_37237_n8887# VSS.t2093 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2654 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD110.t61 VDD110.t60 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2655 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_48324_n15585# VSS.t1765 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2656 a_31512_6115# CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 a_31352_6115# VSS.t1625 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2657 VDD96 CLK_div_96_mag_0.JK_FF_mag_0.Q CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD96.t222 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2658 CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t7 a_40818_n8887# VSS.t750 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2659 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT CLK.t72 VDD108.t453 VDD108.t452 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2660 CLK_div_90_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT VDD90.t117 VDD90.t116 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X2661 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD105.t135 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2662 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD105.t332 VDD105.t331 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2663 a_47704_n1102# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VSS.t477 VSS.t476 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2664 VDD108 CLK_div_108_new_mag_0.JK_FF_mag_1.Q CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD108.t413 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2665 VSS VDD100.t492 a_51652_2768# VSS.t2415 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2666 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t12 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VSS.t2242 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2667 VDD99 dec3x8_ibr_mag_0.and_3_ibr_5.nand3_mag_ibr_0.OUT VDD.t118 VDD.t117 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2668 a_47264_n17599# VDD110.t499 VSS.t1018 VSS.t1017 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2669 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_45000_9057# VSS.t780 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2670 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VDD100.t21 VDD100.t20 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2671 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD110.t65 VDD110.t64 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2672 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD93.t194 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2673 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t17 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 VSS.t2213 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2674 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 a_49794_1671# VSS.t1965 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2675 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 VDD99.t346 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2676 VDD110 RST.t108 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VDD110.t395 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2677 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_27170_6159# VSS.t134 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2678 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.t7 a_51641_n9064# VSS.t1190 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2679 a_54621_10154# CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t18 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VSS.t2216 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2680 VSS CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS.t2149 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X2681 a_45564_9057# CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t7 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VSS.t1072 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2682 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD100.t219 VDD100.t218 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2683 a_35184_n1822# Vdiv93.t3 VSS.t2289 VSS.t2288 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2684 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD105.t414 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2685 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 VDD100.t347 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2686 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD99.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2687 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD93.t436 VDD93.t435 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2688 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VDD90.t41 VDD90.t40 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2689 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 a_49488_n13383# VSS.t1733 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2690 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK VSS.t1747 VSS.t1746 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2691 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t19 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN VDD105.t460 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2692 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 a_36103_n10028# VSS.t283 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2693 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.t7 VDD90.t449 VDD90.t448 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2694 a_50157_n1146# CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 a_49997_n1146# VSS.t880 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2695 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 VSS.t554 VSS.t553 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X2696 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD100.t168 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2697 VSS CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT a_25619_n7107# VSS.t1527 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2698 a_46259_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t137 VSS.t136 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2699 a_28657_n18723# CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS.t1407 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2700 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K VDD105.t362 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2701 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 a_24307_5062# VSS.t1624 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2702 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VDD110.t260 VDD110.t259 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2703 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VDD99.t331 VDD99.t330 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2704 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.t0 VDD108.t335 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2705 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t1 VDD105.t365 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2706 VDD Vdiv96.t3 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT VDD.t28 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2707 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 VDD93.t344 VDD93.t343 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2708 VSS CLK_div_90_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 VSS.t81 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2709 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_52293_n17599# VSS.t1892 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2710 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT RST.t109 VDD99.t359 VDD99.t358 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2711 VSS CLK.t73 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 VSS.t2521 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2712 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 a_46735_10154# VSS.t1139 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2713 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT VSS.t163 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2714 a_29270_n743# RST.t110 a_29110_n743# VSS.t2027 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2715 a_23691_9000# CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.t9 CLK_div_90_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS.t1183 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2716 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD90.t429 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2717 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_32794_5062# VSS.t1023 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2718 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VSS.t291 VSS.t290 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2719 a_29341_n16634# RST.t111 a_29181_n16634# VSS.t2026 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2720 VDD108 RST.t112 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD108.t344 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2721 VSS CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_32789_10099# VSS.t302 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2722 VSS CLK.t74 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 VSS.t2524 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2723 VSS CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t15 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VSS.t1127 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2724 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 VDD99.t323 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2725 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD105.t334 VDD105.t333 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2726 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD100.t463 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2727 a_35192_n17626# CLK.t75 a_35032_n17626# VSS.t2527 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2728 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 a_40972_n9984# VSS.t1940 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2729 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 VDD108.t126 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2730 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_40254_n8887# VSS.t704 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2731 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t20 a_45899_7960# VSS.t492 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2732 a_22466_n8743# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS.t1664 VSS.t1663 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2733 a_54947_n5721# CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t1662 VSS.t1661 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2734 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.t8 a_29862_n9832# VSS.t122 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2735 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_54302_n1102# VSS.t97 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2736 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD108.t273 VDD108.t272 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2737 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD108.t162 VDD108.t161 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2738 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 F1.t17 VSS.t1216 VSS.t1215 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2739 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 a_24391_n20290# VDD99.t406 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X2740 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 a_23956_n14213# VSS.t1576 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2741 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_50447_n18696# VSS.t1891 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2742 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT VSS.t768 VSS.t767 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X2743 VDD99 VDD99.t40 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD99.t41 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2744 a_39690_n8887# CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS.t1570 VSS.t1569 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2745 CLK_div_96_mag_0.JK_FF_mag_3.QB CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD96.t52 VDD96.t51 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2746 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 VSS.t791 VSS.t790 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X2747 VDD108 RST.t113 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD108.t341 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2748 a_50763_n10161# CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT VSS.t1904 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2749 VDD F2.t10 dec3x8_ibr_mag_0.and_3_ibr_2.nand3_mag_ibr_0.OUT VDD.t83 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2750 a_29680_398# CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t1879 VSS.t1878 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2751 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K VDD110.t244 VDD110.t243 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2752 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_43229_n10116# VSS.t78 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2753 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD110.t12 VDD110.t14 VDD110.t13 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2754 a_25488_n15535# CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t24 a_25328_n15535# VSS.t1253 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2755 a_23594_n8743# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t712 VSS.t711 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2756 CLK_div_100_mag_0.CLK_div_10_mag_1.CLK CLK_div_100_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 VSS.t461 VSS.t460 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X2757 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT VDD110.t365 VDD110.t364 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2758 a_32295_n16632# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT VSS.t1668 VSS.t1667 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2759 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t25 a_30210_n13332# VSS.t1254 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2760 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD100.t197 VDD100.t196 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2761 a_47988_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VSS.t978 VSS.t977 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2762 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_36024_n15495# VSS.t1368 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2763 a_26226_n9831# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS.t1925 VSS.t1924 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2764 a_25508_n8734# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS.t1371 VSS.t1370 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2765 VSS CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_25076_n18723# VSS.t1599 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2766 a_49122_n18696# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VSS.t620 VSS.t619 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2767 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT VDD110.t120 VDD110.t119 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2768 dec3x8_ibr_mag_0.and_3_ibr_6.nand3_mag_ibr_0.OUT dec3x8_ibr_mag_0.and_3_ibr_6.IN3 VDD.t46 VDD.t45 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2769 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_50304_n16724# VSS.t398 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2770 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 a_50353_n9020# VSS.t1901 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2771 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 Vdiv100.t0 VSS.t370 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X2772 a_32750_n7675# CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.t9 VDD93.t31 VDD93.t30 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X2773 a_30163_n17626# CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.t7 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K VSS.t1075 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2774 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB a_28016_n8779# VSS.t202 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2775 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD100.t118 VDD100.t117 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2776 VSS CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_25055_n7107# VSS.t1705 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2777 a_54775_9057# CLK_div_105_mag_0.CLK_div_10_mag_1.CLK a_54615_9057# VSS.t1556 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2778 VDD90 RST.t114 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VDD90.t225 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2779 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_53129_n19793# VSS.t1322 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2780 VSS CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN VSS.t1579 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X2781 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD110.t286 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2782 a_47252_6240# CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 a_47092_6240# VSS.t2112 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2783 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t26 VSS.t1256 VSS.t1255 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2784 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD105.t167 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2785 a_49789_n9020# CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.t7 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.t2 VSS.t2268 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2786 a_44229_5143# CLK.t76 a_44069_5143# VSS.t2528 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2787 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 VDD100.t396 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2788 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT VDD99.t12 VDD99.t11 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2789 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_52923_9057# VSS.t1429 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2790 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_36827_n10028# VSS.t1044 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2791 a_28010_n9876# CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t15 a_27850_n9876# VSS.t1006 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2792 mux_8x1_ibr_0.mux_2x1_ibr_0.I1 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 VDD.t4 VDD.t3 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2793 a_53168_n2243# CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 a_53008_n2243# VSS.t2455 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2794 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K VDD110.t240 VDD110.t239 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2795 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 a_49635_n10117# VSS.t1285 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2796 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 VDD108.t63 VDD108.t62 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2797 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_93_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS.t772 VSS.t771 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2798 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VDD100.t280 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X2799 a_49794_1671# CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t1 VSS.t1837 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2800 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 CLK_div_96_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD96.t362 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2801 a_27170_6159# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VSS.t89 VSS.t88 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2802 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 VDD96.t361 VDD96.t360 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2803 VDD90 CLK.t77 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VDD90.t462 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2804 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t1 VDD99.t219 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2805 VDD105 CLK.t78 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD105.t473 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2806 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t2 VDD96.t310 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2807 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t8 VDD108.t230 VDD108.t229 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2808 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN VSS.t559 VSS.t558 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2809 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD105.t328 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2810 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT a_50204_2768# VSS.t2182 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2811 VDD96 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD96.t258 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2812 VDD105 RST.t115 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VDD105.t387 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2813 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 VDD110.t206 VDD110.t205 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2814 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VDD110.t32 VDD110.t31 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X2815 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT VDD99.t261 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2816 VDD93 VDD93.t76 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD93.t77 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2817 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_45131_n17599# VSS.t2161 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2818 VSS CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_27529_n18723# VSS.t935 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2819 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD96.t146 VDD96.t148 VDD96.t147 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2820 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD96.t88 VDD96.t87 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2821 VSS VDD108.t466 a_54664_n10161# VSS.t526 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2822 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 VDD99.t422 VDD99.t421 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2823 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD108.t192 VDD108.t191 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2824 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.t0 VDD99.t284 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2825 a_38454_6265# F2.t11 a_38294_6265# VSS.t1206 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2826 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN VSS.t1365 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X2827 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT VDD93.t73 VDD93.t75 VDD93.t74 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2828 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS.t102 VSS.t101 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2829 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_23589_6159# VSS.t2254 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2830 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT a_35747_880# VSS.t1276 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2831 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 VDD.t32 VDD.t31 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2832 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t8 VDD93.t245 VDD93.t244 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2833 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_53819_n5721# VSS.t1058 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2834 a_48783_n13424# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_48623_n13424# VSS.t1801 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2835 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK VSS.t541 VSS.t540 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2836 mux_8x1_ibr_0.mux_2x1_ibr_0.I1 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT a_37999_880# VSS.t15 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2837 VSS CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_23403_10099# VSS.t112 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2838 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 VDD105.t413 VDD105.t412 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2839 a_32794_5062# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS.t471 VSS.t470 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2840 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 VSS.t2454 VSS.t2453 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2841 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD99.t202 VDD99.t201 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2842 a_54746_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS.t108 VSS.t107 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2843 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t8 a_53174_n1146# VSS.t1177 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2844 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD110.t306 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2845 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN CLK.t79 a_31129_n6271# VSS.t411 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2846 VSS CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_30727_n17626# VSS.t1147 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2847 VSS CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.CLK VSS.t2223 nfet_03v3 ad=86.8f pd=0.92u as=86.8f ps=0.92u w=0.22u l=0.28u
X2848 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD96.t15 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2849 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 a_55310_n17599# VSS.t2105 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2850 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN VDD93.t27 VDD93.t26 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X2851 a_31128_n7028# CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 VSS.t1508 VSS.t1507 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2852 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT VDD99.t7 VDD99.t6 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2853 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t0 VDD108.t7 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2854 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t16 VDD100.t431 VDD100.t430 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2855 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_45039_n5176# VSS.t145 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2856 a_54907_297# CLK_div_100_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 VDD100.t124 VDD100.t123 pfet_03v3 ad=0.624p pd=2.92u as=1.06p ps=5.68u w=2.4u l=0.28u
X2857 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 a_30209_7256# VSS.t2259 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2858 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 a_53280_5143# VSS.t1948 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2859 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 VDD110.t319 VDD110.t318 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2860 dec3x8_ibr_mag_0.and_3_ibr_2.nand3_mag_ibr_0.OUT dec3x8_ibr_mag_0.and_3_ibr_6.IN3 VDD.t44 VDD.t43 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2861 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD105.t353 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2862 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_96_mag_0.JK_FF_mag_0.Q VDD96.t221 VDD96.t220 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2863 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK.t80 VDD110.t488 VDD110.t487 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2864 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 VDD99.t420 VDD99.t418 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2865 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 VDD90.t428 VDD90.t427 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2866 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_0.Q VSS.t1692 VSS.t1691 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2867 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD93.t17 VDD93.t16 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2868 VDD96 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT VDD96.t190 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2869 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 a_25529_n743# VSS.t2548 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2870 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VDD110.t202 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2871 a_23249_11196# CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS.t1313 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2872 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I1 VDD.t154 VDD.t153 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2873 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_47994_n18696# VSS.t1996 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2874 VSS CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS.t2226 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X2875 a_21841_n6009# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VSS.t2017 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2876 a_53844_5143# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS.t1446 VSS.t1445 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2877 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t13 VDD108.t387 VDD108.t386 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2878 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS.t1041 VSS.t1040 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2879 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I1 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT a_36873_880# VSS.t1186 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2880 a_38454_6821# F2.t12 a_38294_6821# VSS.t1206 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2881 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_32865_n15491# VSS.t1396 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2882 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t14 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VDD108.t388 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2883 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 F0.t21 VDD.t185 VDD.t184 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2884 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_52161_n19793# VSS.t868 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2885 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I1 VDD.t142 VDD.t141 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2886 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 VDD93.t334 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2887 a_47092_6240# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t8 VSS.t861 VSS.t860 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2888 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD105.t283 VDD105.t282 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2889 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 VDD105.t378 VDD105.t377 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2890 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 a_28489_5018# VSS.t218 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2891 VDD93 CLK.t81 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 VDD93.t466 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2892 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD90.t21 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2893 a_44069_5143# VDD105.t493 VSS.t1116 VSS.t1115 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2894 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD100.t68 VDD100.t70 VDD100.t69 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2895 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 F0.t22 VSS.t2448 VSS.t2447 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2896 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 VDD110.t292 VDD110.t291 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2897 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_22620_n9884# VSS.t708 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2898 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD93.t202 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2899 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 VDD99.t190 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2900 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD110.t59 VDD110.t58 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2901 a_22711_n14504# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 a_22551_n14504# VSS.t1578 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2902 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT VDD99.t415 VDD99.t414 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2903 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD93.t70 VDD93.t72 VDD93.t71 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2904 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K VSS.t1945 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2905 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_51575_n18696# VSS.t831 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2906 a_25535_354# CLK_div_96_mag_0.JK_FF_mag_3.Q a_25375_354# VSS.t435 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2907 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN VSS.t1984 VSS.t1983 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X2908 a_53813_n6862# CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS.t153 VSS.t152 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2909 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t13 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VDD90.t262 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2910 a_29053_5018# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VSS.t1589 VSS.t1588 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2911 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN VSS.t1845 VSS.t1844 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2912 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 a_42083_n15712# VDD110.t163 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X2913 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK.t82 VDD90.t466 VDD90.t465 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2914 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB VDD90.t86 VDD90.t85 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2915 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_26253_n743# VSS.t173 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2916 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD105.t35 VDD105.t37 VDD105.t36 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2917 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 VSS.t1797 VSS.t1796 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X2918 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 VDD90.t426 VDD90.t425 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2919 a_55101_n6818# CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t297 VSS.t296 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2920 a_29116_398# CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS.t640 VSS.t639 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2921 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_25662_n9875# VSS.t1923 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X2922 a_25364_n19822# CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.t10 CLK_div_99_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS.t2360 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2923 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VDD108.t263 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2924 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT RST.t116 VDD90.t246 VDD90.t245 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2925 a_23973_11196# CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.t8 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS.t2387 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2926 a_29307_n1855# CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VSS.t594 VSS.t593 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2927 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VDD99.t30 VDD99.t29 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2928 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD90.t107 VDD90.t106 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2929 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 VDD110.t141 VDD110.t140 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2930 a_29905_n16590# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT VSS.t1281 VSS.t1280 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2931 VDD100 CLK.t83 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD100.t473 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2932 VDD110 RST.t117 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT VDD110.t392 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2933 VDD mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_2x1_ibr_0.I1 VDD.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2934 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB VDD93.t191 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2935 a_48747_10154# CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t15 a_48587_10154# VSS.t1229 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2936 a_47492_n5176# RST.t118 a_47332_n5176# VSS.t2025 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2937 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.t8 VDD108.t218 VDD108.t217 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2938 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD90.t49 VDD90.t51 VDD90.t50 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2939 VSS CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_34462_n18723# VSS.t2294 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2940 a_53304_n18696# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K VSS.t690 VSS.t689 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2941 a_38294_6265# dec3x8_ibr_mag_0.and_3_ibr_6.IN3 VSS.t785 VSS.t783 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2942 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 VDD110.t430 VDD110.t429 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2943 a_47299_10154# CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 VSS.t1137 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2944 a_23589_6159# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t949 VSS.t948 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2945 VDD mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 VDD.t40 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2946 VSS CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS.t721 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X2947 a_48478_n16682# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT VSS.t1672 VSS.t1671 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2948 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t15 VDD108.t392 VDD108.t391 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2949 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_45449_n6273# VSS.t146 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2950 a_50880_10154# CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT VSS.t1590 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2951 a_45452_1671# CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t7 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VSS.t536 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2952 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB VDD99.t258 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2953 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB VDD100.t277 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2954 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t8 a_33429_n15491# VSS.t1197 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2955 VDD99 dec3x8_ibr_mag_0.and_3_ibr_5.nand3_mag_ibr_0.OUT VSS.t1340 VSS.t279 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2956 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK.t84 VDD93.t470 VDD93.t469 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2957 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT RST.t119 VDD93.t393 VDD93.t392 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2958 a_37999_n1222# mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 VSS.t796 VSS.t795 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2959 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD110.t275 VDD110.t274 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2960 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VDD99.t34 VDD99.t33 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2961 a_29708_n8735# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 VSS.t2345 VSS.t2344 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2962 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K VDD99.t21 VDD99.t20 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2963 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD93.t154 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2964 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD93.t366 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2965 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 VSS.t1319 VSS.t1318 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2966 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK.t85 VDD110.t490 VDD110.t489 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X2967 VSS CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_22121_11196# VSS.t1736 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2968 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD105.t200 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2969 VDD110 CLK.t86 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT VDD110.t491 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2970 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB VDD90.t279 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2971 a_53280_5143# CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 a_53120_5143# VSS.t2111 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2972 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_52139_n18696# VSS.t1890 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2973 VSS CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 a_21431_n7106# VSS.t720 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2974 a_26974_1919# CLK.t87 a_26814_1919# VSS.t2529 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2975 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t14 VDD90.t266 VDD90.t265 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2976 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD110.t338 VDD110.t337 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2977 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_96_mag_0.JK_FF_mag_2.QB VDD96.t344 VDD96.t343 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2978 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD96.t305 VDD96.t304 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2979 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 a_49640_2768# VSS.t1602 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2980 a_53939_1671# CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t1264 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2981 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.t9 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT VDD108.t219 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2982 a_27334_n16588# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t1526 VSS.t1525 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2983 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_55161_n15587# VSS.t1807 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2984 a_39684_n10028# CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS.t1300 VSS.t1299 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2985 a_26349_n6010# CLK.t88 a_26189_n6010# VSS.t2530 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2986 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VDD90.t329 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2987 VSS CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 a_25122_1919# VSS.t337 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2988 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_23552_n1789# VSS.t1646 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2989 CLK_div_96_mag_0.JK_FF_mag_0.QB CLK_div_96_mag_0.JK_FF_mag_0.Q a_24270_n2886# VSS.t1690 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2990 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_24153_6159# VSS.t1019 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2991 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD90.t315 VDD90.t314 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2992 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_45343_n16680# VSS.t1546 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2993 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.t0 VDD108.t231 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X2994 a_38294_6821# dec3x8_ibr_mag_0.and_3_ibr_6.IN3 VSS.t784 VSS.t783 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2995 a_54498_n9064# CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT VSS.t643 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X2996 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT RST.t120 VDD90.t248 VDD90.t247 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X2997 a_49098_5187# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VSS.t1777 VSS.t1776 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X2998 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_51193_n19793# VSS.t868 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2999 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VDD90.t92 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3000 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VDD90.t5 VDD90.t4 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X3001 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VDD105.t132 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X3002 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD99.t299 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X3003 VSS CLK.t89 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VSS.t2531 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X3004 a_28489_5018# CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 a_28329_5018# VSS.t218 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X3005 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 VDD96.t309 VDD96.t308 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3006 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_44413_n18696# VSS.t1316 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X3007 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.t6 VDD93.t164 VDD93.t163 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3008 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VDD90.t319 VDD90.t318 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X3009 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 F0.t23 VDD.t187 VDD.t186 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X3010 VDD108 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD108.t282 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3011 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t12 VDD100.t233 VDD100.t232 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X3012 a_22982_n2930# CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS.t2089 VSS.t2088 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X3013 a_35186_n18723# CLK.t90 a_35026_n18723# VSS.t2534 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X3014 a_53738_n1102# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS.t851 VSS.t850 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X3015 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD108.t10 VDD108.t12 VDD108.t11 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X3016 a_54057_10154# RST.t121 a_53897_10154# VSS.t2024 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X3017 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t0 VDD100.t387 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3018 a_32015_n17626# CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.t8 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VSS.t1076 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X3019 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD110.t9 VDD110.t11 VDD110.t10 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X3020 a_34896_n15539# CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t27 a_34736_n15539# VSS.t1257 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X3021 a_37436_880# mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I1 VSS.t2181 VSS.t2180 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X3022 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_41284_n14596# VSS.t2186 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X3023 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 VSS.t2110 VSS.t2109 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X3024 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD96.t3 VDD96.t2 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X3025 a_29144_n8735# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 VSS.t1231 VSS.t1230 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X3026 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB VDD105.t374 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3027 a_54028_n18696# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS.t691 VSS.t109 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X3028 a_44357_n10160# CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VSS.t1488 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X3029 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_32640_6159# VSS.t1022 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X3030 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t7 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD99.t485 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3031 RST CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN VDD93.t361 VDD93.t360 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X3032 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VDD90.t422 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X3033 CLK_div_108_new_mag_0.JK_FF_mag_1.QB CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD108.t250 VDD108.t249 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X3034 a_47902_n6273# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t1029 VSS.t146 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X3035 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB VDD93.t9 VDD93.t8 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3036 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD90.t345 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X3037 Vdiv96 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VDD96.t50 VDD96.t49 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X3038 a_46810_n10116# CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t361 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X3039 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD100.t160 VDD100.t159 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X3040 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN VSS.t809 VSS.t808 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X3041 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t15 VDD90.t268 VDD90.t267 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X3042 a_36178_n16592# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT VSS.t1379 VSS.t1378 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X3043 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN VDD110.t84 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3044 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_28623_n15537# VSS.t2348 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X3045 VSS CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT Vdiv110.t0 VSS.t1619 nfet_03v3 ad=86.8f pd=0.92u as=86.8f ps=0.92u w=0.22u l=0.28u
X3046 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.t2 VDD108.t155 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3047 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS.t1745 VSS.t1744 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X3048 VSS CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN VSS.t562 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X3049 a_26096_3016# CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT VSS.t1550 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X3050 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t7 a_48252_n9063# VSS.t993 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X3051 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 VDD90.t294 VDD90.t293 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X3052 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD110.t6 VDD110.t5 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X3053 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD108.t47 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3054 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB VDD90.t419 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3055 a_29213_5018# RST.t122 a_29053_5018# VSS.t2023 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X3056 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD96.t271 VDD96.t270 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3057 a_26778_n1855# CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VSS.t2144 VSS.t2143 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X3058 a_27496_n2952# CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VSS.t1699 VSS.t1697 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X3059 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 a_54187_n16728# VSS.t1785 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X3060 VDD110 RST.t123 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT VDD110.t389 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X3061 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.t10 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD90.t242 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X3062 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD99.t245 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3063 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 VDD110.t428 VDD110.t427 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X3064 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_47528_n9019# VSS.t572 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X3065 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD99.t229 VDD99.t228 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X3066 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_37391_n9984# VSS.t2092 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X3067 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 a_29298_n9832# VSS.t2130 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X3068 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_36673_n8887# VSS.t188 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X3069 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB VDD110.t351 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3070 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN VDD93.t186 VDD93.t185 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X3071 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_45907_n16680# VSS.t552 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X3072 VSS CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_52769_10154# VSS.t628 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X3073 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD96.t132 VDD96.t131 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X3074 a_33513_10099# CLK.t91 a_33353_10099# VSS.t2535 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X3075 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD100.t25 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3076 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VDD90.t153 VDD90.t152 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X3077 a_28392_354# CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 VSS.t2547 VSS.t2546 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X3078 CLK_div_108_new_mag_0.CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.t10 VDD108.t223 VDD108.t222 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X3079 a_30165_n6282# CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 VSS.t2301 VSS.t450 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X3080 a_44235_6240# CLK.t92 a_44075_6240# VSS.t2536 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X3081 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD100.t440 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X3082 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB VDD110.t347 VDD110.t346 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3083 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 a_30469_n16590# VSS.t2350 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X3084 a_39402_n7788# CLK_div_93_mag_0.CLK_div_3_mag_0.CLK VSS.t695 VSS.t694 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X3085 a_33405_7558# CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT a_33245_7558# VDD90.t408 pfet_03v3 ad=0.624p pd=2.92u as=0.624p ps=2.92u w=2.4u l=0.28u
X3086 VDD96 CLK_div_96_mag_0.JK_FF_mag_5.Q.t12 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD96.t120 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X3087 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 VDD99.t419 VDD99.t418 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X3088 a_47816_6284# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VSS.t845 VSS.t844 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X3089 a_36310_880# Vdiv110.t5 VSS.t752 VSS.t751 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X3090 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD108.t175 VDD108.t174 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X3091 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD108.t252 VDD108.t251 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X3092 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_96_mag_0.JK_FF_mag_3.QB a_28743_n1899# VSS.t447 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X3093 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_29461_n2996# VSS.t1610 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X3094 a_50987_5143# RST.t124 a_50827_5143# VSS.t2022 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X3095 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 VDD110.t122 VDD110.t121 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X3096 CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.t8 VSS.t1080 VSS.t1079 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X3097 VDD96 dec3x8_ibr_mag_0.and_3_ibr_1.nand3_mag_ibr_0.OUT VDD.t16 VDD.t15 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X3098 VSS VDD108.t467 a_48258_n10160# VSS.t529 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X3099 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB VDD90.t111 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3100 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VDD110.t183 VDD110.t182 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X3101 a_26072_n8734# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t1922 VSS.t1921 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X3102 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 a_50151_n2243# VSS.t1034 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X3103 a_48712_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VSS.t1995 VSS.t1994 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X3104 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VDD110.t105 VDD110.t104 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X3105 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VSS.t917 VSS.t916 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X3106 a_29241_7256# CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 VSS.t2258 VSS.t2257 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X3107 a_23948_n13382# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 VDD99.t257 VDD99.t256 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X3108 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_2.OUT CLK_div_96_mag_0.JK_FF_mag_4.Q.t11 VDD96.t127 VDD96.t126 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X3109 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VDD93.t472 VDD93.t471 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X3110 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t0 VDD99.t26 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3111 a_22839_10099# CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t112 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X3112 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 a_33812_n13270# VDD99.t345 pfet_03v3 ad=1.06p pd=5.68u as=0.624p ps=2.92u w=2.4u l=0.28u
X3113 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD105.t20 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3114 a_26214_n1855# CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VSS.t1696 VSS.t1695 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X3115 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 F0.t24 a_36310_n1822# VSS.t2436 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X3116 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 VSS.t1623 VSS.t1622 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X3117 VSS CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_46964_n9019# VSS.t1288 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X3118 a_50903_n5# CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 VSS.t879 VSS.t878 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X3119 VSS CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_53939_1671# VSS.t37 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X3120 a_31577_n15535# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K VSS.t2124 VSS.t2123 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X3121 a_28574_n9876# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT VSS.t2165 VSS.t2164 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X3122 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT VDD110.t181 VDD110.t180 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X3123 Vdiv99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT VSS.t1974 VSS.t1973 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X3124 VDD108 RST.t125 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD108.t338 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X3125 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t16 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VDD93.t427 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3126 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_48380_6284# VSS.t1774 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X3127 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t5 VDD110.t448 VDD110.t447 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X3128 VDD96 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VDD96.t204 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3129 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.t8 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT VDD108.t410 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X3130 a_26817_n699# CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS.t177 VSS.t176 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X3131 a_43826_n7684# CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.t8 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN VDD108.t372 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X3132 a_45517_5187# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS.t788 VSS.t787 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X3133 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 VDD108.t360 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3134 a_23869_810# CLK_div_96_mag_0.JK_FF_mag_4.Q.t12 a_23709_810# VSS.t1220 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X3135 a_54503_1671# CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VSS.t983 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X3136 VDD Vdiv100.t5 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT VDD.t155 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3137 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK.t93 VSS.t2538 VSS.t2537 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X3138 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT VSS.t1448 VSS.t1447 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X3139 VDD100 VDD100.t64 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT VDD100.t65 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3140 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT VDD110.t285 VDD110.t284 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X3141 a_48944_6284# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VSS.t87 VSS.t86 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X3142 a_23956_n14213# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 VSS.t1577 VSS.t1576 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X3143 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 F2.t13 VDD.t87 VDD.t86 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X3144 a_35184_880# Vdiv105.t5 VSS.t2379 VSS.t2378 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X3145 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN VDD110.t97 VDD110.t96 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X3146 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VDD93.t262 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3147 a_25650_n1899# CLK_div_96_mag_0.JK_FF_mag_0.Q a_25490_n1899# VSS.t1689 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X3148 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VDD93.t382 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3149 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t16 VDD105.t248 VDD105.t247 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X3150 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 F0.t25 VSS.t2438 VSS.t2437 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X3151 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD110.t424 VDD110.t423 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
R0 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n3 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t3 37.1981
R1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n5 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t4 31.4332
R2 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n4 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t5 30.4613
R3 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n4 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t7 24.7562
R4 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n3 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t2 17.6611
R5 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n5 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t6 15.3826
R6 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n0 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 12.0716
R7 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n5 7.62076
R8 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n6 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 6.09789
R9 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n7 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n2 2.99416
R10 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n2 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t0 2.2755
R11 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n2 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n1 2.2755
R12 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n7 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n6 2.2505
R13 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n0 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 2.24788
R14 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n6 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n0 1.94903
R15 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n4 1.81638
R16 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n3 1.43706
R17 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n7 0.4325
R18 VDD90.n162 VDD90.n15 11185.2
R19 VDD90.n202 VDD90.n195 11185.2
R20 VDD90.n235 VDD90.n227 11185.2
R21 VDD90.n142 VDD90.t83 1105.93
R22 VDD90.t92 VDD90.t98 961.905
R23 VDD90.t85 VDD90.t90 961.905
R24 VDD90.t24 VDD90.t11 961.905
R25 VDD90.t35 VDD90.t277 961.905
R26 VDD90.t120 VDD90.t411 961.905
R27 VDD90.t201 VDD90.t209 961.905
R28 VDD90.t198 VDD90.t176 765.152
R29 VDD90.t337 VDD90.t135 765.152
R30 VDD90.t279 VDD90.t2 765.152
R31 VDD90.t100 VDD90.t368 765.152
R32 VDD90.t334 VDD90.t138 765.152
R33 VDD90.t189 VDD90.t0 765.152
R34 VDD90.t161 VDD90.t376 765.152
R35 VDD90.t323 VDD90.t332 765.152
R36 VDD90.t179 VDD90.t4 765.152
R37 VDD90.t143 VDD90.t220 765.152
R38 VDD90.t326 VDD90.t329 765.152
R39 VDD90.t140 VDD90.t6 765.152
R40 VDD90.t21 VDD90.t30 765.152
R41 VDD90.t314 VDD90.t318 765.152
R42 VDD90.t425 VDD90.t156 765.152
R43 VDD90.t249 VDD90.t308 765.152
R44 VDD90.t106 VDD90.t388 765.152
R45 VDD90.t340 VDD90.t122 765.152
R46 VDD90.t385 VDD90.t242 765.152
R47 VDD90.t391 VDD90.t108 765.152
R48 VDD90.t111 VDD90.t124 765.152
R49 VDD90.t403 VDD90.t27 765.152
R50 VDD90.t287 VDD90.t285 765.152
R51 VDD90.t269 VDD90.t152 765.152
R52 VDD90.t149 VDD90.t445 765.152
R53 VDD90.t290 VDD90.t282 765.152
R54 VDD90.t373 VDD90.t154 765.152
R55 VDD90.t414 VDD90.t417 765.152
R56 VDD90.t196 VDD90.t187 765.152
R57 VDD90.t364 VDD90.t217 765.152
R58 VDD90.t394 VDD90.t211 765.152
R59 VDD90.t128 VDD90.t133 765.152
R60 VDD90.t469 VDD90.t228 765.152
R61 VDD90.t214 VDD90.t437 765.152
R62 VDD90.t131 VDD90.t126 765.152
R63 VDD90.t383 VDD90.t182 765.152
R64 VDD90.t95 VDD90.t409 765.152
R65 VDD90.t45 VDD90.t40 765.152
R66 VDD90.t297 VDD90.t343 765.152
R67 VDD90.n138 VDD90.t396 747.159
R68 VDD90.t47 VDD90.n15 676.191
R69 VDD90.n195 VDD90.t316 676.191
R70 VDD90.n227 VDD90.t194 676.191
R71 VDD90.t114 VDD90.t116 645.307
R72 VDD90.n162 VDD90.t70 485.714
R73 VDD90.n202 VDD90.t230 485.714
R74 VDD90.t57 VDD90.n235 485.714
R75 VDD90 VDD90.n96 429.187
R76 VDD90.n153 VDD90 427.092
R77 VDD90.n148 VDD90 427.092
R78 VDD90 VDD90.n439 426.699
R79 VDD90 VDD90.n503 426.699
R80 VDD90 VDD90.n287 426.699
R81 VDD90.n309 VDD90 426.699
R82 VDD90.t427 VDD90.n162 426.44
R83 VDD90.t366 VDD90.n202 426.44
R84 VDD90.n235 VDD90.t16 426.44
R85 VDD90.n143 VDD90 425.019
R86 VDD90.n395 VDD90 424.618
R87 VDD90.n230 VDD90 424.618
R88 VDD90 VDD90.n397 418.495
R89 VDD90 VDD90.n210 418.495
R90 VDD90.n148 VDD90.t362 386.365
R91 VDD90.n153 VDD90.t293 386.365
R92 VDD90.n439 VDD90.t164 386.365
R93 VDD90.n503 VDD90.t171 386.365
R94 VDD90.n287 VDD90.t400 386.365
R95 VDD90.t235 VDD90.n309 386.365
R96 VDD90.n96 VDD90.t467 386.365
R97 VDD90.t422 VDD90.t85 380.952
R98 VDD90.t359 VDD90.t35 380.952
R99 VDD90.t209 VDD90.t13 380.952
R100 VDD90.t303 VDD90.n143 378.788
R101 VDD90.t434 VDD90.n148 378.788
R102 VDD90.t300 VDD90.n153 378.788
R103 VDD90.n397 VDD90.t174 378.788
R104 VDD90.n210 VDD90.t240 378.788
R105 VDD90.n397 VDD90.t311 322.223
R106 VDD90.t158 VDD90.n210 322.223
R107 VDD90.t219 VDD90.n395 320.635
R108 VDD90.t439 VDD90.n230 320.635
R109 VDD90.t176 VDD90.t450 303.031
R110 VDD90.t247 VDD90.t337 303.031
R111 VDD90.t368 VDD90.t452 303.031
R112 VDD90.t460 VDD90.t161 303.031
R113 VDD90.t220 VDD90.t465 303.031
R114 VDD90.t245 VDD90.t326 303.031
R115 VDD90.t440 VDD90.t314 303.031
R116 VDD90.t345 VDD90.t425 303.031
R117 VDD90.t308 VDD90.t265 303.031
R118 VDD90.t242 VDD90.t257 303.031
R119 VDD90.t443 VDD90.t391 303.031
R120 VDD90.t255 VDD90.t403 303.031
R121 VDD90.t445 VDD90.t267 303.031
R122 VDD90.t275 VDD90.t290 303.031
R123 VDD90.t272 VDD90.t196 303.031
R124 VDD90.t18 VDD90.t364 303.031
R125 VDD90.t228 VDD90.t348 303.031
R126 VDD90.t203 VDD90.t131 303.031
R127 VDD90.t353 VDD90.t383 303.031
R128 VDD90.t225 VDD90.t45 303.031
R129 VDD90.t429 VDD90.t297 303.031
R130 VDD90.t42 VDD90.n15 285.714
R131 VDD90.n195 VDD90.t320 285.714
R132 VDD90.n227 VDD90.t184 285.714
R133 VDD90.n123 VDD90.t87 242.857
R134 VDD90.n124 VDD90.t92 242.857
R135 VDD90.n160 VDD90.t42 242.857
R136 VDD90.n161 VDD90.t422 242.857
R137 VDD90.n163 VDD90.t32 242.857
R138 VDD90.n165 VDD90.t24 242.857
R139 VDD90.t320 VDD90.n168 242.857
R140 VDD90.n201 VDD90.t359 242.857
R141 VDD90.n221 VDD90.t206 242.857
R142 VDD90.n226 VDD90.t411 242.857
R143 VDD90.n237 VDD90.t184 242.857
R144 VDD90.t13 VDD90.n236 242.857
R145 VDD90.n144 VDD90.t303 193.183
R146 VDD90.n149 VDD90.t434 193.183
R147 VDD90.n154 VDD90.t300 193.183
R148 VDD90.n368 VDD90.t419 193.183
R149 VDD90.n370 VDD90.t21 193.183
R150 VDD90.n373 VDD90.t440 193.183
R151 VDD90.n376 VDD90.t345 193.183
R152 VDD90.n175 VDD90.t356 193.183
R153 VDD90.n177 VDD90.t414 193.183
R154 VDD90.n180 VDD90.t272 193.183
R155 VDD90.n183 VDD90.t18 193.183
R156 VDD90.n83 VDD90.t232 193.183
R157 VDD90.n89 VDD90.t211 193.183
R158 VDD90.n90 VDD90.t128 193.183
R159 VDD90.n95 VDD90.t348 193.183
R160 VDD90.n28 VDD90.t380 193.183
R161 VDD90.n30 VDD90.t214 193.183
R162 VDD90.n33 VDD90.t203 193.183
R163 VDD90.n36 VDD90.t353 193.183
R164 VDD90.n99 VDD90.t295 193.183
R165 VDD90.n101 VDD90.t95 193.183
R166 VDD90.n104 VDD90.t225 193.183
R167 VDD90.n107 VDD90.t429 193.183
R168 VDD90.t174 VDD90.n7 191.288
R169 VDD90.t450 VDD90.n422 191.288
R170 VDD90.n423 VDD90.t247 191.288
R171 VDD90.t2 VDD90.n431 191.288
R172 VDD90.n432 VDD90.t169 191.288
R173 VDD90.t452 VDD90.n442 191.288
R174 VDD90.t138 VDD90.n446 191.288
R175 VDD90.t0 VDD90.n451 191.288
R176 VDD90.n452 VDD90.t371 191.288
R177 VDD90.n502 VDD90.t460 191.288
R178 VDD90.n501 VDD90.t332 191.288
R179 VDD90.t4 VDD90.n467 191.288
R180 VDD90.n469 VDD90.t167 191.288
R181 VDD90.t465 VDD90.n480 191.288
R182 VDD90.n481 VDD90.t245 191.288
R183 VDD90.t6 VDD90.n489 191.288
R184 VDD90.n490 VDD90.t223 191.288
R185 VDD90.t240 VDD90.n208 191.288
R186 VDD90.t265 VDD90.n296 191.288
R187 VDD90.n297 VDD90.t106 191.288
R188 VDD90.t122 VDD90.n303 191.288
R189 VDD90.n304 VDD90.t306 191.288
R190 VDD90.t257 VDD90.n271 191.288
R191 VDD90.n272 VDD90.t443 191.288
R192 VDD90.t124 VDD90.n280 191.288
R193 VDD90.n281 VDD90.t238 191.288
R194 VDD90.n348 VDD90.t255 191.288
R195 VDD90.n347 VDD90.t285 191.288
R196 VDD90.t152 VDD90.n313 191.288
R197 VDD90.n315 VDD90.t398 191.288
R198 VDD90.t267 VDD90.n326 191.288
R199 VDD90.n327 VDD90.t275 191.288
R200 VDD90.t154 VDD90.n335 191.288
R201 VDD90.n336 VDD90.t448 191.288
R202 VDD90.t408 VDD90.t379 175.631
R203 VDD90.t396 VDD90.n3 153.678
R204 VDD90.n396 VDD90.t219 142.857
R205 VDD90.n231 VDD90.t439 142.857
R206 VDD90.t98 VDD90.n123 138.095
R207 VDD90.n124 VDD90.t47 138.095
R208 VDD90.t90 VDD90.n160 138.095
R209 VDD90.t70 VDD90.n161 138.095
R210 VDD90.t11 VDD90.n163 138.095
R211 VDD90.t316 VDD90.n165 138.095
R212 VDD90.t277 VDD90.n168 138.095
R213 VDD90.t230 VDD90.n201 138.095
R214 VDD90.n221 VDD90.t120 138.095
R215 VDD90.t194 VDD90.n226 138.095
R216 VDD90.n237 VDD90.t201 138.095
R217 VDD90.n236 VDD90.t57 138.095
R218 VDD90.n7 VDD90.t454 111.743
R219 VDD90.n422 VDD90.t80 111.743
R220 VDD90.n423 VDD90.t198 111.743
R221 VDD90.n431 VDD90.t135 111.743
R222 VDD90.n432 VDD90.t279 111.743
R223 VDD90.n442 VDD90.t164 111.743
R224 VDD90.n446 VDD90.t100 111.743
R225 VDD90.n451 VDD90.t334 111.743
R226 VDD90.n452 VDD90.t189 111.743
R227 VDD90.t171 VDD90.n502 111.743
R228 VDD90.t376 VDD90.n501 111.743
R229 VDD90.n467 VDD90.t323 111.743
R230 VDD90.n469 VDD90.t179 111.743
R231 VDD90.n480 VDD90.t60 111.743
R232 VDD90.n481 VDD90.t143 111.743
R233 VDD90.n489 VDD90.t329 111.743
R234 VDD90.n490 VDD90.t140 111.743
R235 VDD90.n208 VDD90.t259 111.743
R236 VDD90.n296 VDD90.t400 111.743
R237 VDD90.n297 VDD90.t249 111.743
R238 VDD90.n303 VDD90.t388 111.743
R239 VDD90.n304 VDD90.t340 111.743
R240 VDD90.n271 VDD90.t76 111.743
R241 VDD90.n272 VDD90.t385 111.743
R242 VDD90.n280 VDD90.t108 111.743
R243 VDD90.n281 VDD90.t111 111.743
R244 VDD90.n348 VDD90.t235 111.743
R245 VDD90.t27 VDD90.n347 111.743
R246 VDD90.n313 VDD90.t287 111.743
R247 VDD90.n315 VDD90.t269 111.743
R248 VDD90.n326 VDD90.t53 111.743
R249 VDD90.n327 VDD90.t149 111.743
R250 VDD90.n335 VDD90.t282 111.743
R251 VDD90.n336 VDD90.t373 111.743
R252 VDD90.t311 VDD90.n396 111.112
R253 VDD90.n231 VDD90.t158 111.112
R254 VDD90.n144 VDD90.t362 109.849
R255 VDD90.n149 VDD90.t293 109.849
R256 VDD90.n154 VDD90.t432 109.849
R257 VDD90.t30 VDD90.n368 109.849
R258 VDD90.t318 VDD90.n370 109.849
R259 VDD90.t156 VDD90.n373 109.849
R260 VDD90.n376 VDD90.t67 109.849
R261 VDD90.t417 VDD90.n175 109.849
R262 VDD90.t187 VDD90.n177 109.849
R263 VDD90.t217 VDD90.n180 109.849
R264 VDD90.n183 VDD90.t64 109.849
R265 VDD90.n83 VDD90.t394 109.849
R266 VDD90.t133 VDD90.n89 109.849
R267 VDD90.n90 VDD90.t469 109.849
R268 VDD90.t467 VDD90.n95 109.849
R269 VDD90.t437 VDD90.n28 109.849
R270 VDD90.t126 VDD90.n30 109.849
R271 VDD90.t182 VDD90.n33 109.849
R272 VDD90.n36 VDD90.t50 109.849
R273 VDD90.t409 VDD90.n99 109.849
R274 VDD90.t40 VDD90.n101 109.849
R275 VDD90.t343 VDD90.n104 109.849
R276 VDD90.n107 VDD90.t73 109.849
R277 VDD90.n439 VDD90.t457 62.1896
R278 VDD90.n503 VDD90.t462 62.1896
R279 VDD90.n287 VDD90.t262 62.1896
R280 VDD90.n309 VDD90.t252 62.1896
R281 VDD90.n395 VDD90.t37 61.8817
R282 VDD90.n230 VDD90.t103 61.8817
R283 VDD90.n397 VDD90.t146 60.9761
R284 VDD90.n210 VDD90.t8 60.9761
R285 VDD90.n96 VDD90.t351 59.702
R286 VDD90.n148 VDD90.t192 59.4064
R287 VDD90.n153 VDD90.t406 59.4064
R288 VDD90.n143 VDD90.t114 59.1138
R289 VDD90.t83 VDD90.n138 55.0852
R290 VDD90.t116 VDD90.n142 55.0852
R291 VDD90.n409 VDD90.t59 30.9379
R292 VDD90.n261 VDD90.t52 30.9379
R293 VDD90.n37 VDD90.t49 30.9379
R294 VDD90.n39 VDD90.t66 30.9379
R295 VDD90.n60 VDD90.t69 30.721
R296 VDD90.n50 VDD90.t56 30.7203
R297 VDD90.n57 VDD90.t72 30.3459
R298 VDD90.n412 VDD90.t79 30.2877
R299 VDD90.n260 VDD90.t75 30.2877
R300 VDD90.n45 VDD90.t63 30.0062
R301 VDD90.n57 VDD90.t476 24.8618
R302 VDD90.n413 VDD90.t479 24.5101
R303 VDD90.n409 VDD90.t471 24.5101
R304 VDD90.n259 VDD90.t480 24.5101
R305 VDD90.n261 VDD90.t473 24.5101
R306 VDD90.n37 VDD90.t472 24.5101
R307 VDD90.n39 VDD90.t478 24.5101
R308 VDD90.n60 VDD90.t477 24.4816
R309 VDD90.n50 VDD90.t484 24.4814
R310 VDD90.n47 VDD90.t481 24.4392
R311 VDD90.n3 VDD90.t408 21.9544
R312 VDD90 VDD90.t427 10.5649
R313 VDD90.t16 VDD90 10.5649
R314 VDD90 VDD90.t366 10.5649
R315 VDD90.n515 VDD90.n513 8.64529
R316 VDD90.n263 VDD90.n262 8.14231
R317 VDD90.n411 VDD90.n410 8.14083
R318 VDD90.n414 VDD90.n413 8.0005
R319 VDD90.n259 VDD90.n258 8.0005
R320 VDD90.n47 VDD90.n46 8.0005
R321 VDD90 VDD90.n512 7.36838
R322 VDD90.n67 VDD90.n66 6.39748
R323 VDD90 VDD90.n221 6.30459
R324 VDD90.n422 VDD90.n421 6.3005
R325 VDD90.n424 VDD90.n423 6.3005
R326 VDD90.n431 VDD90.n430 6.3005
R327 VDD90.n433 VDD90.n432 6.3005
R328 VDD90.n442 VDD90.n441 6.3005
R329 VDD90.n446 VDD90.n445 6.3005
R330 VDD90.n451 VDD90.n450 6.3005
R331 VDD90.n453 VDD90.n452 6.3005
R332 VDD90.n480 VDD90.n479 6.3005
R333 VDD90.n482 VDD90.n481 6.3005
R334 VDD90.n489 VDD90.n488 6.3005
R335 VDD90.n491 VDD90.n490 6.3005
R336 VDD90.n501 VDD90.n500 6.3005
R337 VDD90.n497 VDD90.n467 6.3005
R338 VDD90.n494 VDD90.n469 6.3005
R339 VDD90.n502 VDD90.n459 6.3005
R340 VDD90.n400 VDD90.n7 6.3005
R341 VDD90.n396 VDD90.n11 6.3005
R342 VDD90.n377 VDD90.n376 6.3005
R343 VDD90.n380 VDD90.n373 6.3005
R344 VDD90.n383 VDD90.n370 6.3005
R345 VDD90.n386 VDD90.n368 6.3005
R346 VDD90.n236 VDD90.n219 6.3005
R347 VDD90.n232 VDD90.n231 6.3005
R348 VDD90.n238 VDD90.n237 6.3005
R349 VDD90.n226 VDD90.n225 6.3005
R350 VDD90.n245 VDD90.n208 6.3005
R351 VDD90.n296 VDD90.n295 6.3005
R352 VDD90.n298 VDD90.n297 6.3005
R353 VDD90.n303 VDD90.n302 6.3005
R354 VDD90.n305 VDD90.n304 6.3005
R355 VDD90.n282 VDD90.n281 6.3005
R356 VDD90.n280 VDD90.n279 6.3005
R357 VDD90.n273 VDD90.n272 6.3005
R358 VDD90.n271 VDD90.n270 6.3005
R359 VDD90.n326 VDD90.n325 6.3005
R360 VDD90.n328 VDD90.n327 6.3005
R361 VDD90.n335 VDD90.n334 6.3005
R362 VDD90.n337 VDD90.n336 6.3005
R363 VDD90.n347 VDD90.n346 6.3005
R364 VDD90.n343 VDD90.n313 6.3005
R365 VDD90.n340 VDD90.n315 6.3005
R366 VDD90.n349 VDD90.n348 6.3005
R367 VDD90.n184 VDD90.n183 6.3005
R368 VDD90.n187 VDD90.n180 6.3005
R369 VDD90.n190 VDD90.n177 6.3005
R370 VDD90.n193 VDD90.n175 6.3005
R371 VDD90.n201 VDD90.n200 6.3005
R372 VDD90.n357 VDD90.n168 6.3005
R373 VDD90.n361 VDD90.n165 6.3005
R374 VDD90.n364 VDD90.n163 6.3005
R375 VDD90.n161 VDD90.n14 6.3005
R376 VDD90.n71 VDD90.n36 6.3005
R377 VDD90.n74 VDD90.n33 6.3005
R378 VDD90.n77 VDD90.n30 6.3005
R379 VDD90.n80 VDD90.n28 6.3005
R380 VDD90.n95 VDD90.n94 6.3005
R381 VDD90.n91 VDD90.n90 6.3005
R382 VDD90.n89 VDD90.n88 6.3005
R383 VDD90.n84 VDD90.n83 6.3005
R384 VDD90.n108 VDD90.n107 6.3005
R385 VDD90.n111 VDD90.n104 6.3005
R386 VDD90.n114 VDD90.n101 6.3005
R387 VDD90.n117 VDD90.n99 6.3005
R388 VDD90.n160 VDD90.n159 6.3005
R389 VDD90.n125 VDD90.n124 6.3005
R390 VDD90.n123 VDD90.n122 6.3005
R391 VDD90.n155 VDD90.n154 6.3005
R392 VDD90.n150 VDD90.n149 6.3005
R393 VDD90.n145 VDD90.n144 6.3005
R394 VDD90.n142 VDD90.n141 6.3005
R395 VDD90.n138 VDD90 6.3005
R396 VDD90.n511 VDD90.n3 6.3005
R397 VDD90.n242 VDD90.n211 5.85007
R398 VDD90.n56 VDD90.n55 5.30657
R399 VDD90.n479 VDD90.n475 5.213
R400 VDD90.n377 VDD90.t68 5.213
R401 VDD90.n325 VDD90.n321 5.213
R402 VDD90.n184 VDD90.t65 5.213
R403 VDD90.n108 VDD90.t74 5.213
R404 VDD90.n234 VDD90.t58 5.16878
R405 VDD90.n239 VDD90.t202 5.16878
R406 VDD90.n209 VDD90.t195 5.16878
R407 VDD90.n356 VDD90.t278 5.16878
R408 VDD90.n366 VDD90.n365 5.16878
R409 VDD90 VDD90.t17 5.16454
R410 VDD90 VDD90.n438 5.16369
R411 VDD90 VDD90.n286 5.16369
R412 VDD90.n4 VDD90.t139 5.15997
R413 VDD90.n299 VDD90.t107 5.15997
R414 VDD90.n171 VDD90.n170 5.15997
R415 VDD90.n140 VDD90.t117 5.14212
R416 VDD90.n458 VDD90.n457 5.13287
R417 VDD90.n407 VDD90.n406 5.13287
R418 VDD90.n426 VDD90.n403 5.13287
R419 VDD90.n429 VDD90.t3 5.13287
R420 VDD90.n428 VDD90.n427 5.13287
R421 VDD90.n434 VDD90.t170 5.13287
R422 VDD90.n440 VDD90.n437 5.13287
R423 VDD90.n444 VDD90.n443 5.13287
R424 VDD90.n448 VDD90.n447 5.13287
R425 VDD90.n449 VDD90.t1 5.13287
R426 VDD90.n436 VDD90.n435 5.13287
R427 VDD90.n454 VDD90.t372 5.13287
R428 VDD90.n465 VDD90.n460 5.13287
R429 VDD90.n499 VDD90.t333 5.13287
R430 VDD90.n498 VDD90.n466 5.13287
R431 VDD90.n496 VDD90.t5 5.13287
R432 VDD90.n495 VDD90.n468 5.13287
R433 VDD90.n493 VDD90.t168 5.13287
R434 VDD90.n474 VDD90.n473 5.13287
R435 VDD90.n484 VDD90.n470 5.13287
R436 VDD90.n487 VDD90.t7 5.13287
R437 VDD90.n486 VDD90.n485 5.13287
R438 VDD90.n492 VDD90.t224 5.13287
R439 VDD90.n401 VDD90.n6 5.13287
R440 VDD90.n399 VDD90.t175 5.13287
R441 VDD90.n379 VDD90.t157 5.13287
R442 VDD90.n382 VDD90.t319 5.13287
R443 VDD90.n384 VDD90.n369 5.13287
R444 VDD90.n385 VDD90.t31 5.13287
R445 VDD90.n387 VDD90.n367 5.13287
R446 VDD90.n246 VDD90.n207 5.13287
R447 VDD90.n244 VDD90.t241 5.13287
R448 VDD90.n224 VDD90.n220 5.13287
R449 VDD90.n223 VDD90.t121 5.13287
R450 VDD90.n215 VDD90.n214 5.13287
R451 VDD90.n251 VDD90.n250 5.13287
R452 VDD90.n288 VDD90.n285 5.13287
R453 VDD90.n293 VDD90.n292 5.13287
R454 VDD90.n300 VDD90.n284 5.13287
R455 VDD90.n301 VDD90.t123 5.13287
R456 VDD90.n306 VDD90.t307 5.13287
R457 VDD90.n257 VDD90.n256 5.13287
R458 VDD90.n275 VDD90.n253 5.13287
R459 VDD90.n278 VDD90.t125 5.13287
R460 VDD90.n277 VDD90.n276 5.13287
R461 VDD90.n283 VDD90.t239 5.13287
R462 VDD90.n311 VDD90.n310 5.13287
R463 VDD90.n345 VDD90.t286 5.13287
R464 VDD90.n344 VDD90.n312 5.13287
R465 VDD90.n342 VDD90.t153 5.13287
R466 VDD90.n341 VDD90.n314 5.13287
R467 VDD90.n339 VDD90.t399 5.13287
R468 VDD90.n320 VDD90.n319 5.13287
R469 VDD90.n330 VDD90.n316 5.13287
R470 VDD90.n333 VDD90.t155 5.13287
R471 VDD90.n332 VDD90.n331 5.13287
R472 VDD90.n338 VDD90.t449 5.13287
R473 VDD90.n205 VDD90.n173 5.13287
R474 VDD90.n186 VDD90.t218 5.13287
R475 VDD90.n189 VDD90.t188 5.13287
R476 VDD90.n191 VDD90.n176 5.13287
R477 VDD90.n192 VDD90.t418 5.13287
R478 VDD90.n194 VDD90.n174 5.13287
R479 VDD90.n199 VDD90.t231 5.13287
R480 VDD90.n358 VDD90.n167 5.13287
R481 VDD90.n359 VDD90.t317 5.13287
R482 VDD90.n362 VDD90.n164 5.13287
R483 VDD90.n363 VDD90.t12 5.13287
R484 VDD90.n390 VDD90.t71 5.13287
R485 VDD90.n20 VDD90.t468 5.13287
R486 VDD90.n92 VDD90.t470 5.13287
R487 VDD90.n24 VDD90.n23 5.13287
R488 VDD90.n87 VDD90.t134 5.13287
R489 VDD90.n86 VDD90.n25 5.13287
R490 VDD90.n85 VDD90.t395 5.13287
R491 VDD90.n82 VDD90.n26 5.13287
R492 VDD90.n73 VDD90.t183 5.13287
R493 VDD90.n76 VDD90.t127 5.13287
R494 VDD90.n78 VDD90.n29 5.13287
R495 VDD90.n79 VDD90.t438 5.13287
R496 VDD90.n81 VDD90.n27 5.13287
R497 VDD90.n110 VDD90.t344 5.13287
R498 VDD90.n113 VDD90.t41 5.13287
R499 VDD90.n115 VDD90.n100 5.13287
R500 VDD90.n116 VDD90.t410 5.13287
R501 VDD90.n118 VDD90.n98 5.13287
R502 VDD90.n158 VDD90.t91 5.13287
R503 VDD90.n127 VDD90.n16 5.13287
R504 VDD90.n126 VDD90.t48 5.13287
R505 VDD90.n18 VDD90.n17 5.13287
R506 VDD90.n121 VDD90.t99 5.13287
R507 VDD90.n120 VDD90.n19 5.13287
R508 VDD90.n156 VDD90.t433 5.13287
R509 VDD90.n132 VDD90.n131 5.13287
R510 VDD90.n151 VDD90.t294 5.13287
R511 VDD90.n134 VDD90.n133 5.13287
R512 VDD90.n146 VDD90.t363 5.13287
R513 VDD90.n136 VDD90.n135 5.13287
R514 VDD90 VDD90.n514 5.13104
R515 VDD90.n139 VDD90.t84 5.09693
R516 VDD90.n504 VDD90.n456 5.09407
R517 VDD90.n398 VDD90.n8 5.09407
R518 VDD90.n394 VDD90.n12 5.09407
R519 VDD90.n389 VDD90.t428 5.09407
R520 VDD90.n229 VDD90.n228 5.09407
R521 VDD90.n308 VDD90.n252 5.09407
R522 VDD90.n203 VDD90.t367 5.09407
R523 VDD90.n97 VDD90.t352 5.09407
R524 VDD90.n152 VDD90.t407 5.09407
R525 VDD90.n147 VDD90.t193 5.09407
R526 VDD90.n137 VDD90.t115 5.09407
R527 VDD90.n417 VDD90.n416 4.8755
R528 VDD90.n266 VDD90.n265 4.8755
R529 VDD90.n70 VDD90.t51 4.8755
R530 VDD90.n66 VDD90.n56 4.84121
R531 VDD90.n48 VDD90.n47 4.5005
R532 VDD90.n51 VDD90.n49 4.5005
R533 VDD90.n52 VDD90.n49 4.5005
R534 VDD90.n40 VDD90.n38 4.5005
R535 VDD90.n41 VDD90.n38 4.5005
R536 VDD90.n61 VDD90.n59 4.5005
R537 VDD90.n62 VDD90.n59 4.5005
R538 VDD90.n10 VDD90.n9 4.12326
R539 VDD90.n213 VDD90.n212 4.12326
R540 VDD90.n510 VDD90.t397 3.94862
R541 VDD90.n45 VDD90.n44 3.61662
R542 VDD90.n2 VDD90.n1 2.88497
R543 VDD90.n294 VDD90.n290 2.88497
R544 VDD90.n67 VDD90.n37 2.88182
R545 VDD90.n420 VDD90.n419 2.85787
R546 VDD90.n425 VDD90.n405 2.85787
R547 VDD90.n464 VDD90.n462 2.85787
R548 VDD90.n478 VDD90.n477 2.85787
R549 VDD90.n483 VDD90.n472 2.85787
R550 VDD90.n378 VDD90.n375 2.85787
R551 VDD90.n381 VDD90.n372 2.85787
R552 VDD90.n218 VDD90.n217 2.85787
R553 VDD90.n269 VDD90.n268 2.85787
R554 VDD90.n274 VDD90.n255 2.85787
R555 VDD90.n249 VDD90.n248 2.85787
R556 VDD90.n324 VDD90.n323 2.85787
R557 VDD90.n329 VDD90.n318 2.85787
R558 VDD90.n185 VDD90.n182 2.85787
R559 VDD90.n188 VDD90.n179 2.85787
R560 VDD90.n198 VDD90.n197 2.85787
R561 VDD90.n93 VDD90.n22 2.85787
R562 VDD90.n72 VDD90.n35 2.85787
R563 VDD90.n75 VDD90.n32 2.85787
R564 VDD90.n109 VDD90.n106 2.85787
R565 VDD90.n112 VDD90.n103 2.85787
R566 VDD90.n130 VDD90.n129 2.85787
R567 VDD90 VDD90.n515 2.59663
R568 VDD90.n419 VDD90.t451 2.2755
R569 VDD90.n419 VDD90.n418 2.2755
R570 VDD90.n405 VDD90.t248 2.2755
R571 VDD90.n405 VDD90.n404 2.2755
R572 VDD90.n1 VDD90.t453 2.2755
R573 VDD90.n1 VDD90.n0 2.2755
R574 VDD90.n462 VDD90.t461 2.2755
R575 VDD90.n462 VDD90.n461 2.2755
R576 VDD90.n477 VDD90.t466 2.2755
R577 VDD90.n477 VDD90.n476 2.2755
R578 VDD90.n472 VDD90.t246 2.2755
R579 VDD90.n472 VDD90.n471 2.2755
R580 VDD90.n375 VDD90.t426 2.2755
R581 VDD90.n375 VDD90.n374 2.2755
R582 VDD90.n372 VDD90.t315 2.2755
R583 VDD90.n372 VDD90.n371 2.2755
R584 VDD90.n217 VDD90.t210 2.2755
R585 VDD90.n217 VDD90.n216 2.2755
R586 VDD90.n290 VDD90.t266 2.2755
R587 VDD90.n290 VDD90.n289 2.2755
R588 VDD90.n268 VDD90.t258 2.2755
R589 VDD90.n268 VDD90.n267 2.2755
R590 VDD90.n255 VDD90.t444 2.2755
R591 VDD90.n255 VDD90.n254 2.2755
R592 VDD90.n248 VDD90.t256 2.2755
R593 VDD90.n248 VDD90.n247 2.2755
R594 VDD90.n323 VDD90.t268 2.2755
R595 VDD90.n323 VDD90.n322 2.2755
R596 VDD90.n318 VDD90.t276 2.2755
R597 VDD90.n318 VDD90.n317 2.2755
R598 VDD90.n182 VDD90.t365 2.2755
R599 VDD90.n182 VDD90.n181 2.2755
R600 VDD90.n179 VDD90.t197 2.2755
R601 VDD90.n179 VDD90.n178 2.2755
R602 VDD90.n197 VDD90.t36 2.2755
R603 VDD90.n197 VDD90.n196 2.2755
R604 VDD90.n22 VDD90.t229 2.2755
R605 VDD90.n22 VDD90.n21 2.2755
R606 VDD90.n35 VDD90.t384 2.2755
R607 VDD90.n35 VDD90.n34 2.2755
R608 VDD90.n32 VDD90.t132 2.2755
R609 VDD90.n32 VDD90.n31 2.2755
R610 VDD90.n106 VDD90.t298 2.2755
R611 VDD90.n106 VDD90.n105 2.2755
R612 VDD90.n103 VDD90.t46 2.2755
R613 VDD90.n103 VDD90.n102 2.2755
R614 VDD90.n129 VDD90.t86 2.2755
R615 VDD90.n129 VDD90.n128 2.2755
R616 VDD90.n54 VDD90.n53 2.2439
R617 VDD90.n64 VDD90.n63 2.2439
R618 VDD90.n43 VDD90.n42 2.24362
R619 VDD90.n40 VDD90.n39 2.12257
R620 VDD90.n410 VDD90.n409 2.11346
R621 VDD90.n262 VDD90.n261 2.11346
R622 VDD90.n263 VDD90.n260 1.8236
R623 VDD90.n412 VDD90.n411 1.82345
R624 VDD90 VDD90.n458 1.81843
R625 VDD90.n440 VDD90 1.81843
R626 VDD90 VDD90.n251 1.81843
R627 VDD90.n288 VDD90 1.81843
R628 VDD90.n58 VDD90.n57 1.81789
R629 VDD90.n390 VDD90 1.77285
R630 VDD90 VDD90.n20 1.77285
R631 VDD90 VDD90.n151 1.77285
R632 VDD90 VDD90.n146 1.77285
R633 VDD90 VDD90.n234 1.70433
R634 VDD90.n55 VDD90.n54 1.62565
R635 VDD90.n65 VDD90.n64 1.62565
R636 VDD90.n61 VDD90.n60 1.39782
R637 VDD90.n51 VDD90.n50 1.39728
R638 VDD90.n82 VDD90.n81 1.16167
R639 VDD90.n493 VDD90.n492 1.16051
R640 VDD90.n339 VDD90.n338 1.16051
R641 VDD90.n55 VDD90.n48 1.12171
R642 VDD90.n65 VDD90.n58 1.12171
R643 VDD90.n388 VDD90.n387 1.07428
R644 VDD90.n204 VDD90.n194 1.07428
R645 VDD90.n119 VDD90.n118 1.07428
R646 VDD90.n307 VDD90.n283 1.0737
R647 VDD90.n455 VDD90.n434 1.01824
R648 VDD90.n47 VDD90.n45 0.840632
R649 VDD90.n234 VDD90.n233 0.788255
R650 VDD90.n233 VDD90.n229 0.760634
R651 VDD90.n157 VDD90.n156 0.715235
R652 VDD90.n206 VDD90.n205 0.671656
R653 VDD90.n266 VDD90.n264 0.608132
R654 VDD90.n240 VDD90.n239 0.593661
R655 VDD90.n243 VDD90.n209 0.593661
R656 VDD90.n353 VDD90.n172 0.593661
R657 VDD90.n356 VDD90.n355 0.593661
R658 VDD90.n366 VDD90.n13 0.593661
R659 VDD90.n360 VDD90.n166 0.557288
R660 VDD90.n392 VDD90.n391 0.557288
R661 VDD90.n66 VDD90.n65 0.5228
R662 VDD90.n56 VDD90.n43 0.497812
R663 VDD90.n222 VDD90.n206 0.488955
R664 VDD90.n463 VDD90 0.468385
R665 VDD90 VDD90.n350 0.468385
R666 VDD90.n233 VDD90.n213 0.439524
R667 VDD90.n413 VDD90.n412 0.404541
R668 VDD90.n260 VDD90.n259 0.404541
R669 VDD90.n512 VDD90.n2 0.369535
R670 VDD90.n508 VDD90.n4 0.369535
R671 VDD90.n294 VDD90.n291 0.369535
R672 VDD90.n299 VDD90.n169 0.369535
R673 VDD90.n354 VDD90.n171 0.369535
R674 VDD90.n507 VDD90.n5 0.342778
R675 VDD90.n506 VDD90.n505 0.342778
R676 VDD90.n509 VDD90 0.338387
R677 VDD90.n421 VDD90.n417 0.337997
R678 VDD90.n270 VDD90.n266 0.337997
R679 VDD90.n71 VDD90.n70 0.337997
R680 VDD90.n140 VDD90 0.334577
R681 VDD90.n70 VDD90.n69 0.333658
R682 VDD90.n352 VDD90.n206 0.329033
R683 VDD90.n417 VDD90.n415 0.328132
R684 VDD90.n141 VDD90.n139 0.317357
R685 VDD90.n392 VDD90.n13 0.312894
R686 VDD90.n507 VDD90.n506 0.280925
R687 VDD90.n241 VDD90.n213 0.277085
R688 VDD90.n353 VDD90.n352 0.274194
R689 VDD90.n420 VDD90.n407 0.233919
R690 VDD90.n426 VDD90.n425 0.233919
R691 VDD90.n478 VDD90.n474 0.233919
R692 VDD90.n484 VDD90.n483 0.233919
R693 VDD90.n382 VDD90.n381 0.233919
R694 VDD90.n379 VDD90.n378 0.233919
R695 VDD90.n269 VDD90.n257 0.233919
R696 VDD90.n275 VDD90.n274 0.233919
R697 VDD90.n324 VDD90.n320 0.233919
R698 VDD90.n330 VDD90.n329 0.233919
R699 VDD90.n189 VDD90.n188 0.233919
R700 VDD90.n186 VDD90.n185 0.233919
R701 VDD90.n76 VDD90.n75 0.233919
R702 VDD90.n73 VDD90.n72 0.233919
R703 VDD90.n113 VDD90.n112 0.233919
R704 VDD90.n110 VDD90.n109 0.233919
R705 VDD90.n506 VDD90.n402 0.226218
R706 VDD90.n508 VDD90.n507 0.221851
R707 VDD90.n351 VDD90 0.184731
R708 VDD90.n152 VDD90.n132 0.170231
R709 VDD90.n147 VDD90.n134 0.170231
R710 VDD90.n137 VDD90.n136 0.170231
R711 VDD90.n393 VDD90.n392 0.169866
R712 VDD90.n515 VDD90 0.163082
R713 VDD90.n354 VDD90.n353 0.161388
R714 VDD90.n291 VDD90.n13 0.154438
R715 VDD90.n139 VDD90 0.147133
R716 VDD90.n307 VDD90.n306 0.143967
R717 VDD90.n205 VDD90.n204 0.143501
R718 VDD90.n120 VDD90.n119 0.143501
R719 VDD90.n429 VDD90.n428 0.141016
R720 VDD90.n487 VDD90.n486 0.141016
R721 VDD90.n499 VDD90.n498 0.141016
R722 VDD90.n496 VDD90.n495 0.141016
R723 VDD90.n385 VDD90.n384 0.141016
R724 VDD90.n224 VDD90.n223 0.141016
R725 VDD90.n278 VDD90.n277 0.141016
R726 VDD90.n333 VDD90.n332 0.141016
R727 VDD90.n345 VDD90.n344 0.141016
R728 VDD90.n342 VDD90.n341 0.141016
R729 VDD90.n192 VDD90.n191 0.141016
R730 VDD90.n359 VDD90.n358 0.141016
R731 VDD90.n363 VDD90.n362 0.141016
R732 VDD90.n79 VDD90.n78 0.141016
R733 VDD90.n86 VDD90.n85 0.141016
R734 VDD90.n87 VDD90.n24 0.141016
R735 VDD90.n116 VDD90.n115 0.141016
R736 VDD90.n121 VDD90.n18 0.141016
R737 VDD90.n127 VDD90.n126 0.141016
R738 VDD90.n308 VDD90.n307 0.139745
R739 VDD90.n389 VDD90.n388 0.138896
R740 VDD90.n119 VDD90.n97 0.138896
R741 VDD90.n394 VDD90.n393 0.137219
R742 VDD90.n169 VDD90.n166 0.132199
R743 VDD90.n455 VDD90.n454 0.130793
R744 VDD90.n355 VDD90.n354 0.128029
R745 VDD90 VDD90.n203 0.127858
R746 VDD90.n291 VDD90.n166 0.126986
R747 VDD90.n355 VDD90.n169 0.125597
R748 VDD90.n444 VDD90 0.123016
R749 VDD90.n465 VDD90 0.123016
R750 VDD90 VDD90.n293 0.123016
R751 VDD90.n311 VDD90 0.123016
R752 VDD90 VDD90.n92 0.122435
R753 VDD90 VDD90.n402 0.122231
R754 VDD90.n218 VDD90 0.111984
R755 VDD90.n198 VDD90 0.111984
R756 VDD90.n93 VDD90 0.111984
R757 VDD90 VDD90.n130 0.111984
R758 VDD90 VDD90.n464 0.111403
R759 VDD90 VDD90.n249 0.111403
R760 VDD90.n58 VDD90 0.110941
R761 VDD90.n410 VDD90 0.107393
R762 VDD90.n262 VDD90 0.107393
R763 VDD90.n430 VDD90.n429 0.107339
R764 VDD90.n434 VDD90.n433 0.107339
R765 VDD90.n450 VDD90.n449 0.107339
R766 VDD90.n454 VDD90.n453 0.107339
R767 VDD90.n488 VDD90.n487 0.107339
R768 VDD90.n492 VDD90.n491 0.107339
R769 VDD90.n500 VDD90.n499 0.107339
R770 VDD90.n497 VDD90.n496 0.107339
R771 VDD90.n494 VDD90.n493 0.107339
R772 VDD90.n387 VDD90.n386 0.107339
R773 VDD90.n384 VDD90.n383 0.107339
R774 VDD90.n238 VDD90.n215 0.107339
R775 VDD90.n225 VDD90.n224 0.107339
R776 VDD90.n302 VDD90.n301 0.107339
R777 VDD90.n306 VDD90.n305 0.107339
R778 VDD90.n279 VDD90.n278 0.107339
R779 VDD90.n283 VDD90.n282 0.107339
R780 VDD90.n334 VDD90.n333 0.107339
R781 VDD90.n338 VDD90.n337 0.107339
R782 VDD90.n346 VDD90.n345 0.107339
R783 VDD90.n343 VDD90.n342 0.107339
R784 VDD90.n340 VDD90.n339 0.107339
R785 VDD90.n194 VDD90.n193 0.107339
R786 VDD90.n191 VDD90.n190 0.107339
R787 VDD90.n362 VDD90.n361 0.107339
R788 VDD90.n358 VDD90.n357 0.107339
R789 VDD90.n81 VDD90.n80 0.107339
R790 VDD90.n78 VDD90.n77 0.107339
R791 VDD90.n84 VDD90.n82 0.107339
R792 VDD90.n88 VDD90.n86 0.107339
R793 VDD90.n91 VDD90.n24 0.107339
R794 VDD90.n118 VDD90.n117 0.107339
R795 VDD90.n115 VDD90.n114 0.107339
R796 VDD90.n122 VDD90.n120 0.107339
R797 VDD90.n125 VDD90.n18 0.107339
R798 VDD90.n159 VDD90.n127 0.107339
R799 VDD90.n155 VDD90.n132 0.107339
R800 VDD90.n150 VDD90.n134 0.107339
R801 VDD90.n145 VDD90.n136 0.107339
R802 VDD90 VDD90.n420 0.106758
R803 VDD90.n425 VDD90 0.106758
R804 VDD90 VDD90.n478 0.106758
R805 VDD90.n483 VDD90 0.106758
R806 VDD90 VDD90.n269 0.106758
R807 VDD90.n274 VDD90 0.106758
R808 VDD90 VDD90.n324 0.106758
R809 VDD90.n329 VDD90 0.106758
R810 VDD90.n381 VDD90 0.106177
R811 VDD90.n378 VDD90 0.106177
R812 VDD90 VDD90.n218 0.106177
R813 VDD90.n188 VDD90 0.106177
R814 VDD90.n185 VDD90 0.106177
R815 VDD90 VDD90.n198 0.106177
R816 VDD90.n130 VDD90 0.106177
R817 VDD90.n75 VDD90 0.106177
R818 VDD90.n72 VDD90 0.106177
R819 VDD90 VDD90.n93 0.106177
R820 VDD90.n112 VDD90 0.106177
R821 VDD90.n109 VDD90 0.106177
R822 VDD90.n393 VDD90.n11 0.1004
R823 VDD90.n258 VDD90 0.100075
R824 VDD90.n509 VDD90.n508 0.0980478
R825 VDD90 VDD90.n10 0.0975258
R826 VDD90.n46 VDD90 0.0839415
R827 VDD90.n215 VDD90.n209 0.0835323
R828 VDD90.n157 VDD90 0.082371
R829 VDD90.n52 VDD90 0.0816915
R830 VDD90.n424 VDD90.n407 0.080629
R831 VDD90.n441 VDD90.n440 0.080629
R832 VDD90.n482 VDD90.n474 0.080629
R833 VDD90.n380 VDD90.n379 0.080629
R834 VDD90.n295 VDD90.n288 0.080629
R835 VDD90.n273 VDD90.n257 0.080629
R836 VDD90.n328 VDD90.n320 0.080629
R837 VDD90.n187 VDD90.n186 0.080629
R838 VDD90.n200 VDD90.n199 0.080629
R839 VDD90.n74 VDD90.n73 0.080629
R840 VDD90.n94 VDD90.n20 0.080629
R841 VDD90.n111 VDD90.n110 0.080629
R842 VDD90.n62 VDD90 0.0805665
R843 VDD90.n402 VDD90.n401 0.0795385
R844 VDD90 VDD90.n385 0.0794677
R845 VDD90 VDD90.n382 0.0794677
R846 VDD90 VDD90.n192 0.0794677
R847 VDD90 VDD90.n189 0.0794677
R848 VDD90 VDD90.n363 0.0794677
R849 VDD90 VDD90.n79 0.0794677
R850 VDD90 VDD90.n76 0.0794677
R851 VDD90.n85 VDD90 0.0794677
R852 VDD90 VDD90.n87 0.0794677
R853 VDD90.n92 VDD90 0.0794677
R854 VDD90 VDD90.n116 0.0794677
R855 VDD90 VDD90.n113 0.0794677
R856 VDD90 VDD90.n121 0.0794677
R857 VDD90.n126 VDD90 0.0794677
R858 VDD90 VDD90.n158 0.0794677
R859 VDD90 VDD90.n140 0.0794623
R860 VDD90 VDD90.n426 0.0788871
R861 VDD90.n428 VDD90 0.0788871
R862 VDD90 VDD90.n444 0.0788871
R863 VDD90 VDD90.n448 0.0788871
R864 VDD90 VDD90.n436 0.0788871
R865 VDD90 VDD90.n484 0.0788871
R866 VDD90.n486 VDD90 0.0788871
R867 VDD90 VDD90.n465 0.0788871
R868 VDD90.n498 VDD90 0.0788871
R869 VDD90.n495 VDD90 0.0788871
R870 VDD90.n293 VDD90 0.0788871
R871 VDD90 VDD90.n300 0.0788871
R872 VDD90 VDD90.n275 0.0788871
R873 VDD90.n277 VDD90 0.0788871
R874 VDD90 VDD90.n330 0.0788871
R875 VDD90.n332 VDD90 0.0788871
R876 VDD90 VDD90.n311 0.0788871
R877 VDD90.n344 VDD90 0.0788871
R878 VDD90.n341 VDD90 0.0788871
R879 VDD90.n156 VDD90 0.0759839
R880 VDD90.n151 VDD90 0.0759839
R881 VDD90.n146 VDD90 0.0759839
R882 VDD90.n436 VDD90.n5 0.0754032
R883 VDD90.n366 VDD90.n364 0.0748226
R884 VDD90.n41 VDD90 0.0738165
R885 VDD90.n299 VDD90.n298 0.0730806
R886 VDD90.n69 VDD90.n67 0.0725
R887 VDD90 VDD90.n172 0.0717592
R888 VDD90.n241 VDD90.n240 0.071388
R889 VDD90 VDD90.n389 0.0709717
R890 VDD90.n203 VDD90 0.0709717
R891 VDD90.n97 VDD90 0.0709717
R892 VDD90 VDD90.n152 0.0709717
R893 VDD90 VDD90.n147 0.0709717
R894 VDD90 VDD90.n137 0.0709717
R895 VDD90.n505 VDD90.n455 0.0708636
R896 VDD90.n399 VDD90.n398 0.0704581
R897 VDD90 VDD90.n394 0.0701226
R898 VDD90 VDD90.n229 0.0701226
R899 VDD90 VDD90.n308 0.0701226
R900 VDD90.n68 VDD90 0.0700455
R901 VDD90.n360 VDD90.n359 0.0695968
R902 VDD90.n408 VDD90 0.0690714
R903 VDD90.n449 VDD90.n5 0.0661129
R904 VDD90 VDD90.n510 0.0659817
R905 VDD90.n243 VDD90 0.0656
R906 VDD90.n388 VDD90.n366 0.0639524
R907 VDD90 VDD90.n294 0.0614677
R908 VDD90.n242 VDD90.n241 0.0611
R909 VDD90.n301 VDD90.n171 0.0608871
R910 VDD90.n239 VDD90 0.0603065
R911 VDD90.n391 VDD90.n390 0.0562419
R912 VDD90.n400 VDD90.n399 0.0557
R913 VDD90.n245 VDD90.n244 0.0557
R914 VDD90.n463 VDD90.n458 0.0556613
R915 VDD90.n350 VDD90.n251 0.0556613
R916 VDD90 VDD90.n356 0.0556613
R917 VDD90.n445 VDD90.n4 0.0550806
R918 VDD90.n504 VDD90 0.0546389
R919 VDD90.n223 VDD90.n222 0.0515968
R920 VDD90 VDD90.n2 0.0510161
R921 VDD90.n415 VDD90.n408 0.0471071
R922 VDD90.n69 VDD90.n68 0.0455
R923 VDD90 VDD90.n10 0.0437
R924 VDD90.n510 VDD90 0.0432575
R925 VDD90.n505 VDD90.n504 0.0430455
R926 VDD90.n448 VDD90.n4 0.0428871
R927 VDD90.n464 VDD90.n463 0.0417258
R928 VDD90.n350 VDD90.n249 0.0417258
R929 VDD90.n158 VDD90.n157 0.0405645
R930 VDD90.n401 VDD90 0.0392
R931 VDD90.n246 VDD90 0.0392
R932 VDD90.n414 VDD90.n411 0.0387493
R933 VDD90.n199 VDD90.n172 0.0382419
R934 VDD90.n351 VDD90.n246 0.038
R935 VDD90.n234 VDD90.n219 0.0370806
R936 VDD90.n415 VDD90.n414 0.0358571
R937 VDD90.n264 VDD90.n263 0.0344878
R938 VDD90.n356 VDD90 0.0341774
R939 VDD90.n244 VDD90.n243 0.0311
R940 VDD90.n239 VDD90 0.0295323
R941 VDD90.n53 VDD90.n52 0.0275
R942 VDD90.n46 VDD90.n44 0.0275
R943 VDD90.n63 VDD90.n62 0.026375
R944 VDD90.n54 VDD90.n49 0.025705
R945 VDD90.n64 VDD90.n59 0.025705
R946 VDD90 VDD90.n209 0.0248871
R947 VDD90.n300 VDD90.n299 0.0248871
R948 VDD90.n391 VDD90.n14 0.0248871
R949 VDD90.n398 VDD90 0.0243065
R950 VDD90.n222 VDD90 0.0242273
R951 VDD90.n240 VDD90 0.0234344
R952 VDD90 VDD90.n509 0.0211312
R953 VDD90.n42 VDD90.n41 0.02075
R954 VDD90.n463 VDD90.n459 0.0206923
R955 VDD90.n350 VDD90.n349 0.0206923
R956 VDD90.n233 VDD90.n232 0.017527
R957 VDD90.n43 VDD90.n38 0.0169383
R958 VDD90 VDD90.n2 0.0167581
R959 VDD90.n352 VDD90.n351 0.0157185
R960 VDD90.n264 VDD90.n258 0.0119894
R961 VDD90.n204 VDD90 0.0115377
R962 VDD90 VDD90.n360 0.010371
R963 VDD90.n42 VDD90.n40 0.0095
R964 VDD90.n408 VDD90 0.00907143
R965 VDD90 VDD90.n171 0.00862903
R966 VDD90.n294 VDD90 0.00630645
R967 VDD90 VDD90.n155 0.00514516
R968 VDD90 VDD90.n150 0.00514516
R969 VDD90 VDD90.n145 0.00514516
R970 VDD90.n68 VDD90 0.00459091
R971 VDD90.n63 VDD90.n61 0.003875
R972 VDD90.n512 VDD90.n511 0.00378904
R973 VDD90 VDD90.n400 0.0032
R974 VDD90 VDD90.n245 0.0032
R975 VDD90.n232 VDD90 0.00293243
R976 VDD90.n53 VDD90.n51 0.00275
R977 VDD90.n11 VDD90 0.0026
R978 VDD90.n430 VDD90 0.00224194
R979 VDD90.n433 VDD90 0.00224194
R980 VDD90.n445 VDD90 0.00224194
R981 VDD90.n450 VDD90 0.00224194
R982 VDD90.n453 VDD90 0.00224194
R983 VDD90.n488 VDD90 0.00224194
R984 VDD90.n491 VDD90 0.00224194
R985 VDD90.n500 VDD90 0.00224194
R986 VDD90 VDD90.n497 0.00224194
R987 VDD90 VDD90.n494 0.00224194
R988 VDD90.n298 VDD90 0.00224194
R989 VDD90.n302 VDD90 0.00224194
R990 VDD90.n305 VDD90 0.00224194
R991 VDD90.n279 VDD90 0.00224194
R992 VDD90.n282 VDD90 0.00224194
R993 VDD90.n334 VDD90 0.00224194
R994 VDD90.n337 VDD90 0.00224194
R995 VDD90.n346 VDD90 0.00224194
R996 VDD90 VDD90.n343 0.00224194
R997 VDD90 VDD90.n340 0.00224194
R998 VDD90.n141 VDD90 0.00219811
R999 VDD90.n386 VDD90 0.00166129
R1000 VDD90.n383 VDD90 0.00166129
R1001 VDD90 VDD90.n380 0.00166129
R1002 VDD90 VDD90.n377 0.00166129
R1003 VDD90.n219 VDD90 0.00166129
R1004 VDD90 VDD90.n238 0.00166129
R1005 VDD90.n225 VDD90 0.00166129
R1006 VDD90.n193 VDD90 0.00166129
R1007 VDD90.n190 VDD90 0.00166129
R1008 VDD90 VDD90.n187 0.00166129
R1009 VDD90 VDD90.n184 0.00166129
R1010 VDD90.n200 VDD90 0.00166129
R1011 VDD90.n361 VDD90 0.00166129
R1012 VDD90.n357 VDD90 0.00166129
R1013 VDD90.n364 VDD90 0.00166129
R1014 VDD90 VDD90.n14 0.00166129
R1015 VDD90.n80 VDD90 0.00166129
R1016 VDD90.n77 VDD90 0.00166129
R1017 VDD90 VDD90.n74 0.00166129
R1018 VDD90 VDD90.n71 0.00166129
R1019 VDD90 VDD90.n84 0.00166129
R1020 VDD90.n88 VDD90 0.00166129
R1021 VDD90 VDD90.n91 0.00166129
R1022 VDD90.n94 VDD90 0.00166129
R1023 VDD90.n117 VDD90 0.00166129
R1024 VDD90.n114 VDD90 0.00166129
R1025 VDD90 VDD90.n111 0.00166129
R1026 VDD90 VDD90.n108 0.00166129
R1027 VDD90.n122 VDD90 0.00166129
R1028 VDD90 VDD90.n125 0.00166129
R1029 VDD90.n159 VDD90 0.00166129
R1030 VDD90.n48 VDD90.n44 0.001625
R1031 VDD90 VDD90.n242 0.0011
R1032 VDD90.n421 VDD90 0.00108064
R1033 VDD90 VDD90.n424 0.00108064
R1034 VDD90.n441 VDD90 0.00108064
R1035 VDD90.n479 VDD90 0.00108064
R1036 VDD90 VDD90.n482 0.00108064
R1037 VDD90.n295 VDD90 0.00108064
R1038 VDD90.n270 VDD90 0.00108064
R1039 VDD90 VDD90.n273 0.00108064
R1040 VDD90.n325 VDD90 0.00108064
R1041 VDD90 VDD90.n328 0.00108064
R1042 VDD90.n459 VDD90 0.00107692
R1043 VDD90.n349 VDD90 0.00107692
R1044 VDD90.n511 VDD90 0.000799003
R1045 VDD.t9 VDD.n13 765.153
R1046 VDD.t7 VDD.t59 765.152
R1047 VDD.t13 VDD.t15 765.152
R1048 VDD.t11 VDD.t26 765.152
R1049 VDD.t117 VDD.t61 765.152
R1050 VDD.t5 VDD.t67 765.152
R1051 VDD.t73 VDD.t148 763.259
R1052 VDD.t104 VDD.t3 763.259
R1053 VDD.t150 VDD.t153 763.259
R1054 VDD.t181 VDD.t143 763.259
R1055 VDD.t114 VDD.t38 763.259
R1056 VDD.t166 VDD.t129 763.259
R1057 VDD.t107 VDD.t131 763.259
R1058 VDD.t141 VDD.t188 763.259
R1059 VDD.t139 VDD.t171 763.259
R1060 VDD.t40 VDD.t162 763.259
R1061 VDD.t176 VDD.t119 763.259
R1062 VDD.t0 VDD.t145 761.365
R1063 VDD.n23 VDD.t78 759.471
R1064 VDD.n29 VDD.t43 759.471
R1065 VDD.n35 VDD.t22 759.471
R1066 VDD.n39 VDD.t20 759.471
R1067 VDD.t45 VDD.n222 759.471
R1068 VDD.t24 VDD.n220 759.471
R1069 VDD.t50 VDD.n218 759.471
R1070 VDD.t169 VDD.t57 749.85
R1071 VDD.n191 VDD.t76 587.121
R1072 VDD.n224 VDD.t174 505.683
R1073 VDD.n104 VDD.t127 386.348
R1074 VDD.n85 VDD.t186 365.673
R1075 VDD.n112 VDD.t88 365.673
R1076 VDD.n122 VDD.t179 363.185
R1077 VDD.n121 VDD.t63 362.418
R1078 VDD.n104 VDD.t86 362.409
R1079 VDD.n83 VDD.t65 360.012
R1080 VDD.n111 VDD.t90 360.012
R1081 VDD.n85 VDD.n84 322.221
R1082 VDD.n105 VDD.n104 319.75
R1083 VDD.n86 VDD.n85 319.733
R1084 VDD.n123 VDD.n122 319.733
R1085 VDD.n113 VDD.n112 319.733
R1086 VDD.t101 VDD.t9 303.031
R1087 VDD.t83 VDD.t7 303.031
R1088 VDD.t95 VDD.t13 303.031
R1089 VDD.t47 VDD.t11 303.031
R1090 VDD.t98 VDD.t169 303.031
R1091 VDD.t174 VDD.t80 303.031
R1092 VDD.t61 VDD.t92 303.031
R1093 VDD.t67 VDD.t17 303.031
R1094 VDD.n18 VDD.t101 193.183
R1095 VDD.n26 VDD.t83 193.183
R1096 VDD.n34 VDD.t95 193.183
R1097 VDD.n38 VDD.t47 193.183
R1098 VDD.n64 VDD.t123 193.183
R1099 VDD.n67 VDD.t73 193.183
R1100 VDD.n69 VDD.t0 193.183
R1101 VDD.n72 VDD.t104 193.183
R1102 VDD.n74 VDD.t150 193.183
R1103 VDD.n77 VDD.t181 193.183
R1104 VDD.n79 VDD.t114 193.183
R1105 VDD.n169 VDD.t166 193.183
R1106 VDD.n103 VDD.t136 193.183
R1107 VDD.n144 VDD.t133 193.183
R1108 VDD.n145 VDD.t107 193.183
R1109 VDD.n157 VDD.t171 193.183
R1110 VDD.n158 VDD.t40 193.183
R1111 VDD.n159 VDD.t176 193.183
R1112 VDD.n61 VDD.t98 193.183
R1113 VDD.t80 VDD.n223 193.183
R1114 VDD.t92 VDD.n221 193.183
R1115 VDD.t17 VDD.n219 193.183
R1116 VDD.n82 VDD.t112 192.236
R1117 VDD.n120 VDD.t31 192.236
R1118 VDD.n110 VDD.t52 192.236
R1119 VDD.t78 VDD.n18 109.849
R1120 VDD.t43 VDD.n26 109.849
R1121 VDD.t22 VDD.n34 109.849
R1122 VDD.t20 VDD.n38 109.849
R1123 VDD.t148 VDD.n64 109.849
R1124 VDD.t145 VDD.n67 109.849
R1125 VDD.t3 VDD.n69 109.849
R1126 VDD.t153 VDD.n72 109.849
R1127 VDD.t143 VDD.n74 109.849
R1128 VDD.t38 VDD.n77 109.849
R1129 VDD.t129 VDD.n79 109.849
R1130 VDD.n169 VDD.t164 109.849
R1131 VDD.t127 VDD.n103 109.849
R1132 VDD.t131 VDD.n144 109.849
R1133 VDD.n145 VDD.t141 109.849
R1134 VDD.n149 VDD.t139 109.849
R1135 VDD.t162 VDD.n157 109.849
R1136 VDD.t119 VDD.n158 109.849
R1137 VDD.n159 VDD.t160 109.849
R1138 VDD.t76 VDD.n61 109.849
R1139 VDD.n223 VDD.t45 109.849
R1140 VDD.n221 VDD.t24 109.849
R1141 VDD.n219 VDD.t50 109.849
R1142 VDD.n81 VDD.t155 96.5914
R1143 VDD.n117 VDD.t28 96.5914
R1144 VDD.n109 VDD.t54 96.5914
R1145 VDD.t112 VDD.n81 54.9247
R1146 VDD.t31 VDD.n117 54.9247
R1147 VDD.t52 VDD.n109 54.9247
R1148 VDD VDD.n53 27.6957
R1149 VDD.n138 VDD 18.0631
R1150 VDD.n101 VDD 11.7877
R1151 VDD.n13 VDD.n12 8.19491
R1152 VDD.n196 VDD.n192 7.963
R1153 VDD.n233 VDD.n232 6.8813
R1154 VDD.n40 VDD.n39 6.3005
R1155 VDD.n42 VDD.n38 6.3005
R1156 VDD.n45 VDD.n35 6.3005
R1157 VDD.n34 VDD.n33 6.3005
R1158 VDD.n29 VDD.n28 6.3005
R1159 VDD.n26 VDD.n25 6.3005
R1160 VDD.n23 VDD.n22 6.3005
R1161 VDD.n18 VDD.n17 6.3005
R1162 VDD.n160 VDD.n159 6.3005
R1163 VDD.n157 VDD.n156 6.3005
R1164 VDD.n150 VDD.n149 6.3005
R1165 VDD.n146 VDD.n145 6.3005
R1166 VDD.n144 VDD.n143 6.3005
R1167 VDD.n103 VDD.n102 6.3005
R1168 VDD.n188 VDD.n67 6.3005
R1169 VDD.n185 VDD.n69 6.3005
R1170 VDD.n182 VDD.n72 6.3005
R1171 VDD.n179 VDD.n74 6.3005
R1172 VDD.n176 VDD.n77 6.3005
R1173 VDD.n173 VDD.n79 6.3005
R1174 VDD.n170 VDD.n169 6.3005
R1175 VDD.n231 VDD.n64 6.3005
R1176 VDD.n218 VDD.n217 6.3005
R1177 VDD.n219 VDD.n215 6.3005
R1178 VDD.n220 VDD.n210 6.3005
R1179 VDD.n221 VDD.n208 6.3005
R1180 VDD.n222 VDD.n203 6.3005
R1181 VDD.n223 VDD.n201 6.3005
R1182 VDD.n226 VDD.n225 6.3005
R1183 VDD.n225 VDD.n224 6.3005
R1184 VDD.n192 VDD.n190 6.3005
R1185 VDD.n192 VDD.n191 6.3005
R1186 VDD.n234 VDD.n61 6.3005
R1187 VDD.n229 VDD.n228 6.1422
R1188 VDD.n10 VDD.t34 5.28166
R1189 VDD VDD.n93 5.23855
R1190 VDD VDD.n99 5.23855
R1191 VDD.n170 VDD.t165 5.21701
R1192 VDD.n160 VDD.t161 5.21701
R1193 VDD.n40 VDD.t72 5.19258
R1194 VDD.n86 VDD.t187 5.19258
R1195 VDD.n84 VDD.t66 5.19258
R1196 VDD.n217 VDD.t111 5.19258
R1197 VDD.n106 VDD.t87 5.1858
R1198 VDD.n2 VDD.t79 5.17202
R1199 VDD.n20 VDD.t60 5.14855
R1200 VDD.n129 VDD.t180 5.14703
R1201 VDD.n124 VDD.t64 5.14703
R1202 VDD.n136 VDD.t91 5.14703
R1203 VDD.n114 VDD.t89 5.14703
R1204 VDD.n213 VDD.t6 5.14703
R1205 VDD.n206 VDD.t118 5.14703
R1206 VDD.n227 VDD.t37 5.14703
R1207 VDD.n56 VDD.t185 5.14703
R1208 VDD.n236 VDD.t58 5.14703
R1209 VDD.n27 VDD.t16 5.14491
R1210 VDD.n44 VDD.t27 5.14046
R1211 VDD.n232 VDD.n63 5.13751
R1212 VDD.n175 VDD.t39 5.13746
R1213 VDD.n181 VDD.t154 5.13746
R1214 VDD.n187 VDD.t146 5.13746
R1215 VDD.n147 VDD.t142 5.13746
R1216 VDD.n155 VDD.t163 5.13746
R1217 VDD.n41 VDD.t21 5.13287
R1218 VDD.n9 VDD.t23 5.13287
R1219 VDD.n171 VDD.n168 5.13287
R1220 VDD.n174 VDD.n78 5.13287
R1221 VDD.n177 VDD.n76 5.13287
R1222 VDD.n180 VDD.n73 5.13287
R1223 VDD.n183 VDD.n71 5.13287
R1224 VDD.n186 VDD.n68 5.13287
R1225 VDD.n189 VDD.n66 5.13287
R1226 VDD.n107 VDD.n97 5.13287
R1227 VDD.n107 VDD.n98 5.13287
R1228 VDD.n95 VDD.n94 5.13287
R1229 VDD.n148 VDD.n92 5.13287
R1230 VDD.n152 VDD.n90 5.13287
R1231 VDD.n154 VDD.n153 5.13287
R1232 VDD.n134 VDD.n115 5.13287
R1233 VDD.n134 VDD.n116 5.13287
R1234 VDD.n127 VDD.n125 5.13287
R1235 VDD.n127 VDD.n126 5.13287
R1236 VDD.n161 VDD.n89 5.13287
R1237 VDD.n216 VDD.t51 5.13287
R1238 VDD.n209 VDD.t25 5.13287
R1239 VDD.n202 VDD.t46 5.13287
R1240 VDD.n62 VDD.t77 5.13287
R1241 VDD.n24 VDD.t44 5.12141
R1242 VDD.n54 VDD.t184 4.96868
R1243 VDD.n194 VDD.n193 4.5005
R1244 VDD.n196 VDD.n194 4.113
R1245 VDD.n167 VDD.t130 3.91303
R1246 VDD.n75 VDD.t144 3.91303
R1247 VDD.n70 VDD.t4 3.91303
R1248 VDD.n65 VDD.t149 3.91303
R1249 VDD.n91 VDD.t140 3.9128
R1250 VDD.n163 VDD.t120 3.9128
R1251 VDD.n141 VDD.t132 3.91277
R1252 VDD.n141 VDD.n140 3.87701
R1253 VDD.n164 VDD.n163 3.87649
R1254 VDD.n119 VDD.n91 3.87641
R1255 VDD.n167 VDD.n166 3.87623
R1256 VDD.n118 VDD.n75 3.87623
R1257 VDD.n96 VDD.n70 3.87623
R1258 VDD.n100 VDD.n65 3.87523
R1259 VDD.n100 VDD.t128 3.51093
R1260 VDD.n166 VDD.t113 3.51093
R1261 VDD.n118 VDD.t35 3.51093
R1262 VDD.n96 VDD.t126 3.51093
R1263 VDD.n164 VDD.t147 3.51079
R1264 VDD.n140 VDD.t53 3.51063
R1265 VDD.n119 VDD.t32 3.51063
R1266 VDD.n107 VDD.n106 3.45802
R1267 VDD.n109 VDD.n108 3.15287
R1268 VDD.n133 VDD.n117 3.1505
R1269 VDD.n81 VDD.n80 3.1505
R1270 VDD.n197 VDD.n196 3.1505
R1271 VDD.n196 VDD.n195 3.1505
R1272 VDD.n237 VDD.n57 3.1505
R1273 VDD.n60 VDD.n57 3.1505
R1274 VDD.n55 VDD.n54 3.1505
R1275 VDD.n6 VDD.n5 2.88349
R1276 VDD.n43 VDD.n37 2.85787
R1277 VDD.n214 VDD.n212 2.85787
R1278 VDD.n207 VDD.n205 2.85787
R1279 VDD.n200 VDD.n199 2.85787
R1280 VDD.n235 VDD.n59 2.85787
R1281 VDD.n32 VDD.n31 2.85561
R1282 VDD.n16 VDD.n15 2.84433
R1283 VDD.n37 VDD.t12 2.2755
R1284 VDD.n37 VDD.n36 2.2755
R1285 VDD.n31 VDD.t14 2.2755
R1286 VDD.n31 VDD.n30 2.2755
R1287 VDD.n5 VDD.t8 2.2755
R1288 VDD.n5 VDD.n4 2.2755
R1289 VDD.n15 VDD.t10 2.2755
R1290 VDD.n15 VDD.n14 2.2755
R1291 VDD.n212 VDD.t68 2.2755
R1292 VDD.n212 VDD.n211 2.2755
R1293 VDD.n205 VDD.t62 2.2755
R1294 VDD.n205 VDD.n204 2.2755
R1295 VDD.n199 VDD.t175 2.2755
R1296 VDD.n199 VDD.n198 2.2755
R1297 VDD.n59 VDD.t170 2.2755
R1298 VDD.n59 VDD.n58 2.2755
R1299 VDD.t59 VDD.n23 1.89444
R1300 VDD.t15 VDD.n29 1.89444
R1301 VDD.t26 VDD.n35 1.89444
R1302 VDD.n39 VDD.t71 1.89444
R1303 VDD.n195 VDD.t36 1.89444
R1304 VDD.n222 VDD.t117 1.89444
R1305 VDD.n220 VDD.t5 1.89444
R1306 VDD.n218 VDD.t110 1.89444
R1307 VDD.t57 VDD.n60 1.81868
R1308 VDD.n48 VDD.n7 1.41965
R1309 VDD.n49 VDD.n6 1.41813
R1310 VDD.n50 VDD.n3 1.41813
R1311 VDD.n51 VDD.n2 1.41813
R1312 VDD.n52 VDD.n1 1.41813
R1313 VDD.n47 VDD.n46 1.41483
R1314 VDD.n53 VDD.n52 1.41139
R1315 VDD.n47 VDD.n8 1.37847
R1316 VDD.n21 VDD.n20 1.31193
R1317 VDD.n10 VDD.n0 1.09386
R1318 VDD.n83 VDD.n82 0.939698
R1319 VDD.n111 VDD.n110 0.939698
R1320 VDD.n121 VDD.n120 0.93954
R1321 VDD.n11 VDD.n10 0.592429
R1322 VDD.n87 VDD 0.412255
R1323 VDD.n131 VDD 0.412255
R1324 VDD.n131 VDD 0.412255
R1325 VDD.n138 VDD 0.411896
R1326 VDD.n87 VDD 0.411255
R1327 VDD.n165 VDD.n164 0.274239
R1328 VDD.n132 VDD.n119 0.273886
R1329 VDD.n140 VDD.n139 0.273886
R1330 VDD.n166 VDD.n165 0.272927
R1331 VDD.n132 VDD.n118 0.272927
R1332 VDD.n139 VDD.n96 0.272927
R1333 VDD.n101 VDD.n100 0.272927
R1334 VDD.n44 VDD.n43 0.230049
R1335 VDD.n214 VDD.n213 0.230049
R1336 VDD.n207 VDD.n206 0.230049
R1337 VDD.n236 VDD.n235 0.230049
R1338 VDD.n172 VDD.n167 0.22389
R1339 VDD.n178 VDD.n75 0.22389
R1340 VDD.n184 VDD.n70 0.22389
R1341 VDD.n230 VDD.n65 0.22389
R1342 VDD.n151 VDD.n91 0.22353
R1343 VDD.n163 VDD.n162 0.22353
R1344 VDD.n142 VDD.n141 0.223424
R1345 VDD.n226 VDD.n200 0.198938
R1346 VDD.n41 VDD 0.181314
R1347 VDD VDD.n216 0.181314
R1348 VDD VDD.n209 0.181314
R1349 VDD VDD.n202 0.181314
R1350 VDD VDD.n56 0.178278
R1351 VDD.n135 VDD.n114 0.176707
R1352 VDD.n27 VDD.n8 0.168501
R1353 VDD.n19 VDD.n6 0.146598
R1354 VDD.n136 VDD.n135 0.143461
R1355 VDD.n46 VDD 0.141701
R1356 VDD.n148 VDD.n147 0.141016
R1357 VDD.n155 VDD.n154 0.141016
R1358 VDD.n181 VDD.n180 0.141016
R1359 VDD.n175 VDD.n174 0.141016
R1360 VDD.n187 VDD.n186 0.140435
R1361 VDD.n128 VDD.n124 0.139013
R1362 VDD.n129 VDD.n128 0.139013
R1363 VDD.n190 VDD.n62 0.131314
R1364 VDD.n43 VDD 0.106177
R1365 VDD VDD.n32 0.106177
R1366 VDD VDD.n16 0.106177
R1367 VDD.n95 VDD 0.106177
R1368 VDD VDD.n148 0.106177
R1369 VDD VDD.n152 0.106177
R1370 VDD.n154 VDD 0.106177
R1371 VDD.n161 VDD 0.106177
R1372 VDD.n189 VDD 0.106177
R1373 VDD.n186 VDD 0.106177
R1374 VDD.n183 VDD 0.106177
R1375 VDD.n180 VDD 0.106177
R1376 VDD.n177 VDD 0.106177
R1377 VDD.n174 VDD 0.106177
R1378 VDD.n171 VDD 0.106177
R1379 VDD VDD.n214 0.106177
R1380 VDD VDD.n207 0.106177
R1381 VDD VDD.n200 0.106177
R1382 VDD.n235 VDD 0.106177
R1383 VDD.n232 VDD 0.101532
R1384 VDD.n11 VDD.n1 0.0922419
R1385 VDD.n21 VDD.n2 0.082371
R1386 VDD.n24 VDD.n7 0.0807581
R1387 VDD.n143 VDD.n142 0.0800484
R1388 VDD.n147 VDD.n146 0.0800484
R1389 VDD.n151 VDD.n150 0.0800484
R1390 VDD.n162 VDD.n88 0.0800484
R1391 VDD.n102 VDD.n101 0.0800484
R1392 VDD.n231 VDD.n230 0.0800484
R1393 VDD.n188 VDD.n187 0.0800484
R1394 VDD.n185 VDD.n184 0.0800484
R1395 VDD.n182 VDD.n181 0.0800484
R1396 VDD.n179 VDD.n178 0.0800484
R1397 VDD.n173 VDD.n172 0.0800484
R1398 VDD VDD.n41 0.0794677
R1399 VDD VDD.n24 0.0794677
R1400 VDD.n216 VDD 0.0794677
R1401 VDD.n209 VDD 0.0794677
R1402 VDD.n202 VDD 0.0794677
R1403 VDD VDD.n9 0.0788871
R1404 VDD VDD.n155 0.0788871
R1405 VDD VDD.n175 0.0788871
R1406 VDD.n142 VDD 0.0713387
R1407 VDD VDD.n151 0.0713387
R1408 VDD.n162 VDD 0.0713387
R1409 VDD.n184 VDD 0.0713387
R1410 VDD.n178 VDD 0.0713387
R1411 VDD.n172 VDD 0.0713387
R1412 VDD VDD.n233 0.0713387
R1413 VDD VDD.n95 0.0701774
R1414 VDD.n152 VDD 0.0701774
R1415 VDD VDD.n161 0.0701774
R1416 VDD VDD.n189 0.0701774
R1417 VDD VDD.n183 0.0701774
R1418 VDD VDD.n177 0.0701774
R1419 VDD VDD.n171 0.0701774
R1420 VDD.n12 VDD.n11 0.0655323
R1421 VDD.n32 VDD.n8 0.0620484
R1422 VDD VDD.n21 0.0568226
R1423 VDD.n127 VDD 0.0533387
R1424 VDD VDD.n107 0.0533387
R1425 VDD.n134 VDD 0.0513065
R1426 VDD.n190 VDD 0.0505
R1427 VDD.n53 VDD.n0 0.0493889
R1428 VDD.n45 VDD.n44 0.0460556
R1429 VDD.n28 VDD.n27 0.0460556
R1430 VDD.n114 VDD.n113 0.0460556
R1431 VDD.n137 VDD.n136 0.0460556
R1432 VDD.n124 VDD.n123 0.0460556
R1433 VDD.n130 VDD.n129 0.0460556
R1434 VDD.n213 VDD.n210 0.0460556
R1435 VDD.n206 VDD.n203 0.0460556
R1436 VDD.n56 VDD.n55 0.0460556
R1437 VDD.n237 VDD.n236 0.0460556
R1438 VDD.n230 VDD.n229 0.0423064
R1439 VDD.n46 VDD.n9 0.0405645
R1440 VDD.n133 VDD.n132 0.0402742
R1441 VDD.n165 VDD.n80 0.0402742
R1442 VDD.n139 VDD.n108 0.0402742
R1443 VDD.n20 VDD.n19 0.040161
R1444 VDD.n49 VDD.n48 0.0378171
R1445 VDD.n128 VDD.n127 0.0338871
R1446 VDD.n52 VDD.n51 0.0326951
R1447 VDD.n50 VDD.n49 0.0319634
R1448 VDD VDD.n6 0.0318548
R1449 VDD.n135 VDD.n134 0.0318548
R1450 VDD.n227 VDD.n226 0.0316111
R1451 VDD.n51 VDD.n50 0.0312317
R1452 VDD.n229 VDD 0.0295323
R1453 VDD.n228 VDD.n197 0.0266111
R1454 VDD VDD.n2 0.0243065
R1455 VDD.n139 VDD.n138 0.0239437
R1456 VDD.n132 VDD.n131 0.0225645
R1457 VDD.n165 VDD.n87 0.0225645
R1458 VDD VDD.n47 0.0218659
R1459 VDD.n16 VDD.n1 0.0214032
R1460 VDD.n228 VDD.n227 0.0199444
R1461 VDD.n48 VDD 0.0135244
R1462 VDD.n122 VDD.n121 0.00940791
R1463 VDD.n85 VDD.n83 0.00925055
R1464 VDD.n112 VDD.n111 0.00925055
R1465 VDD.n106 VDD.n105 0.00883333
R1466 VDD.n233 VDD.n62 0.00862903
R1467 VDD.n22 VDD.n3 0.00282258
R1468 VDD VDD.n7 0.00272222
R1469 VDD.n19 VDD.n3 0.00202542
R1470 VDD VDD.n42 0.00166129
R1471 VDD.n42 VDD 0.00166129
R1472 VDD.n33 VDD 0.00166129
R1473 VDD.n33 VDD 0.00166129
R1474 VDD.n25 VDD 0.00166129
R1475 VDD.n25 VDD 0.00166129
R1476 VDD.n17 VDD 0.00166129
R1477 VDD.n17 VDD 0.00166129
R1478 VDD VDD.n0 0.00166129
R1479 VDD.n143 VDD 0.00166129
R1480 VDD.n146 VDD 0.00166129
R1481 VDD.n150 VDD 0.00166129
R1482 VDD.n156 VDD 0.00166129
R1483 VDD.n156 VDD 0.00166129
R1484 VDD VDD.n88 0.00166129
R1485 VDD VDD.n160 0.00166129
R1486 VDD.n102 VDD 0.00166129
R1487 VDD VDD.n231 0.00166129
R1488 VDD VDD.n188 0.00166129
R1489 VDD VDD.n185 0.00166129
R1490 VDD VDD.n182 0.00166129
R1491 VDD VDD.n179 0.00166129
R1492 VDD VDD.n176 0.00166129
R1493 VDD.n176 VDD 0.00166129
R1494 VDD VDD.n173 0.00166129
R1495 VDD VDD.n170 0.00166129
R1496 VDD.n215 VDD 0.00166129
R1497 VDD VDD.n215 0.00166129
R1498 VDD.n208 VDD 0.00166129
R1499 VDD VDD.n208 0.00166129
R1500 VDD.n201 VDD 0.00166129
R1501 VDD VDD.n201 0.00166129
R1502 VDD VDD.n234 0.00166129
R1503 VDD.n234 VDD 0.00166129
R1504 VDD.n22 VDD 0.00108064
R1505 VDD.n12 VDD 0.00108064
R1506 VDD VDD.n133 0.00108064
R1507 VDD VDD.n80 0.00108064
R1508 VDD.n108 VDD 0.00108064
R1509 VDD VDD.n40 0.00105556
R1510 VDD VDD.n45 0.00105556
R1511 VDD.n28 VDD 0.00105556
R1512 VDD.n84 VDD 0.00105556
R1513 VDD VDD.n86 0.00105556
R1514 VDD.n113 VDD 0.00105556
R1515 VDD VDD.n137 0.00105556
R1516 VDD.n123 VDD 0.00105556
R1517 VDD VDD.n130 0.00105556
R1518 VDD.n105 VDD 0.00105556
R1519 VDD.n217 VDD 0.00105556
R1520 VDD.n210 VDD 0.00105556
R1521 VDD.n203 VDD 0.00105556
R1522 VDD.n197 VDD 0.00105556
R1523 VDD.n55 VDD 0.00105556
R1524 VDD VDD.n237 0.00105556
R1525 VDD.n13 VDD.t33 0.00101274
R1526 Vdiv.n4 Vdiv.n1 7.10886
R1527 Vdiv Vdiv.n3 3.25199
R1528 Vdiv.n3 Vdiv.t1 2.2755
R1529 Vdiv.n3 Vdiv.n2 2.2755
R1530 Vdiv Vdiv.n0 2.26888
R1531 Vdiv Vdiv.n4 0.0889483
R1532 Vdiv.n4 Vdiv 0.0067069
R1533 RST.n26 RST.t26 37.2596
R1534 RST.n227 RST.t94 37.2596
R1535 RST.n215 RST.t43 37.2596
R1536 RST.n383 RST.t47 37.2596
R1537 RST.n424 RST.t13 37.2596
R1538 RST.n265 RST.t118 37.2595
R1539 RST.n40 RST.t93 37.2594
R1540 RST.n147 RST.t46 37.1991
R1541 RST.n61 RST.t110 37.1991
R1542 RST.n252 RST.t35 37.1988
R1543 RST.n277 RST.t48 37.1988
R1544 RST.n34 RST.t6 36.935
R1545 RST.n21 RST.t29 36.935
R1546 RST.n12 RST.t104 36.935
R1547 RST.n10 RST.t122 36.935
R1548 RST.n16 RST.t53 36.935
R1549 RST.n235 RST.t62 36.935
R1550 RST.n222 RST.t102 36.935
R1551 RST.n188 RST.t36 36.935
R1552 RST.n198 RST.t111 36.935
R1553 RST.n209 RST.t8 36.935
R1554 RST.n184 RST.t107 36.935
R1555 RST.n142 RST.t15 36.935
R1556 RST.n133 RST.t58 36.935
R1557 RST.n138 RST.t54 36.935
R1558 RST.n112 RST.t80 36.935
R1559 RST.n123 RST.t106 36.935
R1560 RST.n151 RST.t69 36.935
R1561 RST.n406 RST.t78 36.935
R1562 RST.n403 RST.t124 36.935
R1563 RST.n390 RST.t68 36.935
R1564 RST.n369 RST.t3 36.935
R1565 RST.n377 RST.t76 36.935
R1566 RST.n385 RST.t121 36.935
R1567 RST.n447 RST.t70 36.935
R1568 RST.n444 RST.t24 36.935
R1569 RST.n431 RST.t63 36.935
R1570 RST.n410 RST.t52 36.935
R1571 RST.n418 RST.t40 36.935
R1572 RST.n426 RST.t103 36.935
R1573 RST.n346 RST.t72 36.935
R1574 RST.n356 RST.t67 36.935
R1575 RST.n336 RST.t4 36.935
R1576 RST.n303 RST.t105 36.935
R1577 RST.n322 RST.t18 36.935
R1578 RST.n320 RST.t5 36.935
R1579 RST.n316 RST.t98 36.935
R1580 RST.n326 RST.t71 36.935
R1581 RST.n247 RST.t55 36.935
R1582 RST.n259 RST.t22 36.935
R1583 RST.n269 RST.t73 36.935
R1584 RST.n291 RST.t97 36.935
R1585 RST.n286 RST.t96 36.935
R1586 RST.n100 RST.t87 36.935
R1587 RST.n53 RST.t23 36.935
R1588 RST.n67 RST.t66 36.935
R1589 RST.n88 RST.t44 36.935
R1590 RST.n77 RST.t34 36.935
R1591 RST.n73 RST.t86 36.935
R1592 RST.n5 RST.t41 36.859
R1593 RST.n397 RST.t21 36.859
R1594 RST.n438 RST.t20 36.859
R1595 RST.n34 RST.t101 18.1962
R1596 RST.n21 RST.t120 18.1962
R1597 RST.n12 RST.t82 18.1962
R1598 RST.n10 RST.t114 18.1962
R1599 RST.n16 RST.t42 18.1962
R1600 RST.n235 RST.t109 18.1962
R1601 RST.n222 RST.t10 18.1962
R1602 RST.n188 RST.t92 18.1962
R1603 RST.n198 RST.t28 18.1962
R1604 RST.n209 RST.t57 18.1962
R1605 RST.n184 RST.t25 18.1962
R1606 RST.n142 RST.t31 18.1962
R1607 RST.n133 RST.t79 18.1962
R1608 RST.n138 RST.t74 18.1962
R1609 RST.n112 RST.t119 18.1962
R1610 RST.n123 RST.t14 18.1962
R1611 RST.n151 RST.t90 18.1962
R1612 RST.n406 RST.t65 18.1962
R1613 RST.n403 RST.t115 18.1962
R1614 RST.n390 RST.t56 18.1962
R1615 RST.n369 RST.t9 18.1962
R1616 RST.n377 RST.t99 18.1962
R1617 RST.n385 RST.t61 18.1962
R1618 RST.n447 RST.t84 18.1962
R1619 RST.n444 RST.t38 18.1962
R1620 RST.n431 RST.t75 18.1962
R1621 RST.n410 RST.t51 18.1962
R1622 RST.n418 RST.t39 18.1962
R1623 RST.n426 RST.t100 18.1962
R1624 RST.n346 RST.t123 18.1962
R1625 RST.n356 RST.t117 18.1962
R1626 RST.n336 RST.t50 18.1962
R1627 RST.n303 RST.t19 18.1962
R1628 RST.n322 RST.t37 18.1962
R1629 RST.n320 RST.t17 18.1962
R1630 RST.n326 RST.t91 18.1962
R1631 RST.n247 RST.t59 18.1962
R1632 RST.n259 RST.t30 18.1962
R1633 RST.n269 RST.t81 18.1962
R1634 RST.n291 RST.t113 18.1962
R1635 RST.n286 RST.t112 18.1962
R1636 RST.n100 RST.t77 18.1962
R1637 RST.n53 RST.t45 18.1962
R1638 RST.n67 RST.t88 18.1962
R1639 RST.n88 RST.t60 18.1962
R1640 RST.n77 RST.t89 18.1962
R1641 RST.n73 RST.t85 18.1962
R1642 RST.n252 RST.t16 17.6613
R1643 RST.n277 RST.t83 17.6613
R1644 RST.n147 RST.t32 17.66
R1645 RST.n61 RST.t2 17.66
R1646 RST.n26 RST.t116 17.5947
R1647 RST.n227 RST.t7 17.5947
R1648 RST.n215 RST.t95 17.5947
R1649 RST.n383 RST.t64 17.5947
R1650 RST.n424 RST.t11 17.5947
R1651 RST.n40 RST.t49 17.594
R1652 RST.n265 RST.t125 17.5939
R1653 RST.n3 RST.t27 17.236
R1654 RST.n395 RST.t12 17.236
R1655 RST.n436 RST.t33 17.236
R1656 RST.n317 RST.t108 16.3712
R1657 RST.n166 RST.n157 11.4652
R1658 RST.n162 RST.n160 9.33985
R1659 RST.n456 RST.n455 9.19662
R1660 RST.n318 RST.n317 8.0005
R1661 RST.n365 RST.n300 7.49317
R1662 RST.n285 RST.n284 7.32578
R1663 RST.n283 RST.n275 7.18787
R1664 RST.n392 RST.n389 6.72677
R1665 RST.n433 RST.n430 6.72677
R1666 RST.n39 RST.n18 6.53894
R1667 RST.n167 RST.n166 6.23435
R1668 RST.n450 RST.n449 6.09745
R1669 RST.n38 RST.n31 6.06869
R1670 RST.n239 RST.n232 6.06869
R1671 RST.n242 RST 5.86652
R1672 RST.n75 RST.n74 5.63344
R1673 RST.n157 RST.n150 5.63145
R1674 RST.n140 RST.n139 5.42044
R1675 RST.n450 RST.n408 5.40234
R1676 RST.n14 RST.n13 5.39891
R1677 RST.n324 RST.n323 5.39866
R1678 RST.n162 RST.n161 5.17836
R1679 RST.n275 RST.n268 4.99277
R1680 RST.n98 RST.n58 4.84685
R1681 RST.n31 RST.n24 4.82595
R1682 RST.n232 RST.n225 4.82595
R1683 RST.n38 RST.n37 4.82279
R1684 RST.n239 RST.n238 4.82279
R1685 RST.n51 RST.n47 4.71142
R1686 RST.n106 RST.n98 4.63847
R1687 RST.n31 RST.n30 4.5933
R1688 RST.n232 RST.n231 4.5933
R1689 RST.n212 RST.n211 4.54165
R1690 RST.n187 RST.n186 4.52648
R1691 RST.n197 RST.n176 4.51211
R1692 RST.n310 RST.n309 4.51211
R1693 RST.n181 RST.n180 4.51168
R1694 RST.n206 RST.n203 4.51163
R1695 RST.n196 RST.n173 4.50514
R1696 RST.n375 RST.n370 4.50173
R1697 RST.n382 RST.n378 4.50173
R1698 RST.n416 RST.n411 4.50173
R1699 RST.n423 RST.n419 4.50173
R1700 RST.n37 RST.n36 4.5005
R1701 RST.n24 RST.n23 4.5005
R1702 RST.n238 RST.n237 4.5005
R1703 RST.n225 RST.n224 4.5005
R1704 RST.n228 RST.n226 4.5005
R1705 RST.n229 RST.n226 4.5005
R1706 RST.n216 RST.n214 4.5005
R1707 RST.n217 RST.n214 4.5005
R1708 RST.n189 RST.n177 4.5005
R1709 RST.n195 RST.n174 4.5005
R1710 RST.n199 RST.n174 4.5005
R1711 RST.n197 RST.n196 4.5005
R1712 RST.n201 RST.n175 4.5005
R1713 RST.n207 RST.n206 4.5005
R1714 RST.n211 RST.n210 4.5005
R1715 RST.n186 RST.n185 4.5005
R1716 RST.n172 RST.n171 4.5005
R1717 RST.n201 RST.n194 4.5005
R1718 RST.n201 RST.n200 4.5005
R1719 RST.n202 RST.n201 4.5005
R1720 RST.n192 RST.n191 4.5005
R1721 RST.n127 RST.n124 4.5005
R1722 RST.n127 RST.n126 4.5005
R1723 RST.n128 RST.n122 4.5005
R1724 RST.n156 RST.n155 4.5005
R1725 RST.n375 RST.n374 4.5005
R1726 RST.n373 RST.n368 4.5005
R1727 RST.n382 RST.n381 4.5005
R1728 RST.n380 RST.n376 4.5005
R1729 RST.n416 RST.n415 4.5005
R1730 RST.n414 RST.n409 4.5005
R1731 RST.n423 RST.n422 4.5005
R1732 RST.n421 RST.n417 4.5005
R1733 RST.n305 RST.n302 4.5005
R1734 RST.n305 RST.n304 4.5005
R1735 RST.n308 RST.n306 4.5005
R1736 RST.n312 RST.n311 4.5005
R1737 RST.n319 RST.n313 4.5005
R1738 RST.n319 RST.n318 4.5005
R1739 RST.n308 RST.n307 4.5005
R1740 RST.n250 RST.n249 4.5005
R1741 RST.n262 RST.n261 4.5005
R1742 RST.n274 RST.n273 4.5005
R1743 RST.n58 RST.n57 4.5005
R1744 RST.n299 RST.n298 4.46212
R1745 RST.n275 RST.n274 4.4249
R1746 RST.n98 RST.n64 4.41239
R1747 RST.n111 RST.n109 4.22115
R1748 RST.n240 RST.n219 4.15909
R1749 RST.n298 RST.n287 3.94094
R1750 RST.n157 RST.n156 3.78663
R1751 RST.n300 RST.n250 3.78663
R1752 RST.n284 RST.n262 3.78663
R1753 RST.n4 RST.n3 3.60685
R1754 RST.n396 RST.n395 3.60685
R1755 RST.n437 RST.n436 3.60685
R1756 RST.n325 RST.n324 3.52872
R1757 RST.n15 RST.n14 3.52872
R1758 RST.n405 RST.n402 3.52872
R1759 RST.n446 RST.n443 3.52872
R1760 RST.n389 RST.n388 3.52872
R1761 RST.n408 RST.n405 3.52872
R1762 RST.n430 RST.n429 3.52872
R1763 RST.n449 RST.n446 3.52872
R1764 RST.n388 RST.n387 3.52813
R1765 RST.n429 RST.n428 3.52813
R1766 RST.n144 RST.n143 3.49993
R1767 RST.n387 RST 3.47503
R1768 RST.n428 RST 3.47503
R1769 RST RST.n325 3.47469
R1770 RST.n402 RST 3.47443
R1771 RST.n443 RST 3.47443
R1772 RST RST.n241 3.37151
R1773 RST.n365 RST.n364 3.35059
R1774 RST.n282 RST 3.33453
R1775 RST.n85 RST.n84 2.96983
R1776 RST.n6 RST.n5 2.88526
R1777 RST.n398 RST.n397 2.88526
R1778 RST.n439 RST.n438 2.88526
R1779 RST.n46 RST.n45 2.8454
R1780 RST.n285 RST.n256 2.8446
R1781 RST.n282 RST.n281 2.8446
R1782 RST.n168 RST.n167 2.80196
R1783 RST.n47 RST.n46 2.4333
R1784 RST.n163 RST 2.27453
R1785 RST.n153 RST.n152 2.25731
R1786 RST.n271 RST.n270 2.25731
R1787 RST.n55 RST.n54 2.25731
R1788 RST.n181 RST.n178 2.25481
R1789 RST.n183 RST.n182 2.2505
R1790 RST.n117 RST.n115 2.2505
R1791 RST.n129 RST.n128 2.2505
R1792 RST.n359 RST.n358 2.2505
R1793 RST.n35 RST.n33 2.25022
R1794 RST.n22 RST.n20 2.25022
R1795 RST.n236 RST.n234 2.25022
R1796 RST.n223 RST.n221 2.25022
R1797 RST.n248 RST.n246 2.25022
R1798 RST.n260 RST.n258 2.25022
R1799 RST.n234 RST.n233 2.2492
R1800 RST.n221 RST.n220 2.2492
R1801 RST.n176 RST.n173 2.24707
R1802 RST.n344 RST.n310 2.24707
R1803 RST.n80 RST.n79 2.24515
R1804 RST.n455 RST.n452 2.24395
R1805 RST.n45 RST.n43 2.24196
R1806 RST.n30 RST.n29 2.24196
R1807 RST.n231 RST.n230 2.24196
R1808 RST.n219 RST.n218 2.24196
R1809 RST.n268 RST.n267 2.24196
R1810 RST.n150 RST.n149 2.24157
R1811 RST.n256 RST.n255 2.24157
R1812 RST.n281 RST.n280 2.24157
R1813 RST.n64 RST.n63 2.24157
R1814 RST.n287 RST.n286 2.15477
R1815 RST.n139 RST.n138 2.15059
R1816 RST.n74 RST.n73 2.1497
R1817 RST.n143 RST.n142 2.14848
R1818 RST.n323 RST.n322 2.13714
R1819 RST.n321 RST.n320 2.13714
R1820 RST.n13 RST.n12 2.13713
R1821 RST.n407 RST.n406 2.13713
R1822 RST.n448 RST.n447 2.13713
R1823 RST.n11 RST.n10 2.13713
R1824 RST.n404 RST.n403 2.13713
R1825 RST.n445 RST.n444 2.13713
R1826 RST.n386 RST.n385 2.13592
R1827 RST.n427 RST.n426 2.13592
R1828 RST.n327 RST.n326 2.1359
R1829 RST.n17 RST.n16 2.1349
R1830 RST.n391 RST.n390 2.1349
R1831 RST.n432 RST.n431 2.1349
R1832 RST.n153 RST.n151 2.12457
R1833 RST.n271 RST.n269 2.12457
R1834 RST.n55 RST.n53 2.12457
R1835 RST.n78 RST.n77 2.12403
R1836 RST.n35 RST.n34 2.12393
R1837 RST.n22 RST.n21 2.12393
R1838 RST.n236 RST.n235 2.12393
R1839 RST.n223 RST.n222 2.12393
R1840 RST.n248 RST.n247 2.12393
R1841 RST.n260 RST.n259 2.12393
R1842 RST.n189 RST.n188 2.12318
R1843 RST.n199 RST.n198 2.12318
R1844 RST.n347 RST.n346 2.12318
R1845 RST.n304 RST.n303 2.12318
R1846 RST.n113 RST.n112 2.1224
R1847 RST.n210 RST.n209 2.12221
R1848 RST.n337 RST.n336 2.12221
R1849 RST.n185 RST.n184 2.12188
R1850 RST.n124 RST.n123 2.12188
R1851 RST.n357 RST.n356 2.12188
R1852 RST.n292 RST.n291 2.12188
R1853 RST.n101 RST.n100 2.12188
R1854 RST.n68 RST.n67 2.12188
R1855 RST.n89 RST.n88 2.12175
R1856 RST.n134 RST.n133 2.1217
R1857 RST.n370 RST.n369 2.12075
R1858 RST.n378 RST.n377 2.12075
R1859 RST.n411 RST.n410 2.12075
R1860 RST.n419 RST.n418 2.12075
R1861 RST.n316 RST.n315 2.12075
R1862 RST.n109 RST.n108 2.08273
R1863 RST.n167 RST.n132 2.06221
R1864 RST.n98 RST.n97 1.97488
R1865 RST.n192 RST.n187 1.90023
R1866 RST.n353 RST.n352 1.90023
R1867 RST.n194 RST.n193 1.88263
R1868 RST.n351 RST.n345 1.88263
R1869 RST.n408 RST.n407 1.8705
R1870 RST.n449 RST.n448 1.8705
R1871 RST.n14 RST.n11 1.87041
R1872 RST.n405 RST.n404 1.87041
R1873 RST.n446 RST.n445 1.87041
R1874 RST.n324 RST.n321 1.8704
R1875 RST.n387 RST.n384 1.8703
R1876 RST.n428 RST.n425 1.8703
R1877 RST.n203 RST.n202 1.86678
R1878 RST.n343 RST.n342 1.86678
R1879 RST.n329 RST 1.83526
R1880 RST.n317 RST.n316 1.8255
R1881 RST RST.n386 1.81628
R1882 RST RST.n427 1.81628
R1883 RST RST.n17 1.81585
R1884 RST.n167 RST.n144 1.79221
R1885 RST.n298 RST.n297 1.78745
R1886 RST.n132 RST.n119 1.78161
R1887 RST.n392 RST.n391 1.76851
R1888 RST.n433 RST.n432 1.76851
R1889 RST.n328 RST.n327 1.76243
R1890 RST.n18 RST.n15 1.75158
R1891 RST.n144 RST.n141 1.72354
R1892 RST.n18 RST 1.72336
R1893 RST.n283 RST.n282 1.66471
R1894 RST.n299 RST.n285 1.57395
R1895 RST.n132 RST.n131 1.53272
R1896 RST.n371 RST.n368 1.51229
R1897 RST.n412 RST.n409 1.51229
R1898 RST.n8 RST.n7 1.51223
R1899 RST.n400 RST.n399 1.51223
R1900 RST.n441 RST.n440 1.51223
R1901 RST.n314 RST.n311 1.51223
R1902 RST.n379 RST.n376 1.51214
R1903 RST.n420 RST.n417 1.51214
R1904 RST.n164 RST.n163 1.50509
R1905 RST.n51 RST.n50 1.50055
R1906 RST.n179 RST.n178 1.5005
R1907 RST.n208 RST.n172 1.5005
R1908 RST.n205 RST.n204 1.5005
R1909 RST.n339 RST.n338 1.5005
R1910 RST.n341 RST.n340 1.5005
R1911 RST.n362 RST.n361 1.5005
R1912 RST.n294 RST.n293 1.5005
R1913 RST.n296 RST.n295 1.5005
R1914 RST.n83 RST.n82 1.5005
R1915 RST.n91 RST.n90 1.5005
R1916 RST.n94 RST.n93 1.5005
R1917 RST.n70 RST.n69 1.5005
R1918 RST.n104 RST.n103 1.5005
R1919 RST.n106 RST.n105 1.49882
R1920 RST.n243 RST.n170 1.49805
R1921 RST.n458 RST.n111 1.49778
R1922 RST.n384 RST.n383 1.43806
R1923 RST.n425 RST.n424 1.43806
R1924 RST.n97 RST.n72 1.4372
R1925 RST.n97 RST.n96 1.42363
R1926 RST.n41 RST.n40 1.42237
R1927 RST.n27 RST.n26 1.42168
R1928 RST.n228 RST.n227 1.42168
R1929 RST.n216 RST.n215 1.42168
R1930 RST.n266 RST.n265 1.42098
R1931 RST.n253 RST.n252 1.41601
R1932 RST.n278 RST.n277 1.41601
R1933 RST.n148 RST.n147 1.41552
R1934 RST.n62 RST.n61 1.41552
R1935 RST.n46 RST.n39 1.19738
R1936 RST.n193 RST.n177 1.13307
R1937 RST.n351 RST.n350 1.13307
R1938 RST.n141 RST.n137 1.1266
R1939 RST.n284 RST.n283 1.12471
R1940 RST.n72 RST.n71 1.12389
R1941 RST.n15 RST.n9 1.12371
R1942 RST.n402 RST.n401 1.12371
R1943 RST.n443 RST.n442 1.12371
R1944 RST.n389 RST.n375 1.12354
R1945 RST.n430 RST.n416 1.12354
R1946 RST.n325 RST.n319 1.1235
R1947 RST.n388 RST.n382 1.1235
R1948 RST.n429 RST.n423 1.1235
R1949 RST.n300 RST.n299 1.08012
R1950 RST.n460 RST.n459 0.968374
R1951 RST.n119 RST.n118 0.940487
R1952 RST.n191 RST.n190 0.898107
R1953 RST.n349 RST.n348 0.898107
R1954 RST.n136 RST.n135 0.898026
R1955 RST.n457 RST.n456 0.851724
R1956 RST.n330 RST.n329 0.839477
R1957 RST.n170 RST.n168 0.805644
R1958 RST.n158 RST 0.723675
R1959 RST.n241 RST.n240 0.668278
R1960 RST.n213 RST.n212 0.643971
R1961 RST.n366 RST.n365 0.633678
R1962 RST.n331 RST.n330 0.627203
R1963 RST.n166 RST.n165 0.473577
R1964 RST.n456 RST.n244 0.407304
R1965 RST.n329 RST.n328 0.388998
R1966 RST.n240 RST.n239 0.309974
R1967 RST.n451 RST.n450 0.284363
R1968 RST.n241 RST.n213 0.136193
R1969 RST.n39 RST.n38 0.118716
R1970 RST RST.n162 0.109973
R1971 RST.n386 RST 0.0704961
R1972 RST.n427 RST 0.0704961
R1973 RST.n17 RST 0.0687763
R1974 RST.n391 RST 0.0687763
R1975 RST.n432 RST 0.0687763
R1976 RST.n327 RST 0.0687763
R1977 RST.n11 RST 0.06755
R1978 RST.n404 RST 0.06755
R1979 RST.n445 RST 0.06755
R1980 RST.n13 RST 0.0675495
R1981 RST.n407 RST 0.0675495
R1982 RST.n448 RST 0.0675495
R1983 RST.n321 RST 0.0675415
R1984 RST.n323 RST 0.0675409
R1985 RST.n384 RST 0.0659998
R1986 RST.n425 RST 0.0659998
R1987 RST.n154 RST 0.0593097
R1988 RST.n272 RST 0.0593097
R1989 RST.n56 RST 0.0593097
R1990 RST.n32 RST 0.0584663
R1991 RST.n19 RST 0.0584663
R1992 RST.n233 RST 0.0584663
R1993 RST.n220 RST 0.0584663
R1994 RST.n245 RST 0.0584663
R1995 RST.n257 RST 0.0584663
R1996 RST.n143 RST 0.0563307
R1997 RST.n139 RST 0.0558741
R1998 RST.n135 RST 0.0553557
R1999 RST.n328 RST 0.0544779
R2000 RST.n190 RST 0.0518307
R2001 RST.n348 RST 0.0518307
R2002 RST RST.n392 0.0484016
R2003 RST RST.n433 0.0484016
R2004 RST.n287 RST 0.0476942
R2005 RST.n74 RST 0.0445432
R2006 RST.n146 RST 0.0410354
R2007 RST.n264 RST 0.0410354
R2008 RST.n60 RST 0.0410354
R2009 RST.n42 RST 0.0394837
R2010 RST.n28 RST 0.0394837
R2011 RST.n1 RST 0.0394837
R2012 RST.n229 RST 0.0394837
R2013 RST.n217 RST 0.0394837
R2014 RST.n393 RST 0.0394837
R2015 RST.n380 RST 0.0394837
R2016 RST.n434 RST 0.0394837
R2017 RST.n421 RST 0.0394837
R2018 RST.n312 RST 0.0394837
R2019 RST.n254 RST 0.0394837
R2020 RST.n279 RST 0.0394837
R2021 RST.n102 RST 0.0394837
R2022 RST.n66 RST 0.0394837
R2023 RST.n372 RST 0.0383947
R2024 RST.n413 RST 0.0383947
R2025 RST.n87 RST 0.0379319
R2026 RST.n43 RST.n42 0.0377414
R2027 RST.n29 RST.n28 0.0377414
R2028 RST.n230 RST.n229 0.0377414
R2029 RST.n218 RST.n217 0.0377414
R2030 RST.n114 RST 0.0377414
R2031 RST.n255 RST.n254 0.0377414
R2032 RST.n280 RST.n279 0.0377414
R2033 RST.n103 RST.n102 0.0377414
R2034 RST.n374 RST.n371 0.0377319
R2035 RST.n415 RST.n412 0.0377319
R2036 RST.n381 RST.n379 0.0377318
R2037 RST.n422 RST.n420 0.0377318
R2038 RST.n7 RST.n2 0.0367013
R2039 RST.n399 RST.n394 0.0367013
R2040 RST.n440 RST.n435 0.0367013
R2041 RST.n314 RST.n313 0.0367013
R2042 RST.n207 RST 0.0363802
R2043 RST.n335 RST 0.0363802
R2044 RST.n183 RST.n180 0.0361897
R2045 RST.n115 RST.n114 0.0361897
R2046 RST.n149 RST.n146 0.0361897
R2047 RST.n358 RST.n355 0.0361897
R2048 RST.n267 RST.n264 0.0361897
R2049 RST.n293 RST.n290 0.0361897
R2050 RST.n63 RST.n60 0.0361897
R2051 RST.n69 RST.n66 0.0361897
R2052 RST.n90 RST.n87 0.0361897
R2053 RST.n297 RST.n296 0.0358571
R2054 RST.n126 RST 0.0348285
R2055 RST.n208 RST.n207 0.0346379
R2056 RST.n338 RST.n335 0.0346379
R2057 RST.n180 RST 0.031725
R2058 RST.n355 RST 0.031725
R2059 RST.n290 RST 0.031725
R2060 RST.n367 RST.n366 0.0311
R2061 RST.n94 RST.n85 0.0305
R2062 RST.n76 RST 0.0301733
R2063 RST.n96 RST.n95 0.0295625
R2064 RST.n37 RST 0.0293
R2065 RST.n24 RST 0.0293
R2066 RST.n238 RST 0.0293
R2067 RST.n225 RST 0.0293
R2068 RST.n156 RST 0.0293
R2069 RST.n250 RST 0.0293
R2070 RST.n262 RST 0.0293
R2071 RST.n274 RST 0.0293
R2072 RST.n58 RST 0.0293
R2073 RST.n104 RST.n99 0.0285519
R2074 RST.n197 RST.n195 0.028431
R2075 RST.n373 RST.n372 0.028431
R2076 RST.n414 RST.n413 0.028431
R2077 RST.n135 RST.n134 0.0275188
R2078 RST.n165 RST.n164 0.0274231
R2079 RST.n108 RST.n107 0.02675
R2080 RST.n117 RST.n116 0.0267025
R2081 RST.n127 RST.n125 0.0255
R2082 RST.n79 RST.n76 0.0253276
R2083 RST.n190 RST.n189 0.0249551
R2084 RST.n348 RST.n347 0.0249551
R2085 RST.n175 RST 0.0239664
R2086 RST.n306 RST 0.0239664
R2087 RST.n50 RST.n48 0.0239404
R2088 RST.n45 RST.n44 0.0238218
R2089 RST.n30 RST.n25 0.0238218
R2090 RST.n231 RST.n226 0.0238218
R2091 RST.n219 RST.n214 0.0238218
R2092 RST.n268 RST.n263 0.0238218
R2093 RST.n91 RST.n86 0.0237584
R2094 RST.n196 RST.n174 0.0236959
R2095 RST.n305 RST.n301 0.0236959
R2096 RST.n121 RST.n120 0.0235
R2097 RST.n150 RST.n145 0.0230258
R2098 RST.n256 RST.n251 0.0230258
R2099 RST.n281 RST.n276 0.0230258
R2100 RST.n64 RST.n59 0.0230258
R2101 RST.n83 RST.n75 0.0221964
R2102 RST.n84 RST.n83 0.0221964
R2103 RST.n295 RST.n288 0.0219286
R2104 RST.n359 RST.n354 0.0218402
R2105 RST.n187 RST.n178 0.0205676
R2106 RST.n364 RST.n363 0.0205676
R2107 RST.n362 RST.n353 0.0205676
R2108 RST.n36 RST.n32 0.0196058
R2109 RST.n23 RST.n19 0.0196058
R2110 RST.n237 RST.n233 0.0196058
R2111 RST.n224 RST.n220 0.0196058
R2112 RST.n249 RST.n245 0.0196058
R2113 RST.n261 RST.n257 0.0196058
R2114 RST.n372 RST 0.0194474
R2115 RST.n413 RST 0.0194474
R2116 RST.n204 RST.n203 0.0193514
R2117 RST.n342 RST.n341 0.0193514
R2118 RST.n155 RST.n154 0.0187743
R2119 RST.n273 RST.n272 0.0187743
R2120 RST.n57 RST.n56 0.0187743
R2121 RST.n206 RST.n205 0.0181289
R2122 RST.n340 RST.n333 0.0181289
R2123 RST.n244 RST.n243 0.01766
R2124 RST.n141 RST.n140 0.0175868
R2125 RST.n51 RST.n0 0.01754
R2126 RST.n452 RST.n451 0.0163335
R2127 RST.n79 RST.n78 0.0160172
R2128 RST.n455 RST.n454 0.0159928
R2129 RST.n202 RST.n173 0.0144865
R2130 RST.n344 RST.n343 0.0144865
R2131 RST.n164 RST.n158 0.0140977
R2132 RST.n201 RST.n176 0.0130264
R2133 RST.n310 RST.n308 0.0130264
R2134 RST.n185 RST.n183 0.0129138
R2135 RST.n358 RST.n357 0.0129138
R2136 RST.n293 RST.n292 0.0129138
R2137 RST.n461 RST.n460 0.01274
R2138 RST.n82 RST.n80 0.0127086
R2139 RST.n70 RST.n65 0.0125591
R2140 RST.n111 RST.n110 0.0120785
R2141 RST.n193 RST.n192 0.0117735
R2142 RST.n352 RST.n351 0.0117735
R2143 RST.n170 RST.n169 0.0116705
R2144 RST.n182 RST.n181 0.0116103
R2145 RST.n107 RST.n106 0.0115492
R2146 RST.n458 RST.n457 0.0107
R2147 RST.n50 RST.n49 0.010313
R2148 RST.n243 RST.n242 0.00992367
R2149 RST.n195 RST.n175 0.00825862
R2150 RST.n200 RST.n199 0.00825862
R2151 RST.n210 RST.n208 0.00825862
R2152 RST.n338 RST.n337 0.00825862
R2153 RST.n90 RST.n89 0.00825862
R2154 RST.n194 RST.n173 0.0077973
R2155 RST.n345 RST.n344 0.0077973
R2156 RST.n459 RST.n458 0.00681423
R2157 RST.n200 RST.n197 0.0067069
R2158 RST.n315 RST.n314 0.00540913
R2159 RST.n294 RST.n289 0.0052523
R2160 RST.n115 RST.n113 0.00515517
R2161 RST.n149 RST.n148 0.00515517
R2162 RST.n267 RST.n266 0.00515517
R2163 RST.n63 RST.n62 0.00515517
R2164 RST.n69 RST.n68 0.00515517
R2165 RST.n7 RST.n6 0.0051456
R2166 RST.n399 RST.n398 0.0051456
R2167 RST.n440 RST.n439 0.0051456
R2168 RST.n211 RST.n172 0.00513918
R2169 RST.n186 RST.n179 0.00513918
R2170 RST.n361 RST.n360 0.00513918
R2171 RST.n339 RST.n334 0.00513918
R2172 RST.n137 RST.n136 0.00494444
R2173 RST.n93 RST.n92 0.00454494
R2174 RST.n379 RST.n378 0.00438036
R2175 RST.n420 RST.n419 0.00438036
R2176 RST.n371 RST.n370 0.00438025
R2177 RST.n412 RST.n411 0.00438025
R2178 RST.n375 RST.n368 0.00391772
R2179 RST.n416 RST.n409 0.00391772
R2180 RST.n9 RST.n8 0.003875
R2181 RST.n401 RST.n400 0.003875
R2182 RST.n382 RST.n376 0.003875
R2183 RST.n442 RST.n441 0.003875
R2184 RST.n423 RST.n417 0.003875
R2185 RST.n319 RST.n311 0.003875
R2186 RST.n118 RST.n117 0.00372575
R2187 RST.n295 RST.n294 0.00371429
R2188 RST.n52 RST.n51 0.00362
R2189 RST.n43 RST.n41 0.00360345
R2190 RST.n29 RST.n27 0.00360345
R2191 RST.n230 RST.n228 0.00360345
R2192 RST.n218 RST.n216 0.00360345
R2193 RST.n255 RST.n253 0.00360345
R2194 RST.n280 RST.n278 0.00360345
R2195 RST.n103 RST.n101 0.00360345
R2196 RST.n71 RST.n70 0.00353371
R2197 RST RST.n461 0.00338
R2198 RST.n155 RST.n153 0.00333412
R2199 RST.n273 RST.n271 0.00333412
R2200 RST.n57 RST.n55 0.00333412
R2201 RST.n191 RST.n177 0.00328351
R2202 RST.n205 RST.n172 0.00328351
R2203 RST.n182 RST.n179 0.00328351
R2204 RST.n350 RST.n349 0.00328351
R2205 RST.n361 RST.n359 0.00328351
R2206 RST.n340 RST.n339 0.00328351
R2207 RST.n105 RST.n104 0.00283766
R2208 RST.n36 RST.n35 0.00255119
R2209 RST.n23 RST.n22 0.00255119
R2210 RST.n237 RST.n236 0.00255119
R2211 RST.n224 RST.n223 0.00255119
R2212 RST.n249 RST.n248 0.00255119
R2213 RST.n261 RST.n260 0.00255119
R2214 RST.n82 RST.n81 0.00245652
R2215 RST RST.n52 0.00242
R2216 RST.n204 RST.n171 0.00232432
R2217 RST.n212 RST.n171 0.00232432
R2218 RST.n363 RST.n362 0.00232432
R2219 RST.n341 RST.n332 0.00232432
R2220 RST.n332 RST.n331 0.00232432
R2221 RST.n163 RST.n159 0.00217441
R2222 RST.n2 RST.n1 0.00205172
R2223 RST.n394 RST.n393 0.00205172
R2224 RST.n374 RST.n373 0.00205172
R2225 RST.n381 RST.n380 0.00205172
R2226 RST.n435 RST.n434 0.00205172
R2227 RST.n415 RST.n414 0.00205172
R2228 RST.n422 RST.n421 0.00205172
R2229 RST.n313 RST.n312 0.00205172
R2230 RST.n6 RST.n4 0.00199457
R2231 RST.n398 RST.n396 0.00199457
R2232 RST.n439 RST.n437 0.00199457
R2233 RST.n318 RST.n315 0.00173095
R2234 RST.n33 RST 0.0017
R2235 RST.n20 RST 0.0017
R2236 RST.n234 RST 0.0017
R2237 RST.n221 RST 0.0017
R2238 RST.n152 RST 0.0017
R2239 RST.n246 RST 0.0017
R2240 RST.n258 RST 0.0017
R2241 RST.n270 RST 0.0017
R2242 RST.n54 RST 0.0017
R2243 RST.n452 RST.n367 0.00158
R2244 RST.n93 RST.n91 0.00151124
R2245 RST.n128 RST.n121 0.0015
R2246 RST.n128 RST.n127 0.0015
R2247 RST.n131 RST.n130 0.0015
R2248 RST.n130 RST.n129 0.0015
R2249 RST.n95 RST.n94 0.0014375
R2250 RST.n201 RST.n174 0.00142783
R2251 RST.n308 RST.n305 0.00142783
R2252 RST.n168 RST 0.00110105
R2253 RST.n109 RST 0.0010568
R2254 RST.n213 RST 0.00104528
R2255 RST.n47 RST 0.00104485
R2256 RST.n330 RST 0.00104041
R2257 RST.n454 RST.n453 0.000945545
R2258 VDD96.n227 VDD96.n226 11185.2
R2259 VDD96.n363 VDD96.n45 2201.41
R2260 VDD96.t235 VDD96.t314 961.905
R2261 VDD96.t233 VDD96.t343 961.905
R2262 VDD96.t139 VDD96.t196 765.152
R2263 VDD96.t270 VDD96.t131 765.152
R2264 VDD96.t308 VDD96.t198 765.152
R2265 VDD96.t136 VDD96.t142 765.152
R2266 VDD96.t272 VDD96.t133 765.152
R2267 VDD96.t329 VDD96.t83 765.152
R2268 VDD96.t89 VDD96.t340 765.152
R2269 VDD96.t190 VDD96.t94 765.152
R2270 VDD96.t97 VDD96.t25 765.152
R2271 VDD96.t105 VDD96.t108 765.152
R2272 VDD96.t13 VDD96.t18 765.152
R2273 VDD96.t368 VDD96.t100 765.152
R2274 VDD96.t248 VDD96.t117 765.152
R2275 VDD96.t264 VDD96.t253 765.152
R2276 VDD96.t41 VDD96.t186 765.152
R2277 VDD96.t212 VDD96.t215 765.152
R2278 VDD96.t276 VDD96.t243 765.152
R2279 VDD96.t220 VDD96.t297 765.152
R2280 VDD96.t0 VDD96.t258 765.152
R2281 VDD96.t204 VDD96.t200 765.152
R2282 VDD96.t81 VDD96.t79 765.152
R2283 VDD96.t261 VDD96.t51 765.152
R2284 VDD96.t202 VDD96.t207 765.152
R2285 VDD96.t58 VDD96.t87 765.152
R2286 VDD96.t238 VDD96.t241 765.152
R2287 VDD96.t304 VDD96.t299 765.152
R2288 VDD96.t319 VDD96.t4 765.152
R2289 VDD96.n226 VDD96.t306 676.191
R2290 VDD96.n227 VDD96.t150 485.714
R2291 VDD96 VDD96.n212 429.187
R2292 VDD96 VDD96.n0 427.092
R2293 VDD96.t225 VDD96.n227 426.44
R2294 VDD96 VDD96.n2 420.935
R2295 VDD96.n212 VDD96.t147 386.365
R2296 VDD96.t343 VDD96.t230 380.952
R2297 VDD96.t362 VDD96.n2 378.788
R2298 VDD96.t360 VDD96.n364 329.546
R2299 VDD96.n364 VDD96.n363 324.075
R2300 VDD96.n2 VDD96.t256 322.223
R2301 VDD96.t313 VDD96.n0 320.635
R2302 VDD96.t294 VDD96.t270 303.031
R2303 VDD96.t68 VDD96.t308 303.031
R2304 VDD96.t73 VDD96.t329 303.031
R2305 VDD96.t340 VDD96.t355 303.031
R2306 VDD96.t286 VDD96.t190 303.031
R2307 VDD96.t291 VDD96.t13 303.031
R2308 VDD96.t62 VDD96.t368 303.031
R2309 VDD96.t117 VDD96.t126 303.031
R2310 VDD96.t284 VDD96.t264 303.031
R2311 VDD96.t278 VDD96.t276 303.031
R2312 VDD96.t110 VDD96.t220 303.031
R2313 VDD96.t79 VDD96.t323 303.031
R2314 VDD96.t280 VDD96.t202 303.031
R2315 VDD96.t316 VDD96.t58 303.031
R2316 VDD96.t288 VDD96.t304 303.031
R2317 VDD96.t222 VDD96.t319 303.031
R2318 VDD96.n226 VDD96.t301 285.714
R2319 VDD96.n218 VDD96.t345 242.857
R2320 VDD96.n219 VDD96.t235 242.857
R2321 VDD96.t301 VDD96.n225 242.857
R2322 VDD96.t230 VDD96.n134 242.857
R2323 VDD96.t128 VDD96.t274 239.583
R2324 VDD96.t267 VDD96.t2 239.583
R2325 VDD96.t22 VDD96.t11 235.35
R2326 VDD96.t193 VDD96.t32 235.35
R2327 VDD96.n4 VDD96.t362 193.183
R2328 VDD96.n14 VDD96.t310 193.183
R2329 VDD96.n16 VDD96.t139 193.183
R2330 VDD96.n19 VDD96.t294 193.183
R2331 VDD96.n22 VDD96.t68 193.183
R2332 VDD96.n37 VDD96.t333 193.183
R2333 VDD96.n38 VDD96.t136 193.183
R2334 VDD96.n44 VDD96.t133 193.183
R2335 VDD96.n365 VDD96.t73 193.183
R2336 VDD96.n121 VDD96.t365 193.183
R2337 VDD96.n123 VDD96.t105 193.183
R2338 VDD96.n126 VDD96.t291 193.183
R2339 VDD96.n129 VDD96.t62 193.183
R2340 VDD96.n305 VDD96.t227 193.183
R2341 VDD96.n307 VDD96.t212 193.183
R2342 VDD96.n310 VDD96.t278 193.183
R2343 VDD96.n313 VDD96.t110 193.183
R2344 VDD96.n199 VDD96.t76 193.183
R2345 VDD96.n205 VDD96.t258 193.183
R2346 VDD96.n206 VDD96.t204 193.183
R2347 VDD96.n211 VDD96.t323 193.183
R2348 VDD96.n173 VDD96.t65 193.183
R2349 VDD96.n175 VDD96.t261 193.183
R2350 VDD96.n178 VDD96.t280 193.183
R2351 VDD96.n181 VDD96.t316 193.183
R2352 VDD96.n140 VDD96.t326 193.183
R2353 VDD96.n142 VDD96.t238 193.183
R2354 VDD96.n145 VDD96.t288 193.183
R2355 VDD96.n148 VDD96.t222 193.183
R2356 VDD96.t355 VDD96.n79 191.288
R2357 VDD96.n80 VDD96.t286 191.288
R2358 VDD96.t25 VDD96.n88 191.288
R2359 VDD96.n89 VDD96.t338 191.288
R2360 VDD96.t126 VDD96.n265 191.288
R2361 VDD96.n266 VDD96.t284 191.288
R2362 VDD96.t186 VDD96.n274 191.288
R2363 VDD96.n275 VDD96.t115 191.288
R2364 VDD96.t38 VDD96.t123 142.993
R2365 VDD96.t209 VDD96.t336 142.993
R2366 VDD96.t120 VDD96.t188 142.993
R2367 VDD96.t113 VDD96.t9 142.993
R2368 VDD96.n1 VDD96.t313 142.857
R2369 VDD96.t350 VDD96.t357 140.465
R2370 VDD96.t102 VDD96.t353 140.465
R2371 VDD96.t53 VDD96.t27 140.465
R2372 VDD96.t60 VDD96.t44 140.465
R2373 VDD96.t314 VDD96.n218 138.095
R2374 VDD96.n219 VDD96.t306 138.095
R2375 VDD96.n225 VDD96.t233 138.095
R2376 VDD96.t150 VDD96.n134 138.095
R2377 VDD96.n364 VDD96.t56 125.001
R2378 VDD96.n79 VDD96.t156 111.743
R2379 VDD96.n80 VDD96.t89 111.743
R2380 VDD96.n88 VDD96.t94 111.743
R2381 VDD96.n89 VDD96.t97 111.743
R2382 VDD96.n265 VDD96.t183 111.743
R2383 VDD96.n266 VDD96.t248 111.743
R2384 VDD96.n274 VDD96.t253 111.743
R2385 VDD96.n275 VDD96.t41 111.743
R2386 VDD96.t256 VDD96.n1 111.112
R2387 VDD96.n4 VDD96.t71 109.849
R2388 VDD96.t196 VDD96.n14 109.849
R2389 VDD96.t131 VDD96.n16 109.849
R2390 VDD96.t198 VDD96.n19 109.849
R2391 VDD96.n22 VDD96.t176 109.849
R2392 VDD96.t142 VDD96.n37 109.849
R2393 VDD96.n38 VDD96.t272 109.849
R2394 VDD96.t83 VDD96.n44 109.849
R2395 VDD96.n365 VDD96.t360 109.849
R2396 VDD96.t108 VDD96.n121 109.849
R2397 VDD96.t18 VDD96.n123 109.849
R2398 VDD96.t100 VDD96.n126 109.849
R2399 VDD96.n129 VDD96.t170 109.849
R2400 VDD96.t215 VDD96.n305 109.849
R2401 VDD96.t243 VDD96.n307 109.849
R2402 VDD96.t297 VDD96.n310 109.849
R2403 VDD96.n313 VDD96.t153 109.849
R2404 VDD96.n199 VDD96.t0 109.849
R2405 VDD96.t200 VDD96.n205 109.849
R2406 VDD96.n206 VDD96.t81 109.849
R2407 VDD96.t147 VDD96.n211 109.849
R2408 VDD96.t51 VDD96.n173 109.849
R2409 VDD96.t207 VDD96.n175 109.849
R2410 VDD96.t87 VDD96.n178 109.849
R2411 VDD96.n181 VDD96.t173 109.849
R2412 VDD96.t241 VDD96.n140 109.849
R2413 VDD96.t299 VDD96.n142 109.849
R2414 VDD96.t4 VDD96.n145 109.849
R2415 VDD96.n148 VDD96.t167 109.849
R2416 VDD96.n230 VDD96.t38 96.5914
R2417 VDD96.n245 VDD96.t120 96.5914
R2418 VDD96.t336 VDD96.n232 95.6444
R2419 VDD96.t9 VDD96.n247 95.6444
R2420 VDD96.n46 VDD96.t350 94.8842
R2421 VDD96.n61 VDD96.t53 94.8842
R2422 VDD96.t353 VDD96.n48 93.954
R2423 VDD96.t44 VDD96.n63 93.954
R2424 VDD96.t179 VDD96.t85 88.0687
R2425 VDD96.n236 VDD96.t6 88.0687
R2426 VDD96.n240 VDD96.t251 88.0687
R2427 VDD96.t217 VDD96.t164 88.0687
R2428 VDD96.t245 VDD96.n238 87.1217
R2429 VDD96.t36 VDD96.n242 87.1217
R2430 VDD96.t160 VDD96.t144 86.5121
R2431 VDD96.n52 VDD96.t46 86.5121
R2432 VDD96.n56 VDD96.t92 86.5121
R2433 VDD96.t29 VDD96.t331 86.5121
R2434 VDD96.t15 VDD96.n54 85.5819
R2435 VDD96.t348 VDD96.n58 85.5819
R2436 VDD96.n212 VDD96.t321 59.702
R2437 VDD96.n0 VDD96.t49 59.4064
R2438 VDD96.n2 VDD96.t34 58.5371
R2439 VDD96.n232 VDD96.t179 55.8717
R2440 VDD96.n238 VDD96.t128 55.8717
R2441 VDD96.n242 VDD96.t267 55.8717
R2442 VDD96.n247 VDD96.t217 55.8717
R2443 VDD96.t85 VDD96.n230 54.9247
R2444 VDD96.t274 VDD96.n236 54.9247
R2445 VDD96.t2 VDD96.n240 54.9247
R2446 VDD96.t164 VDD96.n245 54.9247
R2447 VDD96.n48 VDD96.t160 54.8842
R2448 VDD96.n54 VDD96.t22 54.8842
R2449 VDD96.n58 VDD96.t193 54.8842
R2450 VDD96.n63 VDD96.t29 54.8842
R2451 VDD96.t144 VDD96.n46 53.954
R2452 VDD96.t11 VDD96.n52 53.954
R2453 VDD96.t32 VDD96.n56 53.954
R2454 VDD96.t331 VDD96.n61 53.954
R2455 VDD96.n70 VDD96.t155 30.9379
R2456 VDD96.n72 VDD96.t159 30.9379
R2457 VDD96.n339 VDD96.t175 30.9379
R2458 VDD96.n254 VDD96.t182 30.9379
R2459 VDD96.n256 VDD96.t178 30.9379
R2460 VDD96.n314 VDD96.t163 30.9379
R2461 VDD96.n316 VDD96.t152 30.9379
R2462 VDD96.n183 VDD96.t172 30.9379
R2463 VDD96.n182 VDD96.t146 30.9379
R2464 VDD96.n149 VDD96.t149 30.9379
R2465 VDD96.n150 VDD96.t166 30.9379
R2466 VDD96.n131 VDD96.t169 30.0062
R2467 VDD96.n70 VDD96.t384 24.5101
R2468 VDD96.n72 VDD96.t379 24.5101
R2469 VDD96.n339 VDD96.t371 24.5101
R2470 VDD96.n254 VDD96.t374 24.5101
R2471 VDD96.n256 VDD96.t370 24.5101
R2472 VDD96.n314 VDD96.t372 24.5101
R2473 VDD96.n316 VDD96.t380 24.5101
R2474 VDD96.n183 VDD96.t375 24.5101
R2475 VDD96.n182 VDD96.t385 24.5101
R2476 VDD96.n149 VDD96.t382 24.5101
R2477 VDD96.n150 VDD96.t378 24.5101
R2478 VDD96.n345 VDD96.t377 24.4392
R2479 VDD96 VDD96.t225 10.5649
R2480 VDD96.n377 VDD96.n375 9.16414
R2481 VDD96.t6 VDD96.t209 8.52323
R2482 VDD96.t251 VDD96.t245 8.52323
R2483 VDD96.t188 VDD96.t36 8.52323
R2484 VDD96.t46 VDD96.t102 8.37259
R2485 VDD96.t92 VDD96.t15 8.37259
R2486 VDD96.t27 VDD96.t348 8.37259
R2487 VDD96 VDD96.t113 8.19444
R2488 VDD96 VDD96.t123 8.19444
R2489 VDD96 VDD96.t60 8.16097
R2490 VDD96.n346 VDD96.n345 8.0005
R2491 VDD96.n23 VDD96.n22 6.3005
R2492 VDD96.n26 VDD96.n19 6.3005
R2493 VDD96.n29 VDD96.n16 6.3005
R2494 VDD96.n32 VDD96.n14 6.3005
R2495 VDD96.n79 VDD96.n78 6.3005
R2496 VDD96.n81 VDD96.n80 6.3005
R2497 VDD96.n88 VDD96.n87 6.3005
R2498 VDD96.n90 VDD96.n89 6.3005
R2499 VDD96.n112 VDD96.n48 6.3005
R2500 VDD96.n106 VDD96.n54 6.3005
R2501 VDD96.n100 VDD96.n58 6.3005
R2502 VDD96.n94 VDD96.n63 6.3005
R2503 VDD96.n97 VDD96.n61 6.3005
R2504 VDD96.n103 VDD96.n56 6.3005
R2505 VDD96.n109 VDD96.n52 6.3005
R2506 VDD96.n115 VDD96.n46 6.3005
R2507 VDD96 VDD96.n45 6.3005
R2508 VDD96.n265 VDD96.n264 6.3005
R2509 VDD96.n267 VDD96.n266 6.3005
R2510 VDD96.n274 VDD96.n273 6.3005
R2511 VDD96.n276 VDD96.n275 6.3005
R2512 VDD96.n298 VDD96.n232 6.3005
R2513 VDD96.n292 VDD96.n238 6.3005
R2514 VDD96.n286 VDD96.n242 6.3005
R2515 VDD96.n280 VDD96.n247 6.3005
R2516 VDD96.n283 VDD96.n245 6.3005
R2517 VDD96.n289 VDD96.n240 6.3005
R2518 VDD96.n295 VDD96.n236 6.3005
R2519 VDD96.n301 VDD96.n230 6.3005
R2520 VDD96.n322 VDD96.n313 6.3005
R2521 VDD96.n325 VDD96.n310 6.3005
R2522 VDD96.n328 VDD96.n307 6.3005
R2523 VDD96.n331 VDD96.n305 6.3005
R2524 VDD96.n187 VDD96.n181 6.3005
R2525 VDD96.n190 VDD96.n178 6.3005
R2526 VDD96.n193 VDD96.n175 6.3005
R2527 VDD96.n196 VDD96.n173 6.3005
R2528 VDD96.n200 VDD96.n199 6.3005
R2529 VDD96.n205 VDD96.n204 6.3005
R2530 VDD96.n207 VDD96.n206 6.3005
R2531 VDD96.n211 VDD96.n210 6.3005
R2532 VDD96.n154 VDD96.n148 6.3005
R2533 VDD96.n157 VDD96.n145 6.3005
R2534 VDD96.n160 VDD96.n142 6.3005
R2535 VDD96.n163 VDD96.n140 6.3005
R2536 VDD96.n336 VDD96.n134 6.3005
R2537 VDD96.n218 VDD96.n217 6.3005
R2538 VDD96.n220 VDD96.n219 6.3005
R2539 VDD96.n225 VDD96.n224 6.3005
R2540 VDD96.n350 VDD96.n129 6.3005
R2541 VDD96.n353 VDD96.n126 6.3005
R2542 VDD96.n356 VDD96.n123 6.3005
R2543 VDD96.n359 VDD96.n121 6.3005
R2544 VDD96.n363 VDD96 6.3005
R2545 VDD96.n44 VDD96.n43 6.3005
R2546 VDD96.n39 VDD96.n38 6.3005
R2547 VDD96.n37 VDD96.n36 6.3005
R2548 VDD96.n366 VDD96.n365 6.3005
R2549 VDD96.n369 VDD96.n4 6.3005
R2550 VDD96.n373 VDD96.n1 6.3005
R2551 VDD96.n341 VDD96.n340 5.63356
R2552 VDD96 VDD96.n377 5.233
R2553 VDD96.n23 VDD96.t177 5.213
R2554 VDD96.n119 VDD96.n118 5.19407
R2555 VDD96.n117 VDD96.n116 5.19167
R2556 VDD96.n42 VDD96.t84 5.13287
R2557 VDD96.n41 VDD96.n9 5.13287
R2558 VDD96.n40 VDD96.t273 5.13287
R2559 VDD96.n11 VDD96.n10 5.13287
R2560 VDD96.n35 VDD96.t143 5.13287
R2561 VDD96.n34 VDD96.n12 5.13287
R2562 VDD96.n25 VDD96.t199 5.13287
R2563 VDD96.n28 VDD96.t132 5.13287
R2564 VDD96.n30 VDD96.n15 5.13287
R2565 VDD96.n31 VDD96.t197 5.13287
R2566 VDD96.n33 VDD96.n13 5.13287
R2567 VDD96.n74 VDD96.n69 5.13287
R2568 VDD96.n68 VDD96.n67 5.13287
R2569 VDD96.n83 VDD96.n64 5.13287
R2570 VDD96.n86 VDD96.t26 5.13287
R2571 VDD96.n85 VDD96.n84 5.13287
R2572 VDD96.n91 VDD96.t339 5.13287
R2573 VDD96.n92 VDD96.t45 5.13287
R2574 VDD96.n114 VDD96.n47 5.13287
R2575 VDD96.n107 VDD96.n53 5.13287
R2576 VDD96.n104 VDD96.t93 5.13287
R2577 VDD96.n101 VDD96.n57 5.13287
R2578 VDD96.n98 VDD96.t28 5.13287
R2579 VDD96.n96 VDD96.n62 5.13287
R2580 VDD96.n95 VDD96.t332 5.13287
R2581 VDD96.n102 VDD96.t33 5.13287
R2582 VDD96.n105 VDD96.n55 5.13287
R2583 VDD96.n108 VDD96.t12 5.13287
R2584 VDD96.n111 VDD96.n49 5.13287
R2585 VDD96.n113 VDD96.t145 5.13287
R2586 VDD96.n260 VDD96.n253 5.13287
R2587 VDD96.n252 VDD96.n251 5.13287
R2588 VDD96.n269 VDD96.n248 5.13287
R2589 VDD96.n272 VDD96.t187 5.13287
R2590 VDD96.n271 VDD96.n270 5.13287
R2591 VDD96.n277 VDD96.t116 5.13287
R2592 VDD96.n321 VDD96.t154 5.13287
R2593 VDD96.n324 VDD96.t298 5.13287
R2594 VDD96.n327 VDD96.t244 5.13287
R2595 VDD96.n329 VDD96.n306 5.13287
R2596 VDD96.n330 VDD96.t216 5.13287
R2597 VDD96.n332 VDD96.n304 5.13287
R2598 VDD96.n165 VDD96.t148 5.13287
R2599 VDD96.n208 VDD96.t82 5.13287
R2600 VDD96.n169 VDD96.n168 5.13287
R2601 VDD96.n203 VDD96.t201 5.13287
R2602 VDD96.n202 VDD96.n170 5.13287
R2603 VDD96.n201 VDD96.t1 5.13287
R2604 VDD96.n198 VDD96.n171 5.13287
R2605 VDD96.n186 VDD96.t174 5.13287
R2606 VDD96.n189 VDD96.t88 5.13287
R2607 VDD96.n192 VDD96.t208 5.13287
R2608 VDD96.n194 VDD96.n174 5.13287
R2609 VDD96.n195 VDD96.t52 5.13287
R2610 VDD96.n197 VDD96.n172 5.13287
R2611 VDD96.n153 VDD96.t168 5.13287
R2612 VDD96.n156 VDD96.t5 5.13287
R2613 VDD96.n159 VDD96.t300 5.13287
R2614 VDD96.n161 VDD96.n141 5.13287
R2615 VDD96.n162 VDD96.t242 5.13287
R2616 VDD96.n164 VDD96.n139 5.13287
R2617 VDD96.n335 VDD96.t151 5.13287
R2618 VDD96.n223 VDD96.t234 5.13287
R2619 VDD96.n222 VDD96.n135 5.13287
R2620 VDD96.n221 VDD96.t307 5.13287
R2621 VDD96.n137 VDD96.n136 5.13287
R2622 VDD96.n216 VDD96.t315 5.13287
R2623 VDD96.n215 VDD96.n138 5.13287
R2624 VDD96.n352 VDD96.t101 5.13287
R2625 VDD96.n355 VDD96.t19 5.13287
R2626 VDD96.n357 VDD96.n122 5.13287
R2627 VDD96.n358 VDD96.t109 5.13287
R2628 VDD96.n360 VDD96.n120 5.13287
R2629 VDD96.n5 VDD96.t361 5.13287
R2630 VDD96.n368 VDD96.t72 5.13287
R2631 VDD96.n370 VDD96.n3 5.13287
R2632 VDD96 VDD96.n376 5.118
R2633 VDD96.n300 VDD96.n231 5.11708
R2634 VDD96.n293 VDD96.n237 5.11708
R2635 VDD96.n290 VDD96.t252 5.11708
R2636 VDD96.n287 VDD96.n241 5.11708
R2637 VDD96.n284 VDD96.t189 5.11708
R2638 VDD96.n282 VDD96.n246 5.11708
R2639 VDD96.n279 VDD96.t10 5.11708
R2640 VDD96.n281 VDD96.t165 5.1155
R2641 VDD96.n288 VDD96.t3 5.1155
R2642 VDD96.n291 VDD96.n239 5.1155
R2643 VDD96.n294 VDD96.t275 5.1155
R2644 VDD96.n297 VDD96.n233 5.1155
R2645 VDD96.n299 VDD96.t86 5.1155
R2646 VDD96.n302 VDD96.n229 5.1155
R2647 VDD96 VDD96.t61 5.10312
R2648 VDD96.n303 VDD96.n228 5.09407
R2649 VDD96.n334 VDD96.t226 5.09407
R2650 VDD96.n213 VDD96.t322 5.09407
R2651 VDD96.n371 VDD96.t35 5.09407
R2652 VDD96.n374 VDD96.t50 5.09407
R2653 VDD96.n278 VDD96.t114 5.09264
R2654 VDD96.n362 VDD96.t57 5.09264
R2655 VDD96.n349 VDD96.t171 4.8755
R2656 VDD96.n342 VDD96.n130 4.51383
R2657 VDD96.n345 VDD96.n344 4.5005
R2658 VDD96.n372 VDD96.t257 4.12326
R2659 VDD96.n257 VDD96.n256 4.08796
R2660 VDD96 VDD96.n149 4.08442
R2661 VDD96.n184 VDD96.n183 4.08323
R2662 VDD96.n71 VDD96.n70 4.07925
R2663 VDD96.n151 VDD96.n150 4.07855
R2664 VDD96.n255 VDD96.n254 4.07362
R2665 VDD96.n315 VDD96.n314 4.04647
R2666 VDD96 VDD96.n72 4.04611
R2667 VDD96 VDD96.n182 4.04234
R2668 VDD96.n317 VDD96.n316 4.041
R2669 VDD96.n343 VDD96.n131 3.61662
R2670 VDD96.n259 VDD96.n258 3.13455
R2671 VDD96.n320 VDD96.n315 3.01689
R2672 VDD96.n73 VDD96 3.01101
R2673 VDD96.n152 VDD96 2.99823
R2674 VDD96.n185 VDD96 2.9975
R2675 VDD96.n259 VDD96.n255 2.95902
R2676 VDD96.n73 VDD96.n71 2.91542
R2677 VDD96.n185 VDD96.n184 2.87793
R2678 VDD96.n152 VDD96.n151 2.86761
R2679 VDD96.n8 VDD96.n7 2.85787
R2680 VDD96.n24 VDD96.n21 2.85787
R2681 VDD96.n27 VDD96.n18 2.85787
R2682 VDD96.n77 VDD96.n76 2.85787
R2683 VDD96.n82 VDD96.n66 2.85787
R2684 VDD96.n110 VDD96.n51 2.85787
R2685 VDD96.n99 VDD96.n60 2.85787
R2686 VDD96.n263 VDD96.n262 2.85787
R2687 VDD96.n268 VDD96.n250 2.85787
R2688 VDD96.n323 VDD96.n312 2.85787
R2689 VDD96.n326 VDD96.n309 2.85787
R2690 VDD96.n209 VDD96.n167 2.85787
R2691 VDD96.n188 VDD96.n180 2.85787
R2692 VDD96.n191 VDD96.n177 2.85787
R2693 VDD96.n155 VDD96.n147 2.85787
R2694 VDD96.n158 VDD96.n144 2.85787
R2695 VDD96.n337 VDD96.n133 2.85787
R2696 VDD96.n351 VDD96.n128 2.85787
R2697 VDD96.n354 VDD96.n125 2.85787
R2698 VDD96.n320 VDD96.n319 2.84443
R2699 VDD96.n296 VDD96.n235 2.84208
R2700 VDD96.n285 VDD96.n244 2.8405
R2701 VDD96.n341 VDD96.n338 2.65604
R2702 VDD96.n7 VDD96.t330 2.2755
R2703 VDD96.n7 VDD96.n6 2.2755
R2704 VDD96.n21 VDD96.t309 2.2755
R2705 VDD96.n21 VDD96.n20 2.2755
R2706 VDD96.n18 VDD96.t271 2.2755
R2707 VDD96.n18 VDD96.n17 2.2755
R2708 VDD96.n76 VDD96.t356 2.2755
R2709 VDD96.n76 VDD96.n75 2.2755
R2710 VDD96.n66 VDD96.t287 2.2755
R2711 VDD96.n66 VDD96.n65 2.2755
R2712 VDD96.n51 VDD96.t354 2.2755
R2713 VDD96.n51 VDD96.n50 2.2755
R2714 VDD96.n60 VDD96.t349 2.2755
R2715 VDD96.n60 VDD96.n59 2.2755
R2716 VDD96.n235 VDD96.t337 2.2755
R2717 VDD96.n235 VDD96.n234 2.2755
R2718 VDD96.n262 VDD96.t127 2.2755
R2719 VDD96.n262 VDD96.n261 2.2755
R2720 VDD96.n250 VDD96.t285 2.2755
R2721 VDD96.n250 VDD96.n249 2.2755
R2722 VDD96.n244 VDD96.t37 2.2755
R2723 VDD96.n244 VDD96.n243 2.2755
R2724 VDD96.n312 VDD96.t221 2.2755
R2725 VDD96.n312 VDD96.n311 2.2755
R2726 VDD96.n309 VDD96.t277 2.2755
R2727 VDD96.n309 VDD96.n308 2.2755
R2728 VDD96.n167 VDD96.t80 2.2755
R2729 VDD96.n167 VDD96.n166 2.2755
R2730 VDD96.n180 VDD96.t59 2.2755
R2731 VDD96.n180 VDD96.n179 2.2755
R2732 VDD96.n177 VDD96.t203 2.2755
R2733 VDD96.n177 VDD96.n176 2.2755
R2734 VDD96.n147 VDD96.t320 2.2755
R2735 VDD96.n147 VDD96.n146 2.2755
R2736 VDD96.n144 VDD96.t305 2.2755
R2737 VDD96.n144 VDD96.n143 2.2755
R2738 VDD96.n133 VDD96.t344 2.2755
R2739 VDD96.n133 VDD96.n132 2.2755
R2740 VDD96.n128 VDD96.t369 2.2755
R2741 VDD96.n128 VDD96.n127 2.2755
R2742 VDD96.n125 VDD96.t14 2.2755
R2743 VDD96.n125 VDD96.n124 2.2755
R2744 VDD96.n321 VDD96.n320 2.26792
R2745 VDD96.n74 VDD96.n73 2.26734
R2746 VDD96.n153 VDD96.n152 2.26618
R2747 VDD96.n186 VDD96.n185 2.2656
R2748 VDD96.n260 VDD96.n259 2.26502
R2749 VDD96.n340 VDD96.n339 2.11318
R2750 VDD96.t357 VDD96.n45 1.86097
R2751 VDD96.n344 VDD96.n342 1.54785
R2752 VDD96.n342 VDD96.n341 1.35532
R2753 VDD96.n34 VDD96.n33 1.16167
R2754 VDD96.n198 VDD96.n197 1.16167
R2755 VDD96.n361 VDD96.n360 1.06836
R2756 VDD96.n333 VDD96.n332 1.04079
R2757 VDD96.n278 VDD96.n277 1.03836
R2758 VDD96.n214 VDD96.n164 1.02405
R2759 VDD96.n92 VDD96.n91 0.993021
R2760 VDD96.n345 VDD96.n131 0.840632
R2761 VDD96.n257 VDD96 0.533317
R2762 VDD96 VDD96.n367 0.468962
R2763 VDD96.n350 VDD96.n349 0.337997
R2764 VDD96.n349 VDD96.n348 0.328132
R2765 VDD96.n368 VDD96 0.243482
R2766 VDD96.n28 VDD96.n27 0.233919
R2767 VDD96.n25 VDD96.n24 0.233919
R2768 VDD96.n77 VDD96.n68 0.233919
R2769 VDD96.n83 VDD96.n82 0.233919
R2770 VDD96.n263 VDD96.n252 0.233919
R2771 VDD96.n269 VDD96.n268 0.233919
R2772 VDD96.n327 VDD96.n326 0.233919
R2773 VDD96.n324 VDD96.n323 0.233919
R2774 VDD96.n192 VDD96.n191 0.233919
R2775 VDD96.n189 VDD96.n188 0.233919
R2776 VDD96.n159 VDD96.n158 0.233919
R2777 VDD96.n156 VDD96.n155 0.233919
R2778 VDD96.n355 VDD96.n354 0.233919
R2779 VDD96.n352 VDD96.n351 0.233919
R2780 VDD96.n334 VDD96.n333 0.211434
R2781 VDD96.n335 VDD96 0.182611
R2782 VDD96 VDD96.n165 0.179233
R2783 VDD96 VDD96.n5 0.17738
R2784 VDD96.n374 VDD96.n373 0.16404
R2785 VDD96.n333 VDD96.n303 0.158852
R2786 VDD96.n214 VDD96.n213 0.152441
R2787 VDD96.n372 VDD96 0.147753
R2788 VDD96.n377 VDD96 0.144879
R2789 VDD96.n31 VDD96.n30 0.141016
R2790 VDD96.n86 VDD96.n85 0.141016
R2791 VDD96.n272 VDD96.n271 0.141016
R2792 VDD96.n330 VDD96.n329 0.141016
R2793 VDD96.n195 VDD96.n194 0.141016
R2794 VDD96.n202 VDD96.n201 0.141016
R2795 VDD96.n203 VDD96.n169 0.141016
R2796 VDD96.n162 VDD96.n161 0.141016
R2797 VDD96.n216 VDD96.n137 0.141016
R2798 VDD96.n222 VDD96.n221 0.141016
R2799 VDD96.n358 VDD96.n357 0.141016
R2800 VDD96.n35 VDD96.n11 0.141016
R2801 VDD96.n41 VDD96.n40 0.141016
R2802 VDD96.n215 VDD96.n214 0.131304
R2803 VDD96 VDD96.n208 0.122435
R2804 VDD96.n223 VDD96 0.122435
R2805 VDD96.n42 VDD96 0.122435
R2806 VDD96.n209 VDD96 0.111984
R2807 VDD96 VDD96.n8 0.111984
R2808 VDD96.n33 VDD96.n32 0.107339
R2809 VDD96.n30 VDD96.n29 0.107339
R2810 VDD96.n87 VDD96.n86 0.107339
R2811 VDD96.n91 VDD96.n90 0.107339
R2812 VDD96.n273 VDD96.n272 0.107339
R2813 VDD96.n277 VDD96.n276 0.107339
R2814 VDD96.n332 VDD96.n331 0.107339
R2815 VDD96.n329 VDD96.n328 0.107339
R2816 VDD96.n197 VDD96.n196 0.107339
R2817 VDD96.n194 VDD96.n193 0.107339
R2818 VDD96.n200 VDD96.n198 0.107339
R2819 VDD96.n204 VDD96.n202 0.107339
R2820 VDD96.n207 VDD96.n169 0.107339
R2821 VDD96.n164 VDD96.n163 0.107339
R2822 VDD96.n161 VDD96.n160 0.107339
R2823 VDD96.n217 VDD96.n215 0.107339
R2824 VDD96.n220 VDD96.n137 0.107339
R2825 VDD96.n224 VDD96.n222 0.107339
R2826 VDD96.n360 VDD96.n359 0.107339
R2827 VDD96.n357 VDD96.n356 0.107339
R2828 VDD96.n36 VDD96.n34 0.107339
R2829 VDD96.n39 VDD96.n11 0.107339
R2830 VDD96.n43 VDD96.n41 0.107339
R2831 VDD96.n371 VDD96.n370 0.10725
R2832 VDD96.n340 VDD96 0.106795
R2833 VDD96 VDD96.n77 0.106758
R2834 VDD96.n82 VDD96 0.106758
R2835 VDD96 VDD96.n263 0.106758
R2836 VDD96.n268 VDD96 0.106758
R2837 VDD96.n27 VDD96 0.106177
R2838 VDD96.n24 VDD96 0.106177
R2839 VDD96.n326 VDD96 0.106177
R2840 VDD96.n323 VDD96 0.106177
R2841 VDD96.n191 VDD96 0.106177
R2842 VDD96.n188 VDD96 0.106177
R2843 VDD96 VDD96.n209 0.106177
R2844 VDD96.n158 VDD96 0.106177
R2845 VDD96.n155 VDD96 0.106177
R2846 VDD96.n337 VDD96 0.106177
R2847 VDD96.n354 VDD96 0.106177
R2848 VDD96.n351 VDD96 0.106177
R2849 VDD96.n317 VDD96 0.102091
R2850 VDD96.n370 VDD96.n369 0.0854231
R2851 VDD96.n362 VDD96.n361 0.0852977
R2852 VDD96.n338 VDD96.n337 0.0846936
R2853 VDD96.n26 VDD96.n25 0.080629
R2854 VDD96.n78 VDD96.n74 0.080629
R2855 VDD96.n81 VDD96.n68 0.080629
R2856 VDD96.n264 VDD96.n260 0.080629
R2857 VDD96.n267 VDD96.n252 0.080629
R2858 VDD96.n325 VDD96.n324 0.080629
R2859 VDD96.n322 VDD96.n321 0.080629
R2860 VDD96.n190 VDD96.n189 0.080629
R2861 VDD96.n187 VDD96.n186 0.080629
R2862 VDD96.n210 VDD96.n165 0.080629
R2863 VDD96.n157 VDD96.n156 0.080629
R2864 VDD96.n154 VDD96.n153 0.080629
R2865 VDD96.n336 VDD96.n335 0.080629
R2866 VDD96.n353 VDD96.n352 0.080629
R2867 VDD96 VDD96.n31 0.0794677
R2868 VDD96 VDD96.n28 0.0794677
R2869 VDD96 VDD96.n330 0.0794677
R2870 VDD96 VDD96.n327 0.0794677
R2871 VDD96 VDD96.n195 0.0794677
R2872 VDD96 VDD96.n192 0.0794677
R2873 VDD96.n201 VDD96 0.0794677
R2874 VDD96 VDD96.n203 0.0794677
R2875 VDD96.n208 VDD96 0.0794677
R2876 VDD96 VDD96.n162 0.0794677
R2877 VDD96 VDD96.n159 0.0794677
R2878 VDD96 VDD96.n216 0.0794677
R2879 VDD96.n221 VDD96 0.0794677
R2880 VDD96 VDD96.n223 0.0794677
R2881 VDD96 VDD96.n358 0.0794677
R2882 VDD96 VDD96.n355 0.0794677
R2883 VDD96 VDD96.n35 0.0794677
R2884 VDD96.n40 VDD96 0.0794677
R2885 VDD96 VDD96.n42 0.0794677
R2886 VDD96 VDD96.n83 0.0788871
R2887 VDD96.n85 VDD96 0.0788871
R2888 VDD96 VDD96.n269 0.0788871
R2889 VDD96.n271 VDD96 0.0788871
R2890 VDD96.n347 VDD96 0.0733571
R2891 VDD96 VDD96.n372 0.0674231
R2892 VDD96 VDD96.n368 0.0605
R2893 VDD96.n367 VDD96.n5 0.0562419
R2894 VDD96.n361 VDD96.n119 0.0557941
R2895 VDD96.n302 VDD96.n301 0.0505302
R2896 VDD96.n280 VDD96.n279 0.0505302
R2897 VDD96.n105 VDD96.n104 0.0480988
R2898 VDD96.n291 VDD96.n290 0.0478112
R2899 VDD96.n348 VDD96.n347 0.0471071
R2900 VDD96.n110 VDD96.n109 0.0470046
R2901 VDD96.n100 VDD96.n99 0.0470046
R2902 VDD96.n119 VDD96 0.046755
R2903 VDD96 VDD96.n111 0.046731
R2904 VDD96.n296 VDD96.n295 0.0467236
R2905 VDD96.n286 VDD96.n285 0.0467236
R2906 VDD96.n98 VDD96 0.0464574
R2907 VDD96 VDD96.n297 0.0464517
R2908 VDD96.n284 VDD96 0.0461798
R2909 VDD96 VDD96.n334 0.0457727
R2910 VDD96.n213 VDD96 0.0444412
R2911 VDD96 VDD96.n362 0.0438334
R2912 VDD96.n367 VDD96.n8 0.0411452
R2913 VDD96 VDD96.n102 0.0377036
R2914 VDD96 VDD96.n288 0.0374789
R2915 VDD96.n107 VDD96 0.0374301
R2916 VDD96.n293 VDD96 0.0372069
R2917 VDD96 VDD96.n371 0.036939
R2918 VDD96.n346 VDD96.n130 0.0358571
R2919 VDD96.n348 VDD96.n346 0.03425
R2920 VDD96 VDD96.n92 0.0327059
R2921 VDD96 VDD96.n108 0.0325061
R2922 VDD96 VDD96.n294 0.0323127
R2923 VDD96.n101 VDD96 0.0322325
R2924 VDD96.n287 VDD96 0.0320408
R2925 VDD96.n93 VDD96 0.0298382
R2926 VDD96.n338 VDD96 0.0277903
R2927 VDD96.n108 VDD96.n107 0.0262143
R2928 VDD96.n102 VDD96.n101 0.0262143
R2929 VDD96.n294 VDD96.n293 0.0260589
R2930 VDD96.n288 VDD96.n287 0.0260589
R2931 VDD96 VDD96.n278 0.023068
R2932 VDD96.n303 VDD96 0.0227961
R2933 VDD96 VDD96.n374 0.0209098
R2934 VDD96.n113 VDD96.n112 0.020196
R2935 VDD96.n97 VDD96.n96 0.020196
R2936 VDD96.n367 VDD96.n366 0.0201154
R2937 VDD96.n299 VDD96.n298 0.020077
R2938 VDD96.n283 VDD96.n282 0.020077
R2939 VDD96 VDD96.n302 0.0198051
R2940 VDD96 VDD96.n114 0.0196489
R2941 VDD96 VDD96.n300 0.0195332
R2942 VDD96.n279 VDD96 0.0195332
R2943 VDD96.n95 VDD96 0.0193754
R2944 VDD96.n281 VDD96 0.0192613
R2945 VDD96.n114 VDD96.n113 0.0185547
R2946 VDD96.n96 VDD96.n95 0.0185547
R2947 VDD96.n300 VDD96.n299 0.0184456
R2948 VDD96.n282 VDD96.n281 0.0184456
R2949 VDD96.n117 VDD96.n115 0.0144514
R2950 VDD96.n94 VDD96.n93 0.0141778
R2951 VDD96.n319 VDD96.n318 0.0141364
R2952 VDD96.n255 VDD96 0.012875
R2953 VDD96.n258 VDD96 0.00810563
R2954 VDD96.n71 VDD96 0.00725
R2955 VDD96.n318 VDD96.n317 0.00725
R2956 VDD96.n319 VDD96 0.00595455
R2957 VDD96.n318 VDD96 0.00595455
R2958 VDD96.n184 VDD96 0.00543151
R2959 VDD96.n347 VDD96 0.00478571
R2960 VDD96.n93 VDD96 0.00469118
R2961 VDD96.n111 VDD96.n110 0.00432979
R2962 VDD96.n99 VDD96.n98 0.00432979
R2963 VDD96.n297 VDD96.n296 0.00430665
R2964 VDD96.n285 VDD96.n284 0.00430665
R2965 VDD96.n369 VDD96 0.00419231
R2966 VDD96.n373 VDD96 0.00373077
R2967 VDD96.n343 VDD96.n130 0.00371429
R2968 VDD96.n106 VDD96.n105 0.00323556
R2969 VDD96.n104 VDD96.n103 0.00323556
R2970 VDD96.n292 VDD96.n291 0.00321903
R2971 VDD96.n290 VDD96.n289 0.00321903
R2972 VDD96.n151 VDD96 0.00256897
R2973 VDD96.n119 VDD96.n117 0.00229283
R2974 VDD96.n87 VDD96 0.00224194
R2975 VDD96.n90 VDD96 0.00224194
R2976 VDD96.n273 VDD96 0.00224194
R2977 VDD96.n276 VDD96 0.00224194
R2978 VDD96.n344 VDD96.n343 0.00210714
R2979 VDD96.n258 VDD96.n257 0.00176761
R2980 VDD96.n32 VDD96 0.00166129
R2981 VDD96.n29 VDD96 0.00166129
R2982 VDD96 VDD96.n26 0.00166129
R2983 VDD96 VDD96.n23 0.00166129
R2984 VDD96.n331 VDD96 0.00166129
R2985 VDD96.n328 VDD96 0.00166129
R2986 VDD96 VDD96.n325 0.00166129
R2987 VDD96 VDD96.n322 0.00166129
R2988 VDD96.n196 VDD96 0.00166129
R2989 VDD96.n193 VDD96 0.00166129
R2990 VDD96 VDD96.n190 0.00166129
R2991 VDD96 VDD96.n187 0.00166129
R2992 VDD96 VDD96.n200 0.00166129
R2993 VDD96.n204 VDD96 0.00166129
R2994 VDD96 VDD96.n207 0.00166129
R2995 VDD96.n210 VDD96 0.00166129
R2996 VDD96.n163 VDD96 0.00166129
R2997 VDD96.n160 VDD96 0.00166129
R2998 VDD96 VDD96.n157 0.00166129
R2999 VDD96 VDD96.n154 0.00166129
R3000 VDD96.n217 VDD96 0.00166129
R3001 VDD96 VDD96.n220 0.00166129
R3002 VDD96.n224 VDD96 0.00166129
R3003 VDD96 VDD96.n336 0.00166129
R3004 VDD96.n359 VDD96 0.00166129
R3005 VDD96.n356 VDD96 0.00166129
R3006 VDD96 VDD96.n353 0.00166129
R3007 VDD96 VDD96.n350 0.00166129
R3008 VDD96.n36 VDD96 0.00166129
R3009 VDD96 VDD96.n39 0.00166129
R3010 VDD96.n43 VDD96 0.00166129
R3011 VDD96.n315 VDD96 0.00152273
R3012 VDD96 VDD96.n106 0.00132067
R3013 VDD96 VDD96.n100 0.00132067
R3014 VDD96 VDD96.n94 0.00132067
R3015 VDD96 VDD96.n292 0.00131571
R3016 VDD96 VDD96.n286 0.00131571
R3017 VDD96 VDD96.n280 0.00131571
R3018 VDD96.n78 VDD96 0.00108064
R3019 VDD96 VDD96.n81 0.00108064
R3020 VDD96.n264 VDD96 0.00108064
R3021 VDD96 VDD96.n267 0.00108064
R3022 VDD96.n366 VDD96 0.00107692
R3023 VDD96.n115 VDD96 0.00104711
R3024 VDD96.n109 VDD96 0.00104711
R3025 VDD96.n103 VDD96 0.00104711
R3026 VDD96 VDD96.n97 0.00104711
R3027 VDD96.n301 VDD96 0.00104381
R3028 VDD96.n295 VDD96 0.00104381
R3029 VDD96.n289 VDD96 0.00104381
R3030 VDD96 VDD96.n283 0.00104381
R3031 VDD96.n112 VDD96 0.000773556
R3032 VDD96.n298 VDD96 0.000771903
R3033 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.n3 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.t9 40.2519
R3034 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.n0 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.t3 36.935
R3035 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.n4 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.t4 31.528
R3036 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.n1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.t8 31.528
R3037 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.n0 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.t7 18.1962
R3038 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.n3 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.t5 15.3826
R3039 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.n4 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.t6 15.3826
R3040 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.n1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.t2 15.3826
R3041 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.n4 7.63442
R3042 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.n1 6.86134
R3043 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.n2 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 5.01116
R3044 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.n5 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 3.11241
R3045 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.n6 2.25871
R3046 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.n0 2.13398
R3047 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.n3 2.12278
R3048 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.n5 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 2.10026
R3049 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.n6 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.n2 1.37588
R3050 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.n6 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.n5 1.26898
R3051 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.n2 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 1.12056
R3052 VDD93.n454 VDD93.t343 13882.6
R3053 VDD93.n120 VDD93.t45 13882.6
R3054 VDD93.n451 VDD93.t433 12382.6
R3055 VDD93.n108 VDD93.t127 12382.6
R3056 VDD93.n225 VDD93.n224 11185.2
R3057 VDD93.n446 VDD93.t133 7208.33
R3058 VDD93.n97 VDD93.t327 7041.67
R3059 VDD93.t197 VDD93.t232 961.905
R3060 VDD93.t163 VDD93.t341 961.905
R3061 VDD93.t358 VDD93.n93 848.615
R3062 VDD93.t427 VDD93.n94 809.492
R3063 VDD93.t419 VDD93.t131 765.152
R3064 VDD93.t307 VDD93.t337 765.152
R3065 VDD93.t32 VDD93.t425 765.152
R3066 VDD93.t437 VDD93.t422 765.152
R3067 VDD93.t309 VDD93.t334 765.152
R3068 VDD93.t189 VDD93.t63 765.152
R3069 VDD93.t157 VDD93.t16 765.152
R3070 VDD93.t366 VDD93.t362 765.152
R3071 VDD93.t8 VDD93.t315 765.152
R3072 VDD93.t331 VDD93.t324 765.152
R3073 VDD93.t352 VDD93.t122 765.152
R3074 VDD93.t355 VDD93.t345 765.152
R3075 VDD93.t319 VDD93.t282 765.152
R3076 VDD93.t349 VDD93.t124 765.152
R3077 VDD93.t191 VDD93.t347 765.152
R3078 VDD93.t382 VDD93.t236 765.152
R3079 VDD93.t259 VDD93.t265 765.152
R3080 VDD93.t291 VDD93.t385 765.152
R3081 VDD93.t18 VDD93.t458 765.152
R3082 VDD93.t256 VDD93.t262 765.152
R3083 VDD93.t389 VDD93.t387 765.152
R3084 VDD93.t194 VDD93.t226 765.152
R3085 VDD93.t228 VDD93.t168 765.152
R3086 VDD93.t149 VDD93.t61 765.152
R3087 VDD93.t154 VDD93.t250 765.152
R3088 VDD93.t364 VDD93.t369 765.152
R3089 VDD93.t444 VDD93.t313 765.152
R3090 VDD93.t411 VDD93.t129 765.152
R3091 VDD93.t296 VDD93.t56 765.152
R3092 VDD93.t118 VDD93.t120 765.152
R3093 VDD93.t187 VDD93.t223 765.152
R3094 VDD93.t51 VDD93.t47 765.152
R3095 VDD93.t339 VDD93.t242 765.152
R3096 VDD93.t220 VDD93.t377 765.152
R3097 VDD93.t49 VDD93.t54 765.152
R3098 VDD93.t371 VDD93.t311 765.152
R3099 VDD93.n224 VDD93.t230 676.191
R3100 VDD93.t5 VDD93.t254 536.798
R3101 VDD93.t379 VDD93.t430 501.002
R3102 VDD93.t26 VDD93.t13 501.002
R3103 VDD93.t185 VDD93.t175 501.002
R3104 VDD93.n225 VDD93.t95 485.714
R3105 VDD93.n473 VDD93.t244 485.714
R3106 VDD93 VDD93.n454 451.327
R3107 VDD93.n120 VDD93 448.709
R3108 VDD93 VDD93.n451 445.577
R3109 VDD93.n108 VDD93 442.993
R3110 VDD93 VDD93.n446 431.3
R3111 VDD93 VDD93.n175 429.187
R3112 VDD93.n340 VDD93 429.187
R3113 VDD93.n492 VDD93 429.187
R3114 VDD93 VDD93.n97 428.8
R3115 VDD93.n434 VDD93 427.092
R3116 VDD93.n508 VDD93 427.092
R3117 VDD93 VDD93.n154 426.699
R3118 VDD93 VDD93.n203 426.699
R3119 VDD93.t300 VDD93.n225 426.44
R3120 VDD93.t205 VDD93.n473 426.44
R3121 VDD93 VDD93.n440 425.019
R3122 VDD93 VDD93.n510 420.935
R3123 VDD93.t74 VDD93.n340 386.365
R3124 VDD93.n175 VDD93.t81 386.365
R3125 VDD93.t84 VDD93.n154 386.365
R3126 VDD93.t91 VDD93.n203 386.365
R3127 VDD93.t110 VDD93.n492 386.365
R3128 VDD93.t302 VDD93.t163 380.952
R3129 VDD93.t210 VDD93.t170 380.952
R3130 VDD93.n440 VDD93.t461 378.788
R3131 VDD93.n446 VDD93.t141 378.788
R3132 VDD93.t285 VDD93.n451 378.788
R3133 VDD93.t449 VDD93.n454 378.788
R3134 VDD93.t446 VDD93.n97 378.788
R3135 VDD93.t144 VDD93.n108 378.788
R3136 VDD93.t34 VDD93.n120 378.788
R3137 VDD93.n382 VDD93.t178 362.8
R3138 VDD93.n384 VDD93.t294 362.8
R3139 VDD93.n386 VDD93.t21 359.49
R3140 VDD93.n354 VDD93.t200 359.49
R3141 VDD93.n510 VDD93.t246 322.223
R3142 VDD93.t373 VDD93.n508 320.635
R3143 VDD93.t381 VDD93.n434 309.341
R3144 VDD93.t400 VDD93.t307 303.031
R3145 VDD93.t452 VDD93.t32 303.031
R3146 VDD93.t63 VDD93.t439 303.031
R3147 VDD93.t151 VDD93.t8 303.031
R3148 VDD93.t324 VDD93.t469 303.031
R3149 VDD93.t282 VDD93.t464 303.031
R3150 VDD93.t392 VDD93.t349 303.031
R3151 VDD93.t236 VDD93.t269 303.031
R3152 VDD93.t458 VDD93.t275 303.031
R3153 VDD93.t409 VDD93.t256 303.031
R3154 VDD93.t406 VDD93.t228 303.031
R3155 VDD93.t455 VDD93.t149 303.031
R3156 VDD93.t397 VDD93.t364 303.031
R3157 VDD93.t138 VDD93.t444 303.031
R3158 VDD93.t394 VDD93.t296 303.031
R3159 VDD93.t217 VDD93.t118 303.031
R3160 VDD93.t242 VDD93.t202 303.031
R3161 VDD93.t403 VDD93.t49 303.031
R3162 VDD93.t207 VDD93.t371 303.031
R3163 VDD93.n355 VDD93.t2 296.538
R3164 VDD93.n224 VDD93.t165 285.714
R3165 VDD93.t58 VDD93.n84 285.714
R3166 VDD93.n206 VDD93.t160 242.857
R3167 VDD93.n212 VDD93.t197 242.857
R3168 VDD93.t165 VDD93.n216 242.857
R3169 VDD93.n221 VDD93.t302 242.857
R3170 VDD93.n78 VDD93.t172 242.857
R3171 VDD93.n81 VDD93.t414 242.857
R3172 VDD93.n85 VDD93.t58 242.857
R3173 VDD93.n88 VDD93.t210 242.857
R3174 VDD93.t183 VDD93.n356 227.456
R3175 VDD93.n445 VDD93.t461 193.183
R3176 VDD93.n450 VDD93.t141 193.183
R3177 VDD93.n453 VDD93.t285 193.183
R3178 VDD93.n456 VDD93.t449 193.183
R3179 VDD93.n395 VDD93.t37 193.183
R3180 VDD93.n397 VDD93.t419 193.183
R3181 VDD93.n400 VDD93.t400 193.183
R3182 VDD93.n403 VDD93.t452 193.183
R3183 VDD93.n96 VDD93.t427 193.183
R3184 VDD93.n99 VDD93.t446 193.183
R3185 VDD93.n114 VDD93.t144 193.183
R3186 VDD93.n121 VDD93.t34 193.183
R3187 VDD93.n344 VDD93.t65 193.183
R3188 VDD93.t422 VDD93.n343 193.183
R3189 VDD93.t334 VDD93.n342 193.183
R3190 VDD93.t439 VDD93.n341 193.183
R3191 VDD93.n157 VDD93.t10 193.183
R3192 VDD93.n163 VDD93.t157 193.183
R3193 VDD93.n167 VDD93.t366 193.183
R3194 VDD93.n172 VDD93.t151 193.183
R3195 VDD93.n177 VDD93.t135 193.183
R3196 VDD93.n179 VDD93.t194 193.183
R3197 VDD93.n182 VDD93.t406 193.183
R3198 VDD93.n185 VDD93.t455 193.183
R3199 VDD93.n128 VDD93.t288 193.183
R3200 VDD93.n130 VDD93.t154 193.183
R3201 VDD93.n133 VDD93.t397 193.183
R3202 VDD93.n136 VDD93.t138 193.183
R3203 VDD93.n4 VDD93.t115 193.183
R3204 VDD93.n45 VDD93.t112 193.183
R3205 VDD93.n47 VDD93.t411 193.183
R3206 VDD93.n50 VDD93.t394 193.183
R3207 VDD93.n53 VDD93.t217 193.183
R3208 VDD93.n34 VDD93.t239 193.183
R3209 VDD93.n40 VDD93.t223 193.183
R3210 VDD93.n494 VDD93.t51 193.183
R3211 VDD93.t202 VDD93.n493 193.183
R3212 VDD93.n13 VDD93.t374 193.183
R3213 VDD93.n15 VDD93.t220 193.183
R3214 VDD93.n18 VDD93.t403 193.183
R3215 VDD93.n21 VDD93.t207 193.183
R3216 VDD93.t469 VDD93.n159 191.288
R3217 VDD93.t122 VDD93.n166 191.288
R3218 VDD93.t345 VDD93.n169 191.288
R3219 VDD93.n174 VDD93.t322 191.288
R3220 VDD93.t464 VDD93.n298 191.288
R3221 VDD93.n299 VDD93.t392 191.288
R3222 VDD93.t347 VDD93.n307 191.288
R3223 VDD93.n308 VDD93.t271 191.288
R3224 VDD93.t269 VDD93.n208 191.288
R3225 VDD93.t265 VDD93.n215 191.288
R3226 VDD93.t385 VDD93.n218 191.288
R3227 VDD93.n223 VDD93.t234 191.288
R3228 VDD93.t275 VDD93.n242 191.288
R3229 VDD93.n243 VDD93.t409 191.288
R3230 VDD93.t387 VDD93.n251 191.288
R3231 VDD93.n252 VDD93.t305 191.288
R3232 VDD93.n382 VDD93.n356 167.588
R3233 VDD93.n509 VDD93.t373 142.857
R3234 VDD93.t232 VDD93.n206 138.095
R3235 VDD93.t230 VDD93.n212 138.095
R3236 VDD93.t341 VDD93.n216 138.095
R3237 VDD93.t95 VDD93.n221 138.095
R3238 VDD93.n78 VDD93.t417 138.095
R3239 VDD93.n81 VDD93.t298 138.095
R3240 VDD93.n85 VDD93.t24 138.095
R3241 VDD93.t244 VDD93.n88 138.095
R3242 VDD93.n435 VDD93.t381 137.826
R3243 VDD93.n385 VDD93.n384 119.706
R3244 VDD93.n386 VDD93.n385 118.614
R3245 VDD93.n159 VDD93.t84 111.743
R3246 VDD93.n166 VDD93.t331 111.743
R3247 VDD93.n169 VDD93.t352 111.743
R3248 VDD93.n174 VDD93.t355 111.743
R3249 VDD93.n298 VDD93.t107 111.743
R3250 VDD93.n299 VDD93.t319 111.743
R3251 VDD93.n307 VDD93.t124 111.743
R3252 VDD93.n308 VDD93.t191 111.743
R3253 VDD93.n208 VDD93.t91 111.743
R3254 VDD93.n215 VDD93.t382 111.743
R3255 VDD93.n218 VDD93.t259 111.743
R3256 VDD93.n223 VDD93.t291 111.743
R3257 VDD93.n242 VDD93.t77 111.743
R3258 VDD93.n243 VDD93.t18 111.743
R3259 VDD93.n251 VDD93.t262 111.743
R3260 VDD93.n252 VDD93.t389 111.743
R3261 VDD93.t246 VDD93.n509 111.112
R3262 VDD93.t133 VDD93.n445 109.849
R3263 VDD93.t433 VDD93.n450 109.849
R3264 VDD93.t343 VDD93.n453 109.849
R3265 VDD93.n456 VDD93.t277 109.849
R3266 VDD93.t131 VDD93.n395 109.849
R3267 VDD93.t337 VDD93.n397 109.849
R3268 VDD93.t425 VDD93.n400 109.849
R3269 VDD93.n403 VDD93.t104 109.849
R3270 VDD93.t327 VDD93.n96 109.849
R3271 VDD93.t127 VDD93.n99 109.849
R3272 VDD93.t45 VDD93.n114 109.849
R3273 VDD93.n121 VDD93.t273 109.849
R3274 VDD93.n344 VDD93.t437 109.849
R3275 VDD93.n343 VDD93.t309 109.849
R3276 VDD93.n342 VDD93.t189 109.849
R3277 VDD93.n341 VDD93.t74 109.849
R3278 VDD93.t16 VDD93.n157 109.849
R3279 VDD93.t362 VDD93.n163 109.849
R3280 VDD93.t315 VDD93.n167 109.849
R3281 VDD93.t81 VDD93.n172 109.849
R3282 VDD93.t226 VDD93.n177 109.849
R3283 VDD93.t168 VDD93.n179 109.849
R3284 VDD93.t61 VDD93.n182 109.849
R3285 VDD93.n185 VDD93.t71 109.849
R3286 VDD93.t250 VDD93.n128 109.849
R3287 VDD93.t369 VDD93.n130 109.849
R3288 VDD93.t313 VDD93.n133 109.849
R3289 VDD93.n136 VDD93.t98 109.849
R3290 VDD93.n4 VDD93.t213 109.849
R3291 VDD93.t129 VDD93.n45 109.849
R3292 VDD93.t56 VDD93.n47 109.849
R3293 VDD93.t120 VDD93.n50 109.849
R3294 VDD93.n53 VDD93.t88 109.849
R3295 VDD93.n34 VDD93.t187 109.849
R3296 VDD93.t47 VDD93.n40 109.849
R3297 VDD93.n494 VDD93.t339 109.849
R3298 VDD93.n493 VDD93.t110 109.849
R3299 VDD93.t377 VDD93.n13 109.849
R3300 VDD93.t54 VDD93.n15 109.849
R3301 VDD93.t311 VDD93.n18 109.849
R3302 VDD93.n21 VDD93.t101 109.849
R3303 VDD93.n435 VDD93.t30 107.198
R3304 VDD93.n355 VDD93.n354 100.365
R3305 VDD93.n120 VDD93.t43 65.4455
R3306 VDD93.n108 VDD93.t329 64.6
R3307 VDD93.n454 VDD93.t0 62.8277
R3308 VDD93.n97 VDD93.t68 62.5005
R3309 VDD93.n154 VDD93.t466 62.1896
R3310 VDD93.n203 VDD93.t279 62.1896
R3311 VDD93.n451 VDD93.t267 62.016
R3312 VDD93.n446 VDD93.t435 60.0005
R3313 VDD93.n340 VDD93.t442 59.702
R3314 VDD93.n175 VDD93.t147 59.702
R3315 VDD93.n492 VDD93.t215 59.702
R3316 VDD93.n434 VDD93.t471 59.4064
R3317 VDD93.n508 VDD93.t317 59.4064
R3318 VDD93.n440 VDD93.t181 59.1138
R3319 VDD93.n510 VDD93.t248 58.5371
R3320 VDD93.n385 VDD93.n356 47.8826
R3321 VDD93.n406 VDD93.t103 30.9379
R3322 VDD93.n404 VDD93.t73 30.9379
R3323 VDD93.n288 VDD93.t106 30.9379
R3324 VDD93.n290 VDD93.t83 30.9379
R3325 VDD93.n232 VDD93.t76 30.9379
R3326 VDD93.n233 VDD93.t90 30.9379
R3327 VDD93.n186 VDD93.t94 30.9379
R3328 VDD93.n188 VDD93.t70 30.9379
R3329 VDD93.n137 VDD93.t80 30.9379
R3330 VDD93.n139 VDD93.t97 30.9379
R3331 VDD93.n54 VDD93.t100 30.9379
R3332 VDD93.n59 VDD93.t87 30.0062
R3333 VDD93.n391 VDD93.t2 28.139
R3334 VDD93.t254 VDD93.n391 28.139
R3335 VDD93.n392 VDD93.t5 28.139
R3336 VDD93.n392 VDD93.t252 28.139
R3337 VDD93.n406 VDD93.t474 24.5101
R3338 VDD93.n404 VDD93.t484 24.5101
R3339 VDD93.n288 VDD93.t483 24.5101
R3340 VDD93.n290 VDD93.t478 24.5101
R3341 VDD93.n232 VDD93.t480 24.5101
R3342 VDD93.n233 VDD93.t476 24.5101
R3343 VDD93.n186 VDD93.t477 24.5101
R3344 VDD93.n188 VDD93.t485 24.5101
R3345 VDD93.n137 VDD93.t481 24.5101
R3346 VDD93.n139 VDD93.t475 24.5101
R3347 VDD93.n54 VDD93.t487 24.5101
R3348 VDD93.n58 VDD93.t486 24.4392
R3349 VDD93.n367 VDD93.t40 22.0446
R3350 VDD93.n368 VDD93.t379 22.0446
R3351 VDD93.n371 VDD93.t430 22.0446
R3352 VDD93.n372 VDD93.t26 22.0446
R3353 VDD93.n375 VDD93.t13 22.0446
R3354 VDD93.n376 VDD93.t185 22.0446
R3355 VDD93.n379 VDD93.t175 21.0426
R3356 VDD93.n380 VDD93.t183 21.0426
R3357 VDD93.n385 VDD93.n355 18.2487
R3358 VDD93 VDD93.t300 10.5649
R3359 VDD93 VDD93.t205 10.5649
R3360 VDD93.n364 VDD93.t380 8.94586
R3361 VDD93.n362 VDD93.t27 8.94586
R3362 VDD93.n360 VDD93.t186 8.94586
R3363 VDD93.n358 VDD93.t184 8.92336
R3364 VDD93.n56 VDD93.n55 6.98838
R3365 VDD93.n117 VDD93.t44 6.62407
R3366 VDD93.n470 VDD93.n468 6.57033
R3367 VDD93.n457 VDD93.n456 6.3005
R3368 VDD93.n461 VDD93.n453 6.3005
R3369 VDD93.n450 VDD93.n449 6.3005
R3370 VDD93.n445 VDD93.n444 6.3005
R3371 VDD93.n367 VDD93 6.3005
R3372 VDD93 VDD93.n368 6.3005
R3373 VDD93.n371 VDD93 6.3005
R3374 VDD93 VDD93.n372 6.3005
R3375 VDD93.n375 VDD93 6.3005
R3376 VDD93 VDD93.n376 6.3005
R3377 VDD93.n379 VDD93 6.3005
R3378 VDD93 VDD93.n380 6.3005
R3379 VDD93.n384 VDD93 6.3005
R3380 VDD93 VDD93.n382 6.3005
R3381 VDD93.n419 VDD93.n395 6.3005
R3382 VDD93.n416 VDD93.n397 6.3005
R3383 VDD93.n413 VDD93.n400 6.3005
R3384 VDD93.n410 VDD93.n403 6.3005
R3385 VDD93.n242 VDD93.n241 6.3005
R3386 VDD93.n244 VDD93.n243 6.3005
R3387 VDD93.n251 VDD93.n250 6.3005
R3388 VDD93.n253 VDD93.n252 6.3005
R3389 VDD93.n192 VDD93.n185 6.3005
R3390 VDD93.n195 VDD93.n182 6.3005
R3391 VDD93.n198 VDD93.n179 6.3005
R3392 VDD93.n201 VDD93.n177 6.3005
R3393 VDD93.n275 VDD93.n208 6.3005
R3394 VDD93.n268 VDD93.n215 6.3005
R3395 VDD93.n263 VDD93.n218 6.3005
R3396 VDD93.n257 VDD93.n223 6.3005
R3397 VDD93.n260 VDD93.n221 6.3005
R3398 VDD93.n267 VDD93.n216 6.3005
R3399 VDD93.n272 VDD93.n212 6.3005
R3400 VDD93.n278 VDD93.n206 6.3005
R3401 VDD93.n298 VDD93.n297 6.3005
R3402 VDD93.n300 VDD93.n299 6.3005
R3403 VDD93.n307 VDD93.n306 6.3005
R3404 VDD93.n309 VDD93.n308 6.3005
R3405 VDD93.n143 VDD93.n136 6.3005
R3406 VDD93.n146 VDD93.n133 6.3005
R3407 VDD93.n149 VDD93.n130 6.3005
R3408 VDD93.n152 VDD93.n128 6.3005
R3409 VDD93.n332 VDD93.n159 6.3005
R3410 VDD93.n325 VDD93.n166 6.3005
R3411 VDD93.n320 VDD93.n169 6.3005
R3412 VDD93.n314 VDD93.n174 6.3005
R3413 VDD93.n317 VDD93.n172 6.3005
R3414 VDD93.n324 VDD93.n167 6.3005
R3415 VDD93.n329 VDD93.n163 6.3005
R3416 VDD93.n335 VDD93.n157 6.3005
R3417 VDD93.n341 VDD93.n125 6.3005
R3418 VDD93.n122 VDD93.n121 6.3005
R3419 VDD93.n114 VDD93.n113 6.3005
R3420 VDD93.n342 VDD93.n102 6.3005
R3421 VDD93.n343 VDD93.n101 6.3005
R3422 VDD93.n345 VDD93.n344 6.3005
R3423 VDD93.n425 VDD93.n99 6.3005
R3424 VDD93.n429 VDD93.n96 6.3005
R3425 VDD93 VDD93.n93 6.3005
R3426 VDD93 VDD93.n94 6.3005
R3427 VDD93.n436 VDD93.n435 6.3005
R3428 VDD93.n66 VDD93.n53 6.3005
R3429 VDD93.n69 VDD93.n50 6.3005
R3430 VDD93.n72 VDD93.n47 6.3005
R3431 VDD93.n75 VDD93.n45 6.3005
R3432 VDD93.n476 VDD93.n88 6.3005
R3433 VDD93.n479 VDD93.n85 6.3005
R3434 VDD93.n483 VDD93.n81 6.3005
R3435 VDD93.n487 VDD93.n78 6.3005
R3436 VDD93.n493 VDD93.n41 6.3005
R3437 VDD93.n22 VDD93.n21 6.3005
R3438 VDD93.n25 VDD93.n18 6.3005
R3439 VDD93.n28 VDD93.n15 6.3005
R3440 VDD93.n31 VDD93.n13 6.3005
R3441 VDD93.n495 VDD93.n494 6.3005
R3442 VDD93.n40 VDD93.n39 6.3005
R3443 VDD93.n35 VDD93.n34 6.3005
R3444 VDD93.n503 VDD93.n4 6.3005
R3445 VDD93.n509 VDD93.n0 6.3005
R3446 VDD93.n490 VDD93.n43 6.15559
R3447 VDD93.n485 VDD93.n79 6.1505
R3448 VDD93.n480 VDD93.n83 6.13918
R3449 VDD93.n475 VDD93.n472 6.13239
R3450 VDD93.n439 VDD93.n438 6.01749
R3451 VDD93.n255 VDD93.t301 5.85907
R3452 VDD93.n312 VDD93.t148 5.85907
R3453 VDD93.n337 VDD93.n155 5.85007
R3454 VDD93.n280 VDD93.n204 5.85007
R3455 VDD93.n507 VDD93.n506 5.50832
R3456 VDD93 VDD93.n470 5.38904
R3457 VDD93.n501 VDD93.n2 5.32833
R3458 VDD93.n506 VDD93.n505 5.32746
R3459 VDD93.n22 VDD93.t102 5.213
R3460 VDD93 VDD93.t278 5.1878
R3461 VDD93.n366 VDD93.n365 5.15595
R3462 VDD93 VDD93.t128 5.1508
R3463 VDD93.n458 VDD93.n455 5.13287
R3464 VDD93.n460 VDD93.t344 5.13287
R3465 VDD93.n462 VDD93.n452 5.13287
R3466 VDD93.n90 VDD93.t434 5.13287
R3467 VDD93.n448 VDD93.n91 5.13287
R3468 VDD93.n443 VDD93.t134 5.13287
R3469 VDD93.n442 VDD93.n92 5.13287
R3470 VDD93.n409 VDD93.t105 5.13287
R3471 VDD93.n412 VDD93.t426 5.13287
R3472 VDD93.n415 VDD93.t338 5.13287
R3473 VDD93.n417 VDD93.n396 5.13287
R3474 VDD93.n418 VDD93.t132 5.13287
R3475 VDD93.n420 VDD93.n394 5.13287
R3476 VDD93.n346 VDD93.t438 5.13287
R3477 VDD93.n334 VDD93.n158 5.13287
R3478 VDD93.n327 VDD93.n164 5.13287
R3479 VDD93.n323 VDD93.t123 5.13287
R3480 VDD93.n321 VDD93.n168 5.13287
R3481 VDD93.n318 VDD93.t346 5.13287
R3482 VDD93.n316 VDD93.n173 5.13287
R3483 VDD93.n313 VDD93.t323 5.13287
R3484 VDD93.n277 VDD93.n207 5.13287
R3485 VDD93.n270 VDD93.n213 5.13287
R3486 VDD93.n266 VDD93.t266 5.13287
R3487 VDD93.n264 VDD93.n217 5.13287
R3488 VDD93.n261 VDD93.t386 5.13287
R3489 VDD93.n259 VDD93.n222 5.13287
R3490 VDD93.n256 VDD93.t235 5.13287
R3491 VDD93.n237 VDD93.n231 5.13287
R3492 VDD93.n230 VDD93.n229 5.13287
R3493 VDD93.n246 VDD93.n226 5.13287
R3494 VDD93.n249 VDD93.t388 5.13287
R3495 VDD93.n248 VDD93.n247 5.13287
R3496 VDD93.n254 VDD93.t306 5.13287
R3497 VDD93.n258 VDD93.t96 5.13287
R3498 VDD93.n265 VDD93.t342 5.13287
R3499 VDD93.n269 VDD93.n214 5.13287
R3500 VDD93.n271 VDD93.t231 5.13287
R3501 VDD93.n274 VDD93.n209 5.13287
R3502 VDD93.n276 VDD93.t233 5.13287
R3503 VDD93.n279 VDD93.n205 5.13287
R3504 VDD93.n191 VDD93.t72 5.13287
R3505 VDD93.n194 VDD93.t62 5.13287
R3506 VDD93.n197 VDD93.t169 5.13287
R3507 VDD93.n199 VDD93.n178 5.13287
R3508 VDD93.n200 VDD93.t227 5.13287
R3509 VDD93.n202 VDD93.n176 5.13287
R3510 VDD93.n293 VDD93.n287 5.13287
R3511 VDD93.n286 VDD93.n285 5.13287
R3512 VDD93.n302 VDD93.n282 5.13287
R3513 VDD93.n305 VDD93.t348 5.13287
R3514 VDD93.n304 VDD93.n303 5.13287
R3515 VDD93.n310 VDD93.t272 5.13287
R3516 VDD93.n315 VDD93.t82 5.13287
R3517 VDD93.n322 VDD93.t316 5.13287
R3518 VDD93.n326 VDD93.n165 5.13287
R3519 VDD93.n328 VDD93.t363 5.13287
R3520 VDD93.n331 VDD93.n160 5.13287
R3521 VDD93.n333 VDD93.t17 5.13287
R3522 VDD93.n336 VDD93.n156 5.13287
R3523 VDD93.n142 VDD93.t99 5.13287
R3524 VDD93.n145 VDD93.t314 5.13287
R3525 VDD93.n148 VDD93.t370 5.13287
R3526 VDD93.n150 VDD93.n129 5.13287
R3527 VDD93.n151 VDD93.t251 5.13287
R3528 VDD93.n153 VDD93.n127 5.13287
R3529 VDD93.n126 VDD93.t75 5.13287
R3530 VDD93.n106 VDD93.n105 5.13287
R3531 VDD93.n123 VDD93.t274 5.13287
R3532 VDD93.n107 VDD93.t190 5.13287
R3533 VDD93.n111 VDD93.n110 5.13287
R3534 VDD93.n115 VDD93.t46 5.13287
R3535 VDD93.n119 VDD93.n118 5.13287
R3536 VDD93.n116 VDD93.t310 5.13287
R3537 VDD93.n112 VDD93.n109 5.13287
R3538 VDD93.n426 VDD93.n98 5.13287
R3539 VDD93.n430 VDD93.n95 5.13287
R3540 VDD93.n428 VDD93.t328 5.13287
R3541 VDD93.n68 VDD93.t121 5.13287
R3542 VDD93.n71 VDD93.t57 5.13287
R3543 VDD93.n73 VDD93.n46 5.13287
R3544 VDD93.n74 VDD93.t130 5.13287
R3545 VDD93.n76 VDD93.n44 5.13287
R3546 VDD93.n496 VDD93.t340 5.13287
R3547 VDD93.n9 VDD93.n8 5.13287
R3548 VDD93.n38 VDD93.t48 5.13287
R3549 VDD93.n37 VDD93.n10 5.13287
R3550 VDD93.n36 VDD93.t188 5.13287
R3551 VDD93.n33 VDD93.n11 5.13287
R3552 VDD93.n24 VDD93.t312 5.13287
R3553 VDD93.n27 VDD93.t55 5.13287
R3554 VDD93.n29 VDD93.n14 5.13287
R3555 VDD93.n30 VDD93.t378 5.13287
R3556 VDD93.n32 VDD93.n12 5.13287
R3557 VDD93 VDD93.n469 5.13104
R3558 VDD93 VDD93.t206 5.12757
R3559 VDD93.n502 VDD93.t214 5.12339
R3560 VDD93.n504 VDD93.n3 5.12339
R3561 VDD93.n474 VDD93.t245 5.11708
R3562 VDD93.n478 VDD93.t25 5.11708
R3563 VDD93.n481 VDD93.n82 5.11708
R3564 VDD93.n482 VDD93.t299 5.11708
R3565 VDD93.n484 VDD93.n80 5.11708
R3566 VDD93.n486 VDD93.t418 5.11708
R3567 VDD93.n488 VDD93.n77 5.11708
R3568 VDD93.n42 VDD93.t111 5.11708
R3569 VDD93 VDD93.t330 5.10366
R3570 VDD93 VDD93.t318 5.10321
R3571 VDD93.n378 VDD93.n359 5.09836
R3572 VDD93.n374 VDD93.n361 5.09836
R3573 VDD93.n370 VDD93.n363 5.09836
R3574 VDD93.n381 VDD93.n357 5.09836
R3575 VDD93.n383 VDD93.t295 5.09836
R3576 VDD93.n353 VDD93.n352 5.09836
R3577 VDD93.n388 VDD93.t201 5.09836
R3578 VDD93.n389 VDD93.n351 5.09836
R3579 VDD93.n390 VDD93.t255 5.09836
R3580 VDD93.n350 VDD93.n349 5.09836
R3581 VDD93.n393 VDD93.t253 5.09836
R3582 VDD93.n459 VDD93.t1 5.09407
R3583 VDD93.n463 VDD93.t268 5.09407
R3584 VDD93.n447 VDD93.t436 5.09407
R3585 VDD93.n441 VDD93.t182 5.09407
R3586 VDD93.n339 VDD93.t443 5.09407
R3587 VDD93.n427 VDD93.t69 5.09407
R3588 VDD93.n432 VDD93.t361 5.09407
R3589 VDD93.n431 VDD93.t359 5.09407
R3590 VDD93.n433 VDD93.t472 5.09407
R3591 VDD93.n491 VDD93.t216 5.09407
R3592 VDD93.n1 VDD93.t249 5.09407
R3593 VDD93.n380 VDD93.n379 5.01052
R3594 VDD93.n348 VDD93.n347 4.97242
R3595 VDD93.n421 VDD93.n393 4.93241
R3596 VDD93.n65 VDD93.t89 4.8755
R3597 VDD93.n369 VDD93.n362 4.5905
R3598 VDD93.n373 VDD93.n360 4.5905
R3599 VDD93.n377 VDD93.n358 4.5905
R3600 VDD93.n93 VDD93.t360 4.26489
R3601 VDD93.n94 VDD93.t358 4.26489
R3602 VDD93.n437 VDD93.t31 4.12326
R3603 VDD93.n511 VDD93.t247 4.11379
R3604 VDD93.n140 VDD93.n139 4.08741
R3605 VDD93 VDD93.n232 4.08362
R3606 VDD93.n187 VDD93.n186 4.07437
R3607 VDD93.n407 VDD93.n406 4.07346
R3608 VDD93.n189 VDD93.n188 4.06995
R3609 VDD93.n138 VDD93.n137 4.06354
R3610 VDD93 VDD93.n288 4.0592
R3611 VDD93.n405 VDD93.n404 4.05141
R3612 VDD93.n291 VDD93.n290 4.04913
R3613 VDD93.n368 VDD93.n367 4.00852
R3614 VDD93.n372 VDD93.n371 4.00852
R3615 VDD93.n376 VDD93.n375 4.00852
R3616 VDD93.n234 VDD93.n233 4.0005
R3617 VDD93.n60 VDD93.n59 3.61662
R3618 VDD93.n387 VDD93.n386 3.1505
R3619 VDD93.n387 VDD93.n354 3.1505
R3620 VDD93.n391 VDD93 3.1505
R3621 VDD93 VDD93.n392 3.1505
R3622 VDD93.n190 VDD93.n187 3.06712
R3623 VDD93.n141 VDD93.n138 3.0645
R3624 VDD93.n292 VDD93.n291 3.00562
R3625 VDD93.n408 VDD93.n405 2.95066
R3626 VDD93.n471 VDD93 2.93419
R3627 VDD93.n141 VDD93.n140 2.92128
R3628 VDD93.n236 VDD93.n235 2.91332
R3629 VDD93.n411 VDD93.n402 2.85787
R3630 VDD93.n414 VDD93.n399 2.85787
R3631 VDD93.n330 VDD93.n162 2.85787
R3632 VDD93.n273 VDD93.n211 2.85787
R3633 VDD93.n240 VDD93.n239 2.85787
R3634 VDD93.n245 VDD93.n228 2.85787
R3635 VDD93.n262 VDD93.n220 2.85787
R3636 VDD93.n193 VDD93.n184 2.85787
R3637 VDD93.n196 VDD93.n181 2.85787
R3638 VDD93.n296 VDD93.n295 2.85787
R3639 VDD93.n301 VDD93.n284 2.85787
R3640 VDD93.n319 VDD93.n171 2.85787
R3641 VDD93.n144 VDD93.n135 2.85787
R3642 VDD93.n147 VDD93.n132 2.85787
R3643 VDD93.n124 VDD93.n104 2.85787
R3644 VDD93.n67 VDD93.n52 2.85787
R3645 VDD93.n70 VDD93.n49 2.85787
R3646 VDD93.n497 VDD93.n7 2.85787
R3647 VDD93.n23 VDD93.n20 2.85787
R3648 VDD93.n26 VDD93.n17 2.85787
R3649 VDD93.n190 VDD93.n189 2.85553
R3650 VDD93.n477 VDD93.n87 2.84208
R3651 VDD93.n236 VDD93 2.82101
R3652 VDD93.n292 VDD93.n289 2.8124
R3653 VDD93.n408 VDD93.n407 2.79396
R3654 VDD93.n402 VDD93.t33 2.2755
R3655 VDD93.n402 VDD93.n401 2.2755
R3656 VDD93.n399 VDD93.t308 2.2755
R3657 VDD93.n399 VDD93.n398 2.2755
R3658 VDD93.n162 VDD93.t470 2.2755
R3659 VDD93.n162 VDD93.n161 2.2755
R3660 VDD93.n211 VDD93.t270 2.2755
R3661 VDD93.n211 VDD93.n210 2.2755
R3662 VDD93.n239 VDD93.t276 2.2755
R3663 VDD93.n239 VDD93.n238 2.2755
R3664 VDD93.n228 VDD93.t410 2.2755
R3665 VDD93.n228 VDD93.n227 2.2755
R3666 VDD93.n220 VDD93.t164 2.2755
R3667 VDD93.n220 VDD93.n219 2.2755
R3668 VDD93.n184 VDD93.t150 2.2755
R3669 VDD93.n184 VDD93.n183 2.2755
R3670 VDD93.n181 VDD93.t229 2.2755
R3671 VDD93.n181 VDD93.n180 2.2755
R3672 VDD93.n295 VDD93.t465 2.2755
R3673 VDD93.n295 VDD93.n294 2.2755
R3674 VDD93.n284 VDD93.t393 2.2755
R3675 VDD93.n284 VDD93.n283 2.2755
R3676 VDD93.n171 VDD93.t9 2.2755
R3677 VDD93.n171 VDD93.n170 2.2755
R3678 VDD93.n135 VDD93.t445 2.2755
R3679 VDD93.n135 VDD93.n134 2.2755
R3680 VDD93.n132 VDD93.t365 2.2755
R3681 VDD93.n132 VDD93.n131 2.2755
R3682 VDD93.n104 VDD93.t64 2.2755
R3683 VDD93.n104 VDD93.n103 2.2755
R3684 VDD93.n87 VDD93.t171 2.2755
R3685 VDD93.n87 VDD93.n86 2.2755
R3686 VDD93.n52 VDD93.t119 2.2755
R3687 VDD93.n52 VDD93.n51 2.2755
R3688 VDD93.n49 VDD93.t297 2.2755
R3689 VDD93.n49 VDD93.n48 2.2755
R3690 VDD93.n7 VDD93.t243 2.2755
R3691 VDD93.n7 VDD93.n6 2.2755
R3692 VDD93.n20 VDD93.t372 2.2755
R3693 VDD93.n20 VDD93.n19 2.2755
R3694 VDD93.n17 VDD93.t50 2.2755
R3695 VDD93.n17 VDD93.n16 2.2755
R3696 VDD93.n293 VDD93.n292 2.27547
R3697 VDD93.n237 VDD93.n236 2.27315
R3698 VDD93.n142 VDD93.n141 2.26966
R3699 VDD93.n191 VDD93.n190 2.26502
R3700 VDD93.n409 VDD93.n408 2.26153
R3701 VDD93.n55 VDD93.n54 2.11318
R3702 VDD93 VDD93.n387 1.5755
R3703 VDD93.n57 VDD93.n56 1.54785
R3704 VDD93.n438 VDD93 1.37899
R3705 VDD93 VDD93.n254 1.21661
R3706 VDD93.n281 VDD93.n202 1.18347
R3707 VDD93.n33 VDD93.n32 1.16167
R3708 VDD93.n338 VDD93.n153 1.12775
R3709 VDD93.n311 VDD93.n310 1.12407
R3710 VDD93.n489 VDD93.n76 1.01882
R3711 VDD93.n422 VDD93.n421 0.986314
R3712 VDD93.n59 VDD93.n58 0.840632
R3713 VDD93.n499 VDD93.n5 0.7205
R3714 VDD93.n471 VDD93.n467 0.653723
R3715 VDD93.n422 VDD93.n348 0.559447
R3716 VDD93.n500 VDD93 0.492105
R3717 VDD93.n499 VDD93.n498 0.487926
R3718 VDD93.n472 VDD93.n471 0.411399
R3719 VDD93.n500 VDD93.n499 0.392579
R3720 VDD93.n436 VDD93.n433 0.388218
R3721 VDD93 VDD93.n499 0.386682
R3722 VDD93.n467 VDD93.n466 0.341963
R3723 VDD93.n66 VDD93.n65 0.337997
R3724 VDD93.n65 VDD93.n64 0.328132
R3725 VDD93.n348 VDD93.n346 0.279974
R3726 VDD93.n43 VDD93.n2 0.247933
R3727 VDD93.n466 VDD93.n465 0.247664
R3728 VDD93.n415 VDD93.n414 0.233919
R3729 VDD93.n412 VDD93.n411 0.233919
R3730 VDD93.n240 VDD93.n230 0.233919
R3731 VDD93.n246 VDD93.n245 0.233919
R3732 VDD93.n197 VDD93.n196 0.233919
R3733 VDD93.n194 VDD93.n193 0.233919
R3734 VDD93.n296 VDD93.n286 0.233919
R3735 VDD93.n302 VDD93.n301 0.233919
R3736 VDD93.n148 VDD93.n147 0.233919
R3737 VDD93.n145 VDD93.n144 0.233919
R3738 VDD93.n71 VDD93.n70 0.233919
R3739 VDD93.n68 VDD93.n67 0.233919
R3740 VDD93.n27 VDD93.n26 0.233919
R3741 VDD93.n24 VDD93.n23 0.233919
R3742 VDD93.n472 VDD93.n83 0.224828
R3743 VDD93.n465 VDD93 0.213007
R3744 VDD93.n83 VDD93.n79 0.205754
R3745 VDD93.n79 VDD93.n43 0.193664
R3746 VDD93.n311 VDD93.n281 0.178068
R3747 VDD93.n470 VDD93 0.174585
R3748 VDD93.n506 VDD93.n2 0.16653
R3749 VDD93.n511 VDD93 0.162783
R3750 VDD93.n339 VDD93.n338 0.162742
R3751 VDD93 VDD93.n507 0.155173
R3752 VDD93.n369 VDD93 0.143635
R3753 VDD93.n373 VDD93 0.143635
R3754 VDD93.n377 VDD93 0.143635
R3755 VDD93.n418 VDD93.n417 0.141016
R3756 VDD93.n249 VDD93.n248 0.141016
R3757 VDD93.n200 VDD93.n199 0.141016
R3758 VDD93.n305 VDD93.n304 0.141016
R3759 VDD93.n151 VDD93.n150 0.141016
R3760 VDD93.n74 VDD93.n73 0.141016
R3761 VDD93.n30 VDD93.n29 0.141016
R3762 VDD93.n37 VDD93.n36 0.141016
R3763 VDD93.n38 VDD93.n9 0.141016
R3764 VDD93 VDD93.n42 0.13207
R3765 VDD93.n474 VDD93 0.13207
R3766 VDD93.n428 VDD93 0.126036
R3767 VDD93.n432 VDD93 0.125632
R3768 VDD93 VDD93.n496 0.122435
R3769 VDD93 VDD93.n234 0.121547
R3770 VDD93.n443 VDD93.n89 0.121517
R3771 VDD93.n438 VDD93.n437 0.119239
R3772 VDD93.n460 VDD93 0.11887
R3773 VDD93.n467 VDD93 0.112318
R3774 VDD93.n497 VDD93 0.111984
R3775 VDD93.n437 VDD93 0.110164
R3776 VDD93.n420 VDD93.n419 0.107339
R3777 VDD93.n417 VDD93.n416 0.107339
R3778 VDD93.n250 VDD93.n249 0.107339
R3779 VDD93.n254 VDD93.n253 0.107339
R3780 VDD93.n202 VDD93.n201 0.107339
R3781 VDD93.n199 VDD93.n198 0.107339
R3782 VDD93.n306 VDD93.n305 0.107339
R3783 VDD93.n310 VDD93.n309 0.107339
R3784 VDD93.n153 VDD93.n152 0.107339
R3785 VDD93.n150 VDD93.n149 0.107339
R3786 VDD93.n76 VDD93.n75 0.107339
R3787 VDD93.n73 VDD93.n72 0.107339
R3788 VDD93.n32 VDD93.n31 0.107339
R3789 VDD93.n29 VDD93.n28 0.107339
R3790 VDD93.n35 VDD93.n33 0.107339
R3791 VDD93.n39 VDD93.n37 0.107339
R3792 VDD93.n495 VDD93.n9 0.107339
R3793 VDD93.n55 VDD93 0.106795
R3794 VDD93 VDD93.n240 0.106758
R3795 VDD93.n245 VDD93 0.106758
R3796 VDD93 VDD93.n296 0.106758
R3797 VDD93.n301 VDD93 0.106758
R3798 VDD93.n414 VDD93 0.106177
R3799 VDD93.n411 VDD93 0.106177
R3800 VDD93.n196 VDD93 0.106177
R3801 VDD93.n193 VDD93 0.106177
R3802 VDD93.n147 VDD93 0.106177
R3803 VDD93.n144 VDD93 0.106177
R3804 VDD93.n70 VDD93 0.106177
R3805 VDD93.n67 VDD93 0.106177
R3806 VDD93.n26 VDD93 0.106177
R3807 VDD93.n23 VDD93 0.106177
R3808 VDD93.n464 VDD93.n90 0.105286
R3809 VDD93.n390 VDD93.n350 0.102798
R3810 VDD93.n389 VDD93.n388 0.102778
R3811 VDD93.n383 VDD93.n353 0.0987707
R3812 VDD93.n459 VDD93.n458 0.0984239
R3813 VDD93.n482 VDD93.n481 0.0981682
R3814 VDD93.n463 VDD93.n462 0.0962255
R3815 VDD93.n442 VDD93.n441 0.0962255
R3816 VDD93.n431 VDD93.n430 0.0962255
R3817 VDD93.n489 VDD93.n488 0.0925179
R3818 VDD93.n504 VDD93.n503 0.0925
R3819 VDD93.n448 VDD93.n447 0.0917202
R3820 VDD93.n427 VDD93.n426 0.0917202
R3821 VDD93.n423 VDD93.n422 0.0908448
R3822 VDD93.n505 VDD93.n504 0.0888696
R3823 VDD93.n478 VDD93 0.0852534
R3824 VDD93 VDD93.n390 0.0815938
R3825 VDD93 VDD93.n389 0.081125
R3826 VDD93 VDD93.n439 0.0810263
R3827 VDD93 VDD93.n126 0.0808411
R3828 VDD93.n413 VDD93.n412 0.080629
R3829 VDD93.n410 VDD93.n409 0.080629
R3830 VDD93.n241 VDD93.n237 0.080629
R3831 VDD93.n244 VDD93.n230 0.080629
R3832 VDD93.n195 VDD93.n194 0.080629
R3833 VDD93.n192 VDD93.n191 0.080629
R3834 VDD93.n297 VDD93.n293 0.080629
R3835 VDD93.n300 VDD93.n286 0.080629
R3836 VDD93.n146 VDD93.n145 0.080629
R3837 VDD93.n143 VDD93.n142 0.080629
R3838 VDD93.n69 VDD93.n68 0.080629
R3839 VDD93.n25 VDD93.n24 0.080629
R3840 VDD93.n465 VDD93.n464 0.0796304
R3841 VDD93.n466 VDD93.n89 0.0796304
R3842 VDD93 VDD93.n418 0.0794677
R3843 VDD93 VDD93.n415 0.0794677
R3844 VDD93 VDD93.n200 0.0794677
R3845 VDD93 VDD93.n197 0.0794677
R3846 VDD93 VDD93.n151 0.0794677
R3847 VDD93 VDD93.n148 0.0794677
R3848 VDD93 VDD93.n74 0.0794677
R3849 VDD93 VDD93.n71 0.0794677
R3850 VDD93 VDD93.n30 0.0794677
R3851 VDD93 VDD93.n27 0.0794677
R3852 VDD93.n36 VDD93 0.0794677
R3853 VDD93 VDD93.n38 0.0794677
R3854 VDD93.n496 VDD93 0.0794677
R3855 VDD93 VDD93.n246 0.0788871
R3856 VDD93.n248 VDD93 0.0788871
R3857 VDD93 VDD93.n302 0.0788871
R3858 VDD93.n304 VDD93 0.0788871
R3859 VDD93.n458 VDD93.n457 0.0782465
R3860 VDD93 VDD93.n477 0.0779888
R3861 VDD93.n462 VDD93.n461 0.0764633
R3862 VDD93.n444 VDD93.n442 0.0764633
R3863 VDD93.n430 VDD93.n429 0.0764633
R3864 VDD93.n491 VDD93.n490 0.0759709
R3865 VDD93.n488 VDD93.n487 0.0747601
R3866 VDD93.n484 VDD93.n483 0.0747601
R3867 VDD93.n393 VDD93 0.0742915
R3868 VDD93.n477 VDD93 0.0739529
R3869 VDD93.n388 VDD93 0.0739434
R3870 VDD93 VDD93.n350 0.0738649
R3871 VDD93 VDD93.n353 0.0735189
R3872 VDD93.n63 VDD93 0.0733571
R3873 VDD93 VDD93.n511 0.073
R3874 VDD93.n449 VDD93.n448 0.0728144
R3875 VDD93.n426 VDD93.n425 0.0728144
R3876 VDD93 VDD93.n433 0.0709717
R3877 VDD93.n498 VDD93.n497 0.0669867
R3878 VDD93 VDD93.n502 0.0655
R3879 VDD93.n501 VDD93.n500 0.0635
R3880 VDD93.n486 VDD93.n485 0.0610381
R3881 VDD93 VDD93.n383 0.0594773
R3882 VDD93 VDD93.n381 0.0591364
R3883 VDD93 VDD93.n370 0.0582099
R3884 VDD93 VDD93.n374 0.0582099
R3885 VDD93 VDD93.n378 0.0576483
R3886 VDD93 VDD93.n486 0.0553879
R3887 VDD93 VDD93.n482 0.0553879
R3888 VDD93 VDD93.n478 0.0553879
R3889 VDD93.n502 VDD93.n501 0.055
R3890 VDD93 VDD93.n460 0.0541697
R3891 VDD93 VDD93.n443 0.0541697
R3892 VDD93 VDD93.n428 0.0541697
R3893 VDD93.n423 VDD93 0.0523961
R3894 VDD93.n424 VDD93.n423 0.0518793
R3895 VDD93 VDD93.n90 0.0515917
R3896 VDD93.n42 VDD93.n5 0.0501413
R3897 VDD93 VDD93.n100 0.0493571
R3898 VDD93.n64 VDD93.n63 0.0471071
R3899 VDD93.n475 VDD93.n474 0.0452982
R3900 VDD93 VDD93.n124 0.0435288
R3901 VDD93.n421 VDD93.n420 0.0434677
R3902 VDD93.n481 VDD93.n480 0.0428767
R3903 VDD93 VDD93.n1 0.0410978
R3904 VDD93.n281 VDD93 0.0403112
R3905 VDD93.n507 VDD93.n0 0.0395
R3906 VDD93 VDD93.n311 0.0394651
R3907 VDD93.n338 VDD93 0.0394564
R3908 VDD93 VDD93.n116 0.0392961
R3909 VDD93.n336 VDD93.n335 0.038569
R3910 VDD93.n314 VDD93.n313 0.038569
R3911 VDD93.n279 VDD93.n278 0.0377135
R3912 VDD93.n257 VDD93.n256 0.0377135
R3913 VDD93.n485 VDD93.n484 0.03763
R3914 VDD93.n62 VDD93.n61 0.0358571
R3915 VDD93.n381 VDD93 0.0352326
R3916 VDD93.n126 VDD93.n125 0.0350961
R3917 VDD93.n64 VDD93.n62 0.03425
R3918 VDD93 VDD93.n459 0.0339978
R3919 VDD93 VDD93.n491 0.0339978
R3920 VDD93 VDD93.n463 0.0332632
R3921 VDD93.n441 VDD93 0.0332632
R3922 VDD93 VDD93.n431 0.0332632
R3923 VDD93.n119 VDD93.n102 0.0326553
R3924 VDD93.n480 VDD93.n479 0.0323834
R3925 VDD93.n325 VDD93.n324 0.0323621
R3926 VDD93.n447 VDD93 0.0317552
R3927 VDD93 VDD93.n427 0.0317552
R3928 VDD93.n122 VDD93.n107 0.0313824
R3929 VDD93.n271 VDD93.n270 0.0312416
R3930 VDD93.n265 VDD93.n264 0.0312416
R3931 VDD93.n505 VDD93.n1 0.0293587
R3932 VDD93.n328 VDD93.n327 0.0282241
R3933 VDD93.n322 VDD93.n321 0.0282241
R3934 VDD93.n268 VDD93.n267 0.0280056
R3935 VDD93.n330 VDD93.n329 0.0273966
R3936 VDD93.n320 VDD93.n319 0.0273966
R3937 VDD93 VDD93.n331 0.0271897
R3938 VDD93.n318 VDD93 0.0269828
R3939 VDD93.n276 VDD93.n275 0.0267921
R3940 VDD93.n260 VDD93.n259 0.0267921
R3941 VDD93 VDD93.n277 0.0263876
R3942 VDD93.n258 VDD93 0.0261854
R3943 VDD93.n333 VDD93.n332 0.0236724
R3944 VDD93.n317 VDD93.n316 0.0236724
R3945 VDD93 VDD93.n334 0.0232586
R3946 VDD93.n273 VDD93.n272 0.0231517
R3947 VDD93.n263 VDD93.n262 0.0231517
R3948 VDD93.n315 VDD93 0.0230517
R3949 VDD93 VDD93.n274 0.0229494
R3950 VDD93.n106 VDD93 0.0228998
R3951 VDD93.n327 VDD93.n326 0.0228448
R3952 VDD93.n323 VDD93.n322 0.0228448
R3953 VDD93.n261 VDD93 0.0227472
R3954 VDD93.n424 VDD93 0.0222241
R3955 VDD93.n111 VDD93.n100 0.0214709
R3956 VDD93 VDD93.n339 0.0207439
R3957 VDD93.n113 VDD93.n112 0.0205971
R3958 VDD93.n270 VDD93.n269 0.0187022
R3959 VDD93.n266 VDD93.n265 0.0187022
R3960 VDD93.n123 VDD93 0.0186765
R3961 VDD93.n291 VDD93 0.0181958
R3962 VDD93.n464 VDD93 0.0174737
R3963 VDD93 VDD93.n328 0.016431
R3964 VDD93.n321 VDD93 0.0162241
R3965 VDD93.n124 VDD93.n123 0.0162059
R3966 VDD93.n187 VDD93 0.0157113
R3967 VDD93.n235 VDD93 0.0152541
R3968 VDD93.n274 VDD93.n273 0.0150618
R3969 VDD93.n262 VDD93.n261 0.0150618
R3970 VDD93.n407 VDD93 0.0133571
R3971 VDD93.n405 VDD93 0.0132059
R3972 VDD93.n112 VDD93.n111 0.0125583
R3973 VDD93.n116 VDD93.n115 0.0125583
R3974 VDD93.n370 VDD93.n369 0.0125512
R3975 VDD93.n374 VDD93.n373 0.0125512
R3976 VDD93.n378 VDD93.n377 0.0125094
R3977 VDD93 VDD93.n271 0.0124326
R3978 VDD93.n264 VDD93 0.0122303
R3979 VDD93.n115 VDD93 0.0122087
R3980 VDD93.n331 VDD93.n330 0.0116724
R3981 VDD93.n319 VDD93.n318 0.0116724
R3982 VDD93.n476 VDD93.n475 0.0113969
R3983 VDD93 VDD93.n101 0.0111602
R3984 VDD93.n138 VDD93 0.0110882
R3985 VDD93.n346 VDD93.n345 0.0105519
R3986 VDD93.n189 VDD93 0.00981034
R3987 VDD93 VDD93.n266 0.00980337
R3988 VDD93.n269 VDD93 0.00960112
R3989 VDD93 VDD93.n432 0.00839474
R3990 VDD93.n490 VDD93.n489 0.00816816
R3991 VDD93.n41 VDD93.n5 0.00655381
R3992 VDD93.n337 VDD93.n336 0.0065
R3993 VDD93 VDD93.n323 0.0062931
R3994 VDD93.n313 VDD93.n312 0.0062931
R3995 VDD93.n326 VDD93 0.00608621
R3996 VDD93.n334 VDD93.n333 0.00587931
R3997 VDD93.n316 VDD93.n315 0.00587931
R3998 VDD93.n289 VDD93 0.00579412
R3999 VDD93 VDD93.n436 0.00579412
R4000 VDD93 VDD93.n89 0.00501883
R4001 VDD93.n498 VDD93 0.00493946
R4002 VDD93.n63 VDD93 0.00478571
R4003 VDD93.n503 VDD93 0.0045
R4004 VDD93.n235 VDD93.n234 0.00419863
R4005 VDD93.n439 VDD93 0.00400649
R4006 VDD93 VDD93.n0 0.004
R4007 VDD93.n457 VDD93 0.00388028
R4008 VDD93.n461 VDD93 0.00380275
R4009 VDD93.n444 VDD93 0.00380275
R4010 VDD93.n429 VDD93 0.00380275
R4011 VDD93.n61 VDD93.n60 0.00371429
R4012 VDD93.n449 VDD93 0.0036441
R4013 VDD93.n140 VDD93 0.00307143
R4014 VDD93.n280 VDD93.n279 0.00272472
R4015 VDD93.n256 VDD93.n255 0.00252247
R4016 VDD93.n117 VDD93 0.00242233
R4017 VDD93.n250 VDD93 0.00224194
R4018 VDD93.n253 VDD93 0.00224194
R4019 VDD93.n306 VDD93 0.00224194
R4020 VDD93.n309 VDD93 0.00224194
R4021 VDD93.n277 VDD93.n276 0.00211798
R4022 VDD93.n259 VDD93.n258 0.00211798
R4023 VDD93.n60 VDD93.n57 0.00210714
R4024 VDD93.n107 VDD93.n106 0.00208824
R4025 VDD93 VDD93.n122 0.00191176
R4026 VDD93.n113 VDD93 0.00189806
R4027 VDD93 VDD93.n119 0.0017233
R4028 VDD93.n366 VDD93.n364 0.00167963
R4029 VDD93.n423 VDD93.n100 0.00166883
R4030 VDD93.n345 VDD93 0.00166883
R4031 VDD93.n419 VDD93 0.00166129
R4032 VDD93.n416 VDD93 0.00166129
R4033 VDD93 VDD93.n413 0.00166129
R4034 VDD93 VDD93.n410 0.00166129
R4035 VDD93.n201 VDD93 0.00166129
R4036 VDD93.n198 VDD93 0.00166129
R4037 VDD93 VDD93.n195 0.00166129
R4038 VDD93 VDD93.n192 0.00166129
R4039 VDD93.n152 VDD93 0.00166129
R4040 VDD93.n149 VDD93 0.00166129
R4041 VDD93 VDD93.n146 0.00166129
R4042 VDD93 VDD93.n143 0.00166129
R4043 VDD93.n75 VDD93 0.00166129
R4044 VDD93.n72 VDD93 0.00166129
R4045 VDD93 VDD93.n69 0.00166129
R4046 VDD93 VDD93.n66 0.00166129
R4047 VDD93.n31 VDD93 0.00166129
R4048 VDD93.n28 VDD93 0.00166129
R4049 VDD93 VDD93.n25 0.00166129
R4050 VDD93 VDD93.n22 0.00166129
R4051 VDD93 VDD93.n35 0.00166129
R4052 VDD93.n39 VDD93 0.00166129
R4053 VDD93 VDD93.n495 0.00166129
R4054 VDD93.n289 VDD93 0.00155882
R4055 VDD93 VDD93.n358 0.00152662
R4056 VDD93.n41 VDD93 0.00130718
R4057 VDD93.n487 VDD93 0.00130718
R4058 VDD93.n483 VDD93 0.00130718
R4059 VDD93.n479 VDD93 0.00130718
R4060 VDD93 VDD93.n476 0.00130718
R4061 VDD93 VDD93.n364 0.00118702
R4062 VDD93 VDD93.n362 0.00118702
R4063 VDD93 VDD93.n362 0.00118702
R4064 VDD93 VDD93.n360 0.00118702
R4065 VDD93 VDD93.n360 0.00118702
R4066 VDD93 VDD93.n358 0.00118441
R4067 VDD93 VDD93.n325 0.00112069
R4068 VDD93 VDD93.n320 0.00112069
R4069 VDD93 VDD93.n314 0.00112069
R4070 VDD93 VDD93.n268 0.00110674
R4071 VDD93 VDD93.n263 0.00110674
R4072 VDD93 VDD93.n257 0.00110674
R4073 VDD93.n241 VDD93 0.00108064
R4074 VDD93 VDD93.n244 0.00108064
R4075 VDD93.n297 VDD93 0.00108064
R4076 VDD93 VDD93.n300 0.00108064
R4077 VDD93 VDD93.n366 0.00100731
R4078 VDD93.n125 VDD93 0.00100139
R4079 VDD93 VDD93.n337 0.000913793
R4080 VDD93.n335 VDD93 0.000913793
R4081 VDD93.n329 VDD93 0.000913793
R4082 VDD93.n324 VDD93 0.000913793
R4083 VDD93 VDD93.n317 0.000913793
R4084 VDD93.n312 VDD93 0.000913793
R4085 VDD93 VDD93.n280 0.000904494
R4086 VDD93.n278 VDD93 0.000904494
R4087 VDD93.n272 VDD93 0.000904494
R4088 VDD93.n267 VDD93 0.000904494
R4089 VDD93 VDD93.n260 0.000904494
R4090 VDD93.n255 VDD93 0.000904494
R4091 VDD93.n425 VDD93.n424 0.000893013
R4092 VDD93 VDD93.n101 0.000849515
R4093 VDD93 VDD93.n117 0.000849515
R4094 VDD93 VDD93.n102 0.000849515
R4095 VDD93.n332 VDD93 0.000706897
R4096 VDD93.n275 VDD93 0.000702247
R4097 VSS.n3467 VSS.n18 7.8912e+06
R4098 VSS.t420 VSS.n987 4.82147e+06
R4099 VSS.n3467 VSS.n3466 4.7548e+06
R4100 VSS.n2979 VSS.n18 4.745e+06
R4101 VSS.n2617 VSS.n2616 303512
R4102 VSS.n1884 VSS.n1883 291723
R4103 VSS.n1206 VSS.n1205 132150
R4104 VSS.n525 VSS.n510 106315
R4105 VSS.n2846 VSS.t1650 94673.9
R4106 VSS.n3335 VSS.n3334 89067.6
R4107 VSS.n1924 VSS.n1923 87750
R4108 VSS.n1901 VSS.n1900 71260
R4109 VSS.n514 VSS.n513 53002.1
R4110 VSS.n385 VSS.t739 50344.7
R4111 VSS.n3336 VSS.n3335 44326.9
R4112 VSS.t31 VSS.n1924 40776.9
R4113 VSS.n1900 VSS.n1899 39263.5
R4114 VSS.t1337 VSS.n244 38626.7
R4115 VSS.n1218 VSS.n1206 33732.1
R4116 VSS.n3389 VSS.n3384 32328.9
R4117 VSS.n672 VSS.t1956 25318.3
R4118 VSS.t2378 VSS.n1178 23296.6
R4119 VSS.n517 VSS.n516 21267.7
R4120 VSS.t1983 VSS.n2937 21110.5
R4121 VSS.n3271 VSS.n3270 20815.8
R4122 VSS.n3289 VSS.n117 20141.5
R4123 VSS.n1883 VSS.t517 19851.6
R4124 VSS.n1906 VSS.n1223 19564.1
R4125 VSS.n301 VSS.n300 19500
R4126 VSS.t499 VSS.n1904 18875.9
R4127 VSS.t1241 VSS.n3387 18875.9
R4128 VSS.n2080 VSS.n2063 18801.2
R4129 VSS.n1961 VSS.n1960 18801.2
R4130 VSS.n2445 VSS.n2444 18801.2
R4131 VSS.n438 VSS.n416 18801.2
R4132 VSS.n472 VSS.n386 18801.2
R4133 VSS.n1958 VSS.n1956 18801.2
R4134 VSS.n2061 VSS.n2059 18801.2
R4135 VSS.n1057 VSS.t2153 16947.9
R4136 VSS.t2313 VSS.n1463 16930.7
R4137 VSS.n306 VSS.n301 16250
R4138 VSS.t2498 VSS.t1919 16169.8
R4139 VSS.n2595 VSS.t2222 16128.7
R4140 VSS.n685 VSS.t103 15778.8
R4141 VSS.n3167 VSS.n277 15396.1
R4142 VSS.t441 VSS.n2510 15180.4
R4143 VSS.n2939 VSS.n2938 14010
R4144 VSS.n3339 VSS.n3338 13936
R4145 VSS.n457 VSS.n411 13936
R4146 VSS.n986 VSS.n255 13818.6
R4147 VSS.n2594 VSS.n2593 13763.2
R4148 VSS.n2814 VSS.n2813 13000
R4149 VSS.n3421 VSS.t65 12600.2
R4150 VSS.n54 VSS.n53 12212.1
R4151 VSS.n3167 VSS.n3166 11877.7
R4152 VSS.t859 VSS.n1092 11866
R4153 VSS.t1176 VSS.n1292 11866
R4154 VSS.t535 VSS.n1380 11866
R4155 VSS.t1164 VSS.n1004 11866
R4156 VSS.t1071 VSS.n2139 11866
R4157 VSS.t1728 VSS.n3081 11766.3
R4158 VSS.n2222 VSS.n2221 11621.2
R4159 VSS.n2796 VSS.n2795 11423.9
R4160 VSS.n2848 VSS.n2845 11193.5
R4161 VSS.n74 VSS.n68 11109.4
R4162 VSS.n1143 VSS.n1142 11104.2
R4163 VSS.n519 VSS.n517 11072
R4164 VSS.n1222 VSS.n1126 10903.3
R4165 VSS.n1664 VSS.n1663 10712.2
R4166 VSS.n505 VSS.t377 10467.5
R4167 VSS.n1723 VSS.t717 10467.5
R4168 VSS.n207 VSS.n206 9976.39
R4169 VSS.n2847 VSS.n2846 9810.56
R4170 VSS.n299 VSS.n298 9750
R4171 VSS.n1407 VSS.n1387 9589.42
R4172 VSS.n2167 VSS.n2146 9589.42
R4173 VSS.n1661 VSS.n1620 9589.42
R4174 VSS.n2293 VSS.n1090 9584.01
R4175 VSS.n1309 VSS.n1248 9584.01
R4176 VSS.n3211 VSS.n3210 9580.21
R4177 VSS.n540 VSS.n507 9415.54
R4178 VSS.n1754 VSS.t1904 9200.13
R4179 VSS.n2491 VSS.n2490 8900.19
R4180 VSS.n25 VSS.n24 8870.17
R4181 VSS.n2652 VSS.n2651 8793.57
R4182 VSS.n3466 VSS.n19 8734.15
R4183 VSS.n1057 VSS.t2201 8709.27
R4184 VSS.n3057 VSS.n3014 8615.97
R4185 VSS.n281 VSS.n280 8591.3
R4186 VSS.n1326 VSS.n1325 8434.2
R4187 VSS.n914 VSS.n913 8432.89
R4188 VSS.n1057 VSS.n1030 8422.78
R4189 VSS.n386 VSS.n385 7847.56
R4190 VSS.t1860 VSS.n525 7666.92
R4191 VSS.n2552 VSS.n2542 7369.71
R4192 VSS.n2653 VSS.n2652 7059.24
R4193 VSS.n1725 VSS.t553 7006.49
R4194 VSS.n506 VSS.t1978 7006.49
R4195 VSS.n2969 VSS.n2968 6954.93
R4196 VSS.n1221 VSS.n1220 6949.6
R4197 VSS.n2699 VSS.t1807 6878.25
R4198 VSS.n204 VSS.n203 6643.65
R4199 VSS.n205 VSS.n204 6643.65
R4200 VSS.n524 VSS.n523 6266.68
R4201 VSS.n1203 VSS.n1202 6216.55
R4202 VSS.n3316 VSS.n3299 6129.95
R4203 VSS.n1811 VSS.n912 5850
R4204 VSS.n1219 VSS.n1218 5848.08
R4205 VSS.n159 VSS.n158 5785.02
R4206 VSS.n411 VSS.t1381 5604.27
R4207 VSS.n1773 VSS.n1772 5552.94
R4208 VSS.n3466 VSS.n3465 5328.79
R4209 VSS.n2979 VSS.n2978 5250.54
R4210 VSS.n1541 VSS.n1241 5147.52
R4211 VSS.n184 VSS.n125 5117.4
R4212 VSS.n185 VSS.n124 5117.4
R4213 VSS.n1047 VSS.t1480 5069.75
R4214 VSS.n3338 VSS.n3337 5050.96
R4215 VSS.n2588 VSS.t1372 5021.3
R4216 VSS.n3166 VSS.n3164 4981.69
R4217 VSS.n1214 VSS.n1213 4977.02
R4218 VSS.n520 VSS.n515 4933.75
R4219 VSS.n987 VSS.n986 4911.11
R4220 VSS.n183 VSS.n182 4903.12
R4221 VSS.n1203 VSS.n1199 4795.4
R4222 VSS.n977 VSS.n248 4534.77
R4223 VSS.n1177 VSS.n1176 4512.4
R4224 VSS.n3442 VSS.n3441 4433.19
R4225 VSS.n2600 VSS.n2599 4416.33
R4226 VSS.n634 VSS.n603 4416.33
R4227 VSS.n3269 VSS.n3225 4284.75
R4228 VSS.n3135 VSS.n3134 4274.47
R4229 VSS.n3210 VSS.n3209 4247.05
R4230 VSS.n1142 VSS.n1126 4152.78
R4231 VSS.n24 VSS.n23 4152.58
R4232 VSS.n2590 VSS.t750 4127.74
R4233 VSS.n1540 VSS.t2242 4107.43
R4234 VSS.n3224 VSS.n3223 4041.16
R4235 VSS.n240 VSS.n239 4026.42
R4236 VSS.n3391 VSS.n3390 3956.92
R4237 VSS.n2101 VSS.n2100 3893.61
R4238 VSS.n2145 VSS.n2124 3893.61
R4239 VSS.n2340 VSS.n1084 3893.61
R4240 VSS.n2386 VSS.n1071 3893.61
R4241 VSS.n2341 VSS.n1083 3893.61
R4242 VSS.n1386 VSS.n1365 3893.61
R4243 VSS.n1308 VSS.n1242 3893.61
R4244 VSS.n3351 VSS.n3350 3893.61
R4245 VSS.n494 VSS.n493 3893.61
R4246 VSS.n1444 VSS.n1442 3893.61
R4247 VSS.n2236 VSS.n2235 3893.61
R4248 VSS.n2292 VSS.n1091 3893.61
R4249 VSS.n2038 VSS.n2037 3893.61
R4250 VSS.n947 VSS.n946 3893.61
R4251 VSS.n441 VSS.n440 3893.61
R4252 VSS.n1199 VSS.n1198 3871.27
R4253 VSS.n55 VSS.n54 3870.07
R4254 VSS.n220 VSS.n219 3823.53
R4255 VSS.n153 VSS.n152 3823.53
R4256 VSS.n205 VSS.n202 3823.53
R4257 VSS.n201 VSS.n200 3823.53
R4258 VSS.n199 VSS.n198 3823.53
R4259 VSS.n197 VSS.n196 3823.53
R4260 VSS.n195 VSS.n194 3823.53
R4261 VSS.n207 VSS.n205 3823.53
R4262 VSS.n208 VSS.n201 3823.53
R4263 VSS.n209 VSS.n199 3823.53
R4264 VSS.n210 VSS.n197 3823.53
R4265 VSS.n211 VSS.n195 3823.53
R4266 VSS.n212 VSS.n193 3823.53
R4267 VSS.n213 VSS.n192 3823.53
R4268 VSS.n214 VSS.n191 3823.53
R4269 VSS.n215 VSS.n190 3823.53
R4270 VSS.n216 VSS.n189 3823.53
R4271 VSS.n217 VSS.n188 3823.53
R4272 VSS.n218 VSS.n187 3823.53
R4273 VSS.n178 VSS.n142 3823.53
R4274 VSS.n177 VSS.n143 3823.53
R4275 VSS.n176 VSS.n144 3823.53
R4276 VSS.n175 VSS.n145 3823.53
R4277 VSS.n174 VSS.n146 3823.53
R4278 VSS.n173 VSS.n147 3823.53
R4279 VSS.n172 VSS.n148 3823.53
R4280 VSS.n171 VSS.n149 3823.53
R4281 VSS.n165 VSS.n150 3823.53
R4282 VSS.n164 VSS.n151 3823.53
R4283 VSS.n163 VSS.n153 3823.53
R4284 VSS.n162 VSS.n154 3823.53
R4285 VSS.n161 VSS.n155 3823.53
R4286 VSS.n160 VSS.n156 3823.53
R4287 VSS.n159 VSS.n157 3823.53
R4288 VSS.n181 VSS.n180 3823.53
R4289 VSS.n180 VSS.n179 3823.53
R4290 VSS.n3337 VSS.n3317 3791.26
R4291 VSS.n3168 VSS.n3167 3790.3
R4292 VSS.n3211 VSS.t123 3750
R4293 VSS.n2223 VSS.n2222 3613.6
R4294 VSS.n1981 VSS.t862 3606.54
R4295 VSS.t458 VSS.n1275 3606.54
R4296 VSS.n2426 VSS.t236 3606.54
R4297 VSS.n1409 VSS.t2132 3606.54
R4298 VSS.n2169 VSS.t607 3606.54
R4299 VSS.n1603 VSS.t1770 3606.54
R4300 VSS.n3472 VSS.n3471 3567.93
R4301 VSS.n3337 VSS.n3336 3531.55
R4302 VSS.n1744 VSS.n1553 3525.32
R4303 VSS.n330 VSS.n329 3525.32
R4304 VSS.n2623 VSS.n2622 3472.05
R4305 VSS.n512 VSS.n511 3468.77
R4306 VSS.n1176 VSS.n1175 3357.44
R4307 VSS.n1883 VSS.n1240 3355.98
R4308 VSS.n2589 VSS.n914 3353.53
R4309 VSS.n2980 VSS.n2976 3324.29
R4310 VSS.t75 VSS.n404 3289.63
R4311 VSS.t2226 VSS.n650 3289.63
R4312 VSS.n2702 VSS.n2701 3285.76
R4313 VSS.n1047 VSS.t2451 3278.56
R4314 VSS.t1697 VSS.n2555 3265.82
R4315 VSS.n2555 VSS.t1473 3219.67
R4316 VSS.n2932 VSS.n2931 3214.19
R4317 VSS.n3014 VSS.n3013 3205.8
R4318 VSS.t1701 VSS.n3135 3181.7
R4319 VSS.n1980 VSS.t430 3112.87
R4320 VSS.t460 VSS.n1276 3112.87
R4321 VSS.t370 VSS.n1415 3112.87
R4322 VSS.t1499 VSS.n2175 3112.87
R4323 VSS.n1602 VSS.t1772 3112.87
R4324 VSS.n1906 VSS.n1222 3095.47
R4325 VSS.n1958 VSS.n1957 3086.35
R4326 VSS.n2061 VSS.n2060 3086.35
R4327 VSS.n1960 VSS.n1959 3083.79
R4328 VSS.n2063 VSS.n2062 3083.79
R4329 VSS.n3166 VSS.n3165 3077.65
R4330 VSS.n3133 VSS.n281 3077.65
R4331 VSS.t394 VSS.t1597 3055.32
R4332 VSS.t866 VSS.t864 3055.32
R4333 VSS.t352 VSS.t384 3055.32
R4334 VSS.n185 VSS.n184 3042.38
R4335 VSS.n1883 VSS.n1241 3017.86
R4336 VSS.n1572 VSS.n1565 3004.05
R4337 VSS.n1492 VSS.t1188 2999.9
R4338 VSS.n2402 VSS.n2401 2983.23
R4339 VSS.n3405 VSS.n68 2983.21
R4340 VSS.n2615 VSS.t1844 2945.13
R4341 VSS.n3472 VSS.t973 2945.13
R4342 VSS.t2335 VSS.n674 2933.7
R4343 VSS.n521 VSS.t1581 2925
R4344 VSS.n141 VSS.t211 2818.91
R4345 VSS.t2386 VSS.n3405 2810.52
R4346 VSS.t1365 VSS.t802 2781.65
R4347 VSS.t389 VSS.t1796 2781.65
R4348 VSS.t771 VSS.t769 2781.65
R4349 VSS.t199 VSS.t2229 2781.65
R4350 VSS.n2591 VSS.n912 2727.5
R4351 VSS.n1216 VSS.n1215 2702.93
R4352 VSS.n13 VSS.n12 2682.86
R4353 VSS.t742 VSS.n3339 2673.11
R4354 VSS.n457 VSS.t2370 2673.11
R4355 VSS.n1483 VSS.n1482 2491.86
R4356 VSS.n2626 VSS.n2625 2416.67
R4357 VSS.n3275 VSS.n185 2315.72
R4358 VSS.t1566 VSS.t1230 2311.62
R4359 VSS.t202 VSS.t650 2311.62
R4360 VSS.t2418 VSS.t253 2311.62
R4361 VSS.t1661 VSS.t1561 2307.56
R4362 VSS.t1058 VSS.t1055 2307.56
R4363 VSS.t1048 VSS.t1049 2307.56
R4364 VSS.t2267 VSS.t1492 2307.56
R4365 VSS.t1900 VSS.t1901 2307.56
R4366 VSS.t1952 VSS.t1953 2307.56
R4367 VSS.t101 VSS.t2014 2307.56
R4368 VSS.t1040 VSS.t1037 2307.56
R4369 VSS.t97 VSS.t2193 2307.56
R4370 VSS.t228 VSS.t231 2307.56
R4371 VSS.t1177 VSS.t850 2307.56
R4372 VSS.t848 VSS.t2463 2307.56
R4373 VSS.t1284 VSS.t1867 2307.56
R4374 VSS.t432 VSS.t92 2307.56
R4375 VSS.t946 VSS.t168 2307.56
R4376 VSS.t302 VSS.t1670 2307.56
R4377 VSS.t1531 VSS.t483 2307.56
R4378 VSS.t49 VSS.t818 2307.56
R4379 VSS.t2503 VSS.t754 2307.56
R4380 VSS.t1788 VSS.t743 2307.56
R4381 VSS.t1435 VSS.t1438 2307.56
R4382 VSS.t762 VSS.t57 2307.56
R4383 VSS.t325 VSS.t421 2307.56
R4384 VSS.t1551 VSS.t951 2307.56
R4385 VSS.t337 VSS.t336 2307.56
R4386 VSS.t64 VSS.t1277 2307.56
R4387 VSS.t1686 VSS.t1535 2307.56
R4388 VSS.t1646 VSS.t661 2307.56
R4389 VSS.t1968 VSS.t1739 2307.56
R4390 VSS.t416 VSS.t22 2307.56
R4391 VSS.t387 VSS.t2254 2307.56
R4392 VSS.t948 VSS.t794 2307.56
R4393 VSS.t975 VSS.t1020 2307.56
R4394 VSS.t204 VSS.t93 2307.56
R4395 VSS.t299 VSS.t300 2307.56
R4396 VSS.t197 VSS.t193 2307.56
R4397 VSS.t239 VSS.t240 2307.56
R4398 VSS.t216 VSS.t2260 2307.56
R4399 VSS.t110 VSS.t88 2307.56
R4400 VSS.t1268 VSS.t135 2307.56
R4401 VSS.t2175 VSS.t1338 2307.56
R4402 VSS.t1992 VSS.t1022 2307.56
R4403 VSS.t472 VSS.t474 2307.56
R4404 VSS.t2541 VSS.t1159 2307.56
R4405 VSS.t10 VSS.t1828 2307.56
R4406 VSS.t1611 VSS.t1613 2307.56
R4407 VSS.t447 VSS.t593 2307.56
R4408 VSS.t1331 VSS.t1330 2307.56
R4409 VSS.t1878 VSS.t1298 2307.56
R4410 VSS.t639 VSS.t2202 2307.56
R4411 VSS.t2546 VSS.t436 2307.56
R4412 VSS.t1400 VSS.t1051 2307.56
R4413 VSS.t174 VSS.t178 2307.56
R4414 VSS.t2452 VSS.t354 2307.56
R4415 VSS.t1453 VSS.t1527 2307.56
R4416 VSS.t1705 VSS.t295 2307.56
R4417 VSS.t1711 VSS.t1700 2307.56
R4418 VSS.t678 VSS.t711 2307.56
R4419 VSS.t551 VSS.t709 2307.56
R4420 VSS.t1663 VSS.t539 2307.56
R4421 VSS.t1586 VSS.t1368 2307.56
R4422 VSS.t1380 VSS.t2544 2307.56
R4423 VSS.t2170 VSS.t1859 2307.56
R4424 VSS.t2104 VSS.t2100 2307.56
R4425 VSS.t40 VSS.t457 2307.56
R4426 VSS.t1926 VSS.t1921 2307.56
R4427 VSS.t20 VSS.t1370 2307.56
R4428 VSS.t602 VSS.t54 2307.56
R4429 VSS.t1282 VSS.t2139 2307.56
R4430 VSS.t2321 VSS.t2348 2307.56
R4431 VSS.t2366 VSS.t1166 2307.56
R4432 VSS.t1855 VSS.t1857 2307.56
R4433 VSS.t130 VSS.t970 2307.56
R4434 VSS.t2154 VSS.t1698 2307.56
R4435 VSS.t2141 VSS.t2143 2307.56
R4436 VSS.t1695 VSS.t2332 2307.56
R4437 VSS.t466 VSS.t1781 2307.56
R4438 VSS.t1723 VSS.t829 2307.56
R4439 VSS.t2086 VSS.t2361 2307.56
R4440 VSS.t2090 VSS.t1765 2307.56
R4441 VSS.t1673 VSS.t1675 2307.56
R4442 VSS.t1709 VSS.t2191 2307.56
R4443 VSS.t2486 VSS.t2307 2307.56
R4444 VSS.t2309 VSS.t1786 2307.56
R4445 VSS.t1808 VSS.t1988 2307.56
R4446 VSS.t1294 VSS.t2320 2307.56
R4447 VSS.t1392 VSS.t1394 2307.56
R4448 VSS.t643 VSS.t645 2307.56
R4449 VSS.t799 VSS.t1353 2307.56
R4450 VSS.t156 VSS.t841 2307.56
R4451 VSS.t876 VSS.t476 2307.56
R4452 VSS.t2453 VSS.t1174 2307.56
R4453 VSS.t1520 VSS.t1799 2307.56
R4454 VSS.t2247 VSS.t1873 2307.56
R4455 VSS.t37 VSS.t983 2307.56
R4456 VSS.t599 VSS.t1264 2307.56
R4457 VSS.t1881 VSS.t2005 2307.56
R4458 VSS.t1916 VSS.t1838 2307.56
R4459 VSS.t929 VSS.t2185 2307.56
R4460 VSS.t1965 VSS.t1964 2307.56
R4461 VSS.t2277 VSS.t2397 2307.56
R4462 VSS.t2326 VSS.t546 2307.56
R4463 VSS.t118 VSS.t1720 2307.56
R4464 VSS.t943 VSS.t2127 2307.56
R4465 VSS.t1258 VSS.t69 2307.56
R4466 VSS.t536 VSS.t72 2307.56
R4467 VSS.t19 VSS.t1850 2307.56
R4468 VSS.t427 VSS.t1905 2307.56
R4469 VSS.t909 VSS.t1608 2307.56
R4470 VSS.t1835 VSS.t1716 2307.56
R4471 VSS.t858 VSS.t1548 2307.56
R4472 VSS.t60 VSS.t2109 2307.56
R4473 VSS.t1839 VSS.t179 2307.56
R4474 VSS.t2084 VSS.t367 2307.56
R4475 VSS.t686 VSS.t1102 2307.56
R4476 VSS.t86 VSS.t1774 2307.56
R4477 VSS.t1130 VSS.t844 2307.56
R4478 VSS.t860 VSS.t2117 2307.56
R4479 VSS.t813 VSS.t814 2307.56
R4480 VSS.t1742 VSS.t2121 2307.56
R4481 VSS.t1861 VSS.t817 2307.56
R4482 VSS.t1426 VSS.t635 2307.56
R4483 VSS.t1429 VSS.t1960 2307.56
R4484 VSS.t1308 VSS.t1449 2307.56
R4485 VSS.t1591 VSS.t1387 2307.56
R4486 VSS.t613 VSS.t1594 2307.56
R4487 VSS.t1221 VSS.t1099 2307.56
R4488 VSS.t568 VSS.t774 2307.56
R4489 VSS.t1545 VSS.t1538 2307.56
R4490 VSS.t1138 VSS.t185 2307.56
R4491 VSS.t2207 VSS.t777 2307.56
R4492 VSS.t1072 VSS.t780 2307.56
R4493 VSS.t2328 VSS.t321 2307.56
R4494 VSS.t331 VSS.t332 2307.56
R4495 VSS.t833 VSS.t831 2307.56
R4496 VSS.t666 VSS.t1575 2307.56
R4497 VSS.t413 VSS.t1891 2307.56
R4498 VSS.t1007 VSS.t869 2307.56
R4499 VSS.t619 VSS.t396 2307.56
R4500 VSS.t1997 VSS.t1996 2307.56
R4501 VSS.t641 VSS.t895 2307.56
R4502 VSS.t544 VSS.t1351 2307.56
R4503 VSS.t2162 VSS.t1827 2307.56
R4504 VSS.t1316 VSS.t148 2307.56
R4505 VSS.t1547 VSS.t481 2307.56
R4506 VSS.t478 VSS.t837 2307.56
R4507 VSS.t963 VSS.t967 2307.56
R4508 VSS.t737 VSS.t572 2307.56
R4509 VSS.t363 VSS.t362 2307.56
R4510 VSS.t2233 VSS.t504 2307.56
R4511 VSS.t992 VSS.t1485 2307.56
R4512 VSS.t1511 VSS.t1489 2307.56
R4513 VSS.t351 VSS.t1913 2307.56
R4514 VSS.t704 VSS.t633 2307.56
R4515 VSS.t1569 VSS.t747 2307.56
R4516 VSS.t702 VSS.t285 2307.56
R4517 VSS.t2094 VSS.t2093 2307.56
R4518 VSS.t1045 VSS.t188 2307.56
R4519 VSS.t50 VSS.t560 2307.56
R4520 VSS.t2371 VSS.t2476 2307.56
R4521 VSS.t2347 VSS.t2294 2307.56
R4522 VSS.t1270 VSS.t1930 2307.56
R4523 VSS.t1640 VSS.t1642 2307.56
R4524 VSS.t854 VSS.t2468 2307.56
R4525 VSS.t2195 VSS.t2304 2307.56
R4526 VSS.t1793 VSS.t1150 2307.56
R4527 VSS.t328 VSS.t1563 2307.56
R4528 VSS.t2380 VSS.t1127 2307.56
R4529 VSS.t1407 VSS.t932 2307.56
R4530 VSS.t935 VSS.t893 2307.56
R4531 VSS.t281 VSS.t729 2307.56
R4532 VSS.t1124 VSS.t2356 2307.56
R4533 VSS.t2384 VSS.t1599 2307.56
R4534 VSS.t990 VSS.t1813 2307.56
R4535 VSS.t1638 VSS.t1817 2307.56
R4536 VSS.n986 VSS.n277 2268.25
R4537 VSS.n1060 VSS.n1059 2220.72
R4538 VSS.n2627 VSS.n2626 2213.34
R4539 VSS.n458 VSS.n393 2212.13
R4540 VSS.n1061 VSS.t2539 2187.61
R4541 VSS.n2494 VSS.t1160 2176.19
R4542 VSS.n1690 VSS.t468 2166.67
R4543 VSS.n0 VSS.t1971 2166.67
R4544 VSS.t1938 VSS.t2316 2159.54
R4545 VSS.n2496 VSS.n2495 2142.66
R4546 VSS.t1329 VSS.t1554 2090.76
R4547 VSS.t2152 VSS.t1584 2090.76
R4548 VSS.t1053 VSS.t1052 2090.76
R4549 VSS.t2548 VSS.t961 2090.76
R4550 VSS.t1457 VSS.n968 2084.8
R4551 VSS.n2599 VSS.n2598 2083.58
R4552 VSS.n603 VSS.n19 2083.1
R4553 VSS.t969 VSS.n576 2050.53
R4554 VSS.n2617 VSS.t964 2050.53
R4555 VSS.n2653 VSS.t1376 1984.24
R4556 VSS.n2497 VSS.n2496 1983.03
R4557 VSS.n1484 VSS.n1483 1982.69
R4558 VSS.n255 VSS.t1624 1964.74
R4559 VSS.n184 VSS.n183 1964.37
R4560 VSS.n3271 VSS.n3269 1946.67
R4561 VSS.n3225 VSS.n3224 1946.67
R4562 VSS.n2552 VSS.t2333 1930.58
R4563 VSS.n1904 VSS.n1901 1925.44
R4564 VSS.n1903 VSS.n1902 1922.83
R4565 VSS.n2555 VSS.n2554 1893.95
R4566 VSS.n2701 VSS.n2700 1890.55
R4567 VSS.n2444 VSS.t1627 1884.89
R4568 VSS.t1605 VSS.n1408 1878.69
R4569 VSS.t604 VSS.n2168 1878.69
R4570 VSS.t1359 VSS.n1588 1878.69
R4571 VSS.t1246 VSS.n814 1862.04
R4572 VSS.n2492 VSS.n2491 1787.45
R4573 VSS.n1209 VSS.n1208 1777.53
R4574 VSS.n1209 VSS.n1207 1777.53
R4575 VSS.n1211 VSS.n1210 1777.53
R4576 VSS.n2980 VSS.n2979 1764.29
R4577 VSS.t1452 VSS.n33 1741.59
R4578 VSS.t1197 VSS.n540 1731.96
R4579 VSS.t2362 VSS.n825 1731.96
R4580 VSS.n3289 VSS.t1669 1719.24
R4581 VSS.t644 VSS.n1836 1719.24
R4582 VSS.t984 VSS.n2237 1719.24
R4583 VSS.t1837 VSS.n1961 1719.24
R4584 VSS.n1387 VSS.t2327 1719.24
R4585 VSS.t816 VSS.n2014 1719.24
R4586 VSS.n2080 VSS.t1309 1719.24
R4587 VSS.t738 VSS.n1818 1719.24
R4588 VSS.n438 VSS.t2346 1719.24
R4589 VSS.n472 VSS.t1408 1719.24
R4590 VSS.t169 VSS.n1309 1713.53
R4591 VSS.n2489 VSS.t1019 1713.53
R4592 VSS.t238 VSS.n2445 1713.53
R4593 VSS.t134 VSS.n2464 1713.53
R4594 VSS.n1956 VSS.t877 1713.53
R4595 VSS.n1441 VSS.t2248 1713.53
R4596 VSS.t366 VSS.n2293 1713.53
R4597 VSS.n2059 VSS.t1131 1713.53
R4598 VSS.t2122 VSS.n2387 1713.53
R4599 VSS.n1661 VSS.t1890 1713.53
R4600 VSS.n1654 VSS.t894 1713.53
R4601 VSS.t1317 VSS.n2629 1713.53
R4602 VSS.n945 VSS.t561 1713.53
R4603 VSS.n522 VSS.n521 1701.86
R4604 VSS.n2253 VSS.n2252 1694.51
R4605 VSS.n1202 VSS.n1201 1678.53
R4606 VSS.n1493 VSS.n1492 1670.2
R4607 VSS.n3058 VSS.n3057 1665.01
R4608 VSS.n1214 VSS.n1212 1659.82
R4609 VSS.t2351 VSS.n3473 1652.1
R4610 VSS.n2616 VSS.t2188 1652.1
R4611 VSS.n3057 VSS.t21 1641.48
R4612 VSS.n1705 VSS.t715 1635.55
R4613 VSS.n8 VSS.t1135 1635.55
R4614 VSS.n1059 VSS.n1058 1620.32
R4615 VSS.n501 VSS.n500 1619.38
R4616 VSS.t732 VSS.n1541 1601.22
R4617 VSS.n3275 VSS.n3274 1598.84
R4618 VSS.n3083 VSS.n3082 1597.63
R4619 VSS.t415 VSS.n55 1587.87
R4620 VSS.n3079 VSS.n311 1573.59
R4621 VSS.n1833 VSS.t1190 1565.03
R4622 VSS.n1309 VSS.n1308 1565.03
R4623 VSS.n3350 VSS.n3289 1565.03
R4624 VSS.n3339 VSS.n104 1565.03
R4625 VSS.n2464 VSS.n2463 1565.03
R4626 VSS.n1442 VSS.n1441 1565.03
R4627 VSS.n2237 VSS.n2236 1565.03
R4628 VSS.n1961 VSS.n1083 1565.03
R4629 VSS.n1387 VSS.n1386 1565.03
R4630 VSS.n2293 VSS.n2292 1565.03
R4631 VSS.n2059 VSS.n1084 1565.03
R4632 VSS.n2387 VSS.n2386 1565.03
R4633 VSS.n2100 VSS.n2080 1565.03
R4634 VSS.n2146 VSS.n2145 1565.03
R4635 VSS.n1655 VSS.n1654 1565.03
R4636 VSS.n1818 VSS.n1817 1565.03
R4637 VSS.n946 VSS.n945 1565.03
R4638 VSS.n441 VSS.n438 1565.03
R4639 VSS.n458 VSS.n457 1565.03
R4640 VSS.n493 VSS.n472 1565.03
R4641 VSS.n2600 VSS.t965 1564.96
R4642 VSS.t249 VSS.n2932 1552.6
R4643 VSS.n1327 VSS.t1746 1544.05
R4644 VSS.n1847 VSS.n1484 1520.16
R4645 VSS.n3368 VSS.t1078 1519.41
R4646 VSS.t208 VSS.n3368 1519.41
R4647 VSS.n3338 VSS.n3316 1493.4
R4648 VSS.t251 VSS.n3451 1490.78
R4649 VSS.t537 VSS.t1779 1483.3
R4650 VSS.t2436 VSS.t575 1483.3
R4651 VSS.t2290 VSS.t759 1483.3
R4652 VSS.t1343 VSS.t2441 1483.3
R4653 VSS.t24 VSS.t1209 1483.3
R4654 VSS.t1186 VSS.t2180 1483.3
R4655 VSS.t751 VSS.t1276 1483.3
R4656 VSS.t1163 VSS.t1274 1483.3
R4657 VSS.t15 VSS.t1975 1479.61
R4658 VSS.n1956 VSS.n1117 1450.79
R4659 VSS.t526 VSS.n773 1441.52
R4660 VSS.n2650 VSS.t540 1439.29
R4661 VSS.n2700 VSS.n2699 1428.64
R4662 VSS.n1774 VSS.n1773 1425.15
R4663 VSS.n3231 VSS.t2437 1419.35
R4664 VSS.n3273 VSS.n221 1418.02
R4665 VSS.n23 VSS.n20 1413.96
R4666 VSS.n3080 VSS.n309 1405.57
R4667 VSS.n346 VSS.n345 1381.04
R4668 VSS.n160 VSS.n159 1379.01
R4669 VSS.n161 VSS.n160 1379.01
R4670 VSS.n162 VSS.n161 1379.01
R4671 VSS.n163 VSS.n162 1379.01
R4672 VSS.n164 VSS.n163 1379.01
R4673 VSS.n165 VSS.n164 1379.01
R4674 VSS.n166 VSS.n165 1379.01
R4675 VSS.n167 VSS.n166 1379.01
R4676 VSS.n168 VSS.n167 1379.01
R4677 VSS.n169 VSS.n168 1379.01
R4678 VSS.n170 VSS.n169 1379.01
R4679 VSS.n171 VSS.n170 1379.01
R4680 VSS.n172 VSS.n171 1379.01
R4681 VSS.n173 VSS.n172 1379.01
R4682 VSS.n174 VSS.n173 1379.01
R4683 VSS.n175 VSS.n174 1379.01
R4684 VSS.n176 VSS.n175 1379.01
R4685 VSS.n177 VSS.n176 1379.01
R4686 VSS.n178 VSS.n177 1379.01
R4687 VSS.n181 VSS.n178 1379.01
R4688 VSS.n182 VSS.n181 1379.01
R4689 VSS.t1536 VSS.t1198 1367.44
R4690 VSS.t795 VSS.t1207 1367.44
R4691 VSS.t911 VSS.n2223 1347.12
R4692 VSS.n3473 VSS.n3472 1333.48
R4693 VSS.n2616 VSS.n2615 1333.48
R4694 VSS.n3420 VSS.t1062 1321.31
R4695 VSS.n1321 VSS.t2413 1313.71
R4696 VSS.n1847 VSS.t2473 1313.03
R4697 VSS.n1744 VSS.n1725 1310.77
R4698 VSS.t276 VSS.t610 1310.38
R4699 VSS.t275 VSS.t648 1310.38
R4700 VSS.t278 VSS.t279 1310.38
R4701 VSS.t648 VSS.t1203 1303.89
R4702 VSS.t279 VSS.t783 1303.89
R4703 VSS.t99 VSS.t358 1303.89
R4704 VSS.n229 VSS.t34 1291.67
R4705 VSS.n3009 VSS.n3008 1282.2
R4706 VSS.n2960 VSS.t692 1272.1
R4707 VSS.n3163 VSS.t438 1272.1
R4708 VSS.n3156 VSS.t1691 1272.1
R4709 VSS.n509 VSS.t1168 1272.1
R4710 VSS.n1070 VSS.t2508 1272.1
R4711 VSS.n822 VSS.t2482 1272.1
R4712 VSS.n2220 VSS.t1557 1272.1
R4713 VSS.n3169 VSS.t1217 1268.89
R4714 VSS.n540 VSS.n539 1249.34
R4715 VSS.n825 VSS.n824 1249.34
R4716 VSS.t2385 VSS.n3443 1228.43
R4717 VSS.n3465 VSS.t538 1226.37
R4718 VSS.n3211 VSS.n229 1216.67
R4719 VSS.n1427 VSS.t2391 1200.91
R4720 VSS.n1869 VSS.t521 1199.47
R4721 VSS.t744 VSS.n3278 1199.47
R4722 VSS.t1466 VSS.n977 1199.47
R4723 VSS.n3168 VSS.t1482 1199.47
R4724 VSS.t1478 VSS.n32 1199.47
R4725 VSS.n3164 VSS.t2203 1199.47
R4726 VSS.n3009 VSS.t263 1199.47
R4727 VSS.n3449 VSS.t266 1199.47
R4728 VSS.n538 VSS.t2166 1199.47
R4729 VSS.n557 VSS.t2123 1199.47
R4730 VSS.n3019 VSS.t258 1199.47
R4731 VSS.n588 VSS.t181 1199.47
R4732 VSS.n3155 VSS.t1462 1199.47
R4733 VSS.n840 VSS.t1409 1199.47
R4734 VSS.n823 VSS.t1682 1199.47
R4735 VSS.n1845 VSS.t2264 1199.47
R4736 VSS.n1836 VSS.n1835 1199.47
R4737 VSS.n2252 VSS.t2407 1199.47
R4738 VSS.n2400 VSS.t1087 1199.47
R4739 VSS.n2221 VSS.t1112 1199.47
R4740 VSS.n1827 VSS.t993 1199.47
R4741 VSS.t203 VSS.n2980 1155.81
R4742 VSS.n1484 VSS.t1047 1153.78
R4743 VSS.t2268 VSS.n1828 1153.78
R4744 VSS.n1057 VSS.t448 1153.78
R4745 VSS.t2349 VSS.n558 1153.78
R4746 VSS.t2192 VSS.n841 1153.78
R4747 VSS.t2319 VSS.n1870 1153.78
R4748 VSS.t991 VSS.n1811 1153.78
R4749 VSS.n3020 VSS.t454 1152.75
R4750 VSS.t2223 VSS.n1978 1147.84
R4751 VSS.t1730 VSS.n1252 1147.84
R4752 VSS.t1895 VSS.n1416 1147.84
R4753 VSS.t2198 VSS.n2176 1147.84
R4754 VSS.t1619 VSS.n1596 1147.84
R4755 VSS.n3474 VSS.t422 1143.48
R4756 VSS.n1711 VSS.t348 1143.48
R4757 VSS.n1722 VSS.n1554 1139.06
R4758 VSS.n504 VSS.n5 1139.06
R4759 VSS.t103 VSS.n684 1134.57
R4760 VSS.t1919 VSS.n893 1134.57
R4761 VSS.n520 VSS.n519 1130.93
R4762 VSS.n3276 VSS.t2531 1124.37
R4763 VSS.n575 VSS.n574 1119.51
R4764 VSS.n2619 VSS.n2618 1119.51
R4765 VSS.n1176 VSS.n1174 1119.51
R4766 VSS.n3389 VSS.t1236 1108.08
R4767 VSS.n1064 VSS.n1063 1102.37
R4768 VSS.n2595 VSS.n2594 1091.42
R4769 VSS.n2493 VSS.n2492 1090.42
R4770 VSS.t757 VSS.n3351 1089.34
R4771 VSS.t1182 VSS.n3391 1089.34
R4772 VSS.n3351 VSS.t225 1086.77
R4773 VSS.n3391 VSS.t220 1086.77
R4774 VSS.n238 VSS.t473 1084.99
R4775 VSS.n3383 VSS.n104 1073.81
R4776 VSS.n461 VSS.n458 1073.81
R4777 VSS.n3451 VSS.n3449 1067.77
R4778 VSS.n1579 VSS.n1578 1062.21
R4779 VSS.t1254 VSS.t2342 1058.09
R4780 VSS.t403 VSS.t2481 1058.09
R4781 VSS.t2177 VSS.n2417 1048.6
R4782 VSS.n3443 VSS.n3442 1043.27
R4783 VSS.n1884 VSS.n1238 1041.81
R4784 VSS.t753 VSS.t958 1040.41
R4785 VSS.t48 VSS.t1303 1040.41
R4786 VSS.t590 VSS.t1077 1040.41
R4787 VSS.t56 VSS.t587 1040.41
R4788 VSS.t1864 VSS.t1181 1040.41
R4789 VSS.t393 VSS.t345 1040.41
R4790 VSS.t614 VSS.t2387 1040.41
R4791 VSS.t1736 VSS.t652 1040.41
R4792 VSS.n2592 VSS.t1940 1035.1
R4793 VSS.n1541 VSS.n1540 1034.55
R4794 VSS.n3421 VSS.n3420 1030.8
R4795 VSS.n1215 VSS.n1209 1023
R4796 VSS.n1215 VSS.n1211 1023
R4797 VSS.t881 VSS.n1321 993.85
R4798 VSS.n635 VSS.n634 988.177
R4799 VSS.n2600 VSS.n910 988.177
R4800 VSS.t1063 VSS.n3421 973.808
R4801 VSS.n22 VSS.n21 960.539
R4802 VSS.t1292 VSS.t1363 952.793
R4803 VSS.t1803 VSS.t617 952.793
R4804 VSS.n1859 VSS.t515 943.548
R4805 VSS.n2254 VSS.n2253 934.764
R4806 VSS.n316 VSS.t565 927.717
R4807 VSS.n1553 VSS.t1447 927.716
R4808 VSS.n330 VSS.t1973 927.716
R4809 VSS.n1215 VSS.n1214 923.559
R4810 VSS.n309 VSS.t45 919.253
R4811 VSS.n230 VSS.t562 919.253
R4812 VSS.n3273 VSS.n186 918.764
R4813 VSS.n2970 VSS.t2164 918.653
R4814 VSS.t2420 VSS.t202 915.494
R4815 VSS.t2315 VSS.t1048 913.885
R4816 VSS.t2467 VSS.t2267 913.885
R4817 VSS.t2461 VSS.t1177 913.885
R4818 VSS.t168 VSS.t880 913.885
R4819 VSS.t1670 VSS.t2535 913.885
R4820 VSS.t421 VSS.t2529 913.885
R4821 VSS.t2282 VSS.t64 913.885
R4822 VSS.t1066 VSS.t416 913.885
R4823 VSS.t1020 VSS.t95 913.885
R4824 VSS.t2262 VSS.t239 913.885
R4825 VSS.t135 VSS.t1629 913.885
R4826 VSS.t1159 VSS.t1625 913.885
R4827 VSS.t2158 VSS.t447 913.885
R4828 VSS.t435 VSS.t2452 913.885
R4829 VSS.t2507 VSS.t1453 913.885
R4830 VSS.t1170 VSS.t1193 913.885
R4831 VSS.t453 VSS.t20 913.885
R4832 VSS.t970 VSS.t1253 913.885
R4833 VSS.t2332 VSS.t1689 913.885
R4834 VSS.t2361 VSS.t2518 913.885
R4835 VSS.t2191 VSS.t2484 913.885
R4836 VSS.t2506 VSS.t1808 913.885
R4837 VSS.t1748 VSS.t2318 913.885
R4838 VSS.t2513 VSS.t643 913.885
R4839 VSS.t2457 VSS.t876 913.885
R4840 VSS.t2489 VSS.t2247 913.885
R4841 VSS.t983 VSS.t2001 913.885
R4842 VSS.t1838 VSS.t1152 913.885
R4843 VSS.t2276 VSS.t2326 913.885
R4844 VSS.t1158 VSS.t536 913.885
R4845 VSS.t2119 VSS.t858 913.885
R4846 VSS.t367 VSS.t684 913.885
R4847 VSS.t2112 VSS.t1130 913.885
R4848 VSS.t2121 VSS.t2536 913.885
R4849 VSS.t817 VSS.t1556 913.885
R4850 VSS.t2205 VSS.t1308 913.885
R4851 VSS.t1228 VSS.t568 913.885
R4852 VSS.t2212 VSS.t1072 913.885
R4853 VSS.t1891 VSS.t872 913.885
R4854 VSS.t895 VSS.t1320 913.885
R4855 VSS.t542 VSS.t1316 913.885
R4856 VSS.t2480 VSS.t963 913.885
R4857 VSS.t2232 VSS.t737 913.885
R4858 VSS.t2241 VSS.t992 913.885
R4859 VSS.t747 VSS.t696 913.885
R4860 VSS.t560 VSS.t699 913.885
R4861 VSS.t2534 VSS.t2347 913.885
R4862 VSS.t2304 VSS.t2519 913.885
R4863 VSS.t1119 VSS.t1407 913.885
R4864 VSS.t1117 VSS.t2384 913.885
R4865 VSS.n2629 VSS.n2628 902.461
R4866 VSS.t1369 VSS.t727 887.163
R4867 VSS.t1378 VSS.t2543 887.163
R4868 VSS.n316 VSS.n235 879.836
R4869 VSS.n2495 VSS.n2494 864.766
R4870 VSS.n963 VSS.n962 863.635
R4871 VSS.n2588 VSS.n2587 862.682
R4872 VSS.n1220 VSS.n1204 860
R4873 VSS.t2316 VSS.t1749 855.264
R4874 VSS.n2554 VSS.n2553 843.75
R4875 VSS.n2628 VSS.n2627 839.713
R4876 VSS.n1984 VSS.t58 838.187
R4877 VSS.n1259 VSS.t290 838.187
R4878 VSS.n1364 VSS.t1677 838.187
R4879 VSS.n2147 VSS.t1945 838.187
R4880 VSS.n1619 VSS.t581 838.187
R4881 VSS.n494 VSS.t1853 836.591
R4882 VSS.n2542 VSS.t2550 833.202
R4883 VSS.t2027 VSS.t1880 828.027
R4884 VSS.t445 VSS.t2152 828.027
R4885 VSS.t2071 VSS.t173 828.027
R4886 VSS.t443 VSS.t2548 828.027
R4887 VSS.n1220 VSS.n1219 822.424
R4888 VSS.t1404 VSS.t1525 794.981
R4889 VSS.n507 VSS.n505 791.109
R4890 VSS.n1724 VSS.n1723 791.109
R4891 VSS.t152 VSS.t1184 784.35
R4892 VSS.t1746 VSS.n1240 782.221
R4893 VSS.t1562 VSS.t296 779.128
R4894 VSS.n1536 VSS.t2271 776.83
R4895 VSS.n973 VSS.t2149 776.83
R4896 VSS.n405 VSS.t1073 776.83
R4897 VSS.n651 VSS.t2375 776.83
R4898 VSS.n2574 VSS.t1941 776.83
R4899 VSS.n1919 VSS.t2220 776.83
R4900 VSS.n3082 VSS.t1728 771.441
R4901 VSS.n1885 VSS.n1884 763.912
R4902 VSS.n397 VSS.t857 760.976
R4903 VSS.n643 VSS.t2360 760.976
R4904 VSS.n2627 VSS.n814 756.466
R4905 VSS.t1388 VSS.n1862 754.639
R4906 VSS.n234 VSS.t1985 753.193
R4907 VSS.n1218 VSS.n1217 748.63
R4908 VSS.n3273 VSS.n3272 742.952
R4909 VSS.t2521 VSS.n1833 742.532
R4910 VSS.n3155 VSS.n281 738.636
R4911 VSS.n2401 VSS.n2400 738.636
R4912 VSS.n674 VSS.n673 730.396
R4913 VSS.n556 VSS.t1251 730.073
R4914 VSS.n839 VSS.t2494 730.073
R4915 VSS.n3080 VSS.t5 709.049
R4916 VSS.n1868 VSS.t2313 699.654
R4917 VSS.n2553 VSS.n2552 685.413
R4918 VSS.t451 VSS.n19 681.269
R4919 VSS.t1411 VSS.n788 680.952
R4920 VSS.n3212 VSS.n3211 676.096
R4921 VSS.n3081 VSS.n235 673.139
R4922 VSS.n1979 VSS.t2223 671.942
R4923 VSS.n1277 VSS.t1730 671.942
R4924 VSS.n2418 VSS.t2177 671.942
R4925 VSS.n1417 VSS.t1895 671.942
R4926 VSS.n2177 VSS.t2198 671.942
R4927 VSS.n1597 VSS.t1619 671.942
R4928 VSS.n1238 VSS.t511 668.119
R4929 VSS.n909 VSS.t2186 663.793
R4930 VSS.n636 VSS.t2353 663.793
R4931 VSS.n3276 VSS.n3275 663.732
R4932 VSS.n1845 VSS.n773 663.091
R4933 VSS.t610 VSS.n3230 655.191
R4934 VSS.n3269 VSS.t99 655.191
R4935 VSS.t2317 VSS.n1860 650.643
R4936 VSS.n2622 VSS.n2621 650.433
R4937 VSS.n3471 VSS.t273 643.692
R4938 VSS.t832 VSS.t1783 635.715
R4939 VSS.t1894 VSS.t1361 635.715
R4940 VSS.n894 VSS.t2498 631.266
R4941 VSS.n296 VSS.n295 629.365
R4942 VSS.n3115 VSS.n3114 629.365
R4943 VSS.t1355 VSS.n1143 627.63
R4944 VSS.n1198 VSS.t1345 627.63
R4945 VSS.n293 VSS.n292 626.053
R4946 VSS.n3107 VSS.n3106 626.053
R4947 VSS.t150 VSS.t790 624.697
R4948 VSS.n3443 VSS.n32 620.379
R4949 VSS.n117 VSS.n116 619.048
R4950 VSS.n3085 VSS.n3084 616.962
R4951 VSS.n3091 VSS.n3090 616.962
R4952 VSS.n303 VSS.n302 615.048
R4953 VSS.n3099 VSS.n3098 615.048
R4954 VSS.n2958 VSS.t583 601.938
R4955 VSS.n2949 VSS.t84 601.938
R4956 VSS.n2965 VSS.t810 600.457
R4957 VSS.n2038 VSS.t2210 596.681
R4958 VSS.n2101 VSS.t1226 596.681
R4959 VSS.n2124 VSS.t487 596.681
R4960 VSS.n2598 VSS.n2597 596.27
R4961 VSS.n910 VSS.t558 596.024
R4962 VSS.t2245 VSS.n635 596.024
R4963 VSS.t1107 VSS.n2038 595.269
R4964 VSS.t1104 VSS.n2101 595.269
R4965 VSS.n2124 VSS.t1096 595.269
R4966 VSS.n2492 VSS.n2489 588.769
R4967 VSS.n2445 VSS.n1064 582.601
R4968 VSS.n504 VSS.t1134 578.554
R4969 VSS.n1722 VSS.t1733 578.554
R4970 VSS.n2556 VSS.t1697 577.351
R4971 VSS.n3218 VSS.n229 576.442
R4972 VSS.n440 VSS.t2102 574.562
R4973 VSS.t1442 VSS.t2216 569.879
R4974 VSS.t628 VSS.t1959 569.879
R4975 VSS.t1702 VSS.t1227 569.879
R4976 VSS.t1356 VSS.t612 569.879
R4977 VSS.t1422 VSS.t491 569.879
R4978 VSS.t1139 VSS.t1137 569.879
R4979 VSS.t887 VSS.t1824 569.879
R4980 VSS.t2096 VSS.t330 569.879
R4981 VSS.n2554 VSS.n968 567.962
R4982 VSS.n3442 VSS.t2449 565.933
R4983 VSS.n787 VSS.t874 564.287
R4984 VSS.n1536 VSS.t1365 554.879
R4985 VSS.t1796 VSS.n973 554.879
R4986 VSS.n405 VSS.t75 554.879
R4987 VSS.n651 VSS.t2226 554.879
R4988 VSS.t769 VSS.n2574 554.879
R4989 VSS.n1919 VSS.t199 554.879
R4990 VSS.t218 VSS.n3194 553.516
R4991 VSS.n2981 VSS.t203 549.297
R4992 VSS.n2986 VSS.t2131 549.297
R4993 VSS.n2987 VSS.t1566 549.297
R4994 VSS.n2991 VSS.t2420 549.297
R4995 VSS.n1904 VSS.n1903 548.634
R4996 VSS.t1047 VSS.n1481 548.331
R4997 VSS.n1472 VSS.t1058 548.331
R4998 VSS.n1473 VSS.t2315 548.331
R4999 VSS.n1832 VSS.t2467 548.331
R5000 VSS.n1831 VSS.t1900 548.331
R5001 VSS.n1830 VSS.t1952 548.331
R5002 VSS.n1829 VSS.t2268 548.331
R5003 VSS.n1983 VSS.t2012 548.331
R5004 VSS.n1985 VSS.t685 548.331
R5005 VSS.n1987 VSS.t2011 548.331
R5006 VSS.n1258 VSS.t1036 548.331
R5007 VSS.n1260 VSS.t886 548.331
R5008 VSS.n1262 VSS.t1039 548.331
R5009 VSS.n1295 VSS.t1176 548.331
R5010 VSS.n1296 VSS.t97 548.331
R5011 VSS.n1301 VSS.t231 548.331
R5012 VSS.n1302 VSS.t2461 548.331
R5013 VSS.n1312 VSS.t169 548.331
R5014 VSS.n1313 VSS.t1284 548.331
R5015 VSS.n1320 VSS.t880 548.331
R5016 VSS.t483 VSS.n3283 548.331
R5017 VSS.n3284 VSS.t49 548.331
R5018 VSS.t1669 VSS.n3288 548.331
R5019 VSS.n3348 VSS.t2488 548.331
R5020 VSS.t1438 VSS.n3295 548.331
R5021 VSS.t57 VSS.n3297 548.331
R5022 VSS.n3340 VSS.t742 548.331
R5023 VSS.t2529 VSS.n980 548.331
R5024 VSS.t951 VSS.n982 548.331
R5025 VSS.t336 VSS.n984 548.331
R5026 VSS.n988 VSS.t420 548.331
R5027 VSS.n276 VSS.t2282 548.331
R5028 VSS.n275 VSS.t1756 548.331
R5029 VSS.t1535 VSS.n267 548.331
R5030 VSS.n269 VSS.t65 548.331
R5031 VSS.n58 VSS.t415 548.331
R5032 VSS.n59 VSS.t1646 548.331
R5033 VSS.n64 VSS.t1739 548.331
R5034 VSS.n65 VSS.t1066 548.331
R5035 VSS.t1019 VSS.n2488 548.331
R5036 VSS.t2254 VSS.n2487 548.331
R5037 VSS.t794 VSS.n2486 548.331
R5038 VSS.t95 VSS.n2485 548.331
R5039 VSS.n2448 VSS.t238 548.331
R5040 VSS.n2449 VSS.t299 548.331
R5041 VSS.n2454 VSS.t193 548.331
R5042 VSS.n2455 VSS.t2262 548.331
R5043 VSS.n2467 VSS.t134 548.331
R5044 VSS.n2468 VSS.t110 548.331
R5045 VSS.n2471 VSS.t1419 548.331
R5046 VSS.n2476 VSS.t1629 548.331
R5047 VSS.n2430 VSS.t1336 548.331
R5048 VSS.n2433 VSS.t2259 548.331
R5049 VSS.n2435 VSS.t1335 548.331
R5050 VSS.n1005 VSS.t1164 548.331
R5051 VSS.n1010 VSS.t1022 548.331
R5052 VSS.n1011 VSS.t472 548.331
R5053 VSS.n1016 VSS.t1625 548.331
R5054 VSS.t448 VSS.n1029 548.331
R5055 VSS.t1828 VSS.n1028 548.331
R5056 VSS.t1613 VSS.n1027 548.331
R5057 VSS.n1022 VSS.t2158 548.331
R5058 VSS.t2201 VSS.n1056 548.331
R5059 VSS.t1330 VSS.n1055 548.331
R5060 VSS.t1298 VSS.n1054 548.331
R5061 VSS.n1049 VSS.t444 548.331
R5062 VSS.t2451 VSS.n1046 548.331
R5063 VSS.t1051 VSS.n1045 548.331
R5064 VSS.n1039 VSS.t435 548.331
R5065 VSS.n3007 VSS.t2507 548.331
R5066 VSS.t1700 VSS.n2998 548.331
R5067 VSS.n3000 VSS.t1452 548.331
R5068 VSS.t538 VSS.n3464 548.331
R5069 VSS.n26 VSS.t678 548.331
R5070 VSS.n27 VSS.t551 548.331
R5071 VSS.n28 VSS.t1162 548.331
R5072 VSS.n526 VSS.t1860 548.331
R5073 VSS.n531 VSS.t1368 548.331
R5074 VSS.n532 VSS.t1380 548.331
R5075 VSS.n537 VSS.t1257 548.331
R5076 VSS.n541 VSS.t1197 548.331
R5077 VSS.n547 VSS.t1396 548.331
R5078 VSS.n548 VSS.t2104 548.331
R5079 VSS.n551 VSS.t1170 548.331
R5080 VSS.t21 VSS.n3056 548.331
R5081 VSS.t457 VSS.n3055 548.331
R5082 VSS.n3017 VSS.t1926 548.331
R5083 VSS.n3018 VSS.t453 548.331
R5084 VSS.n559 VSS.t2349 548.331
R5085 VSS.n565 VSS.t54 548.331
R5086 VSS.n566 VSS.t1282 548.331
R5087 VSS.n569 VSS.t1248 548.331
R5088 VSS.n577 VSS.t969 548.331
R5089 VSS.n582 VSS.t1523 548.331
R5090 VSS.n583 VSS.t1855 548.331
R5091 VSS.n587 VSS.t1253 548.331
R5092 VSS.t2333 VSS.n2551 548.331
R5093 VSS.n2544 VSS.t2141 548.331
R5094 VSS.n3154 VSS.t1689 548.331
R5095 VSS.n826 VSS.t2362 548.331
R5096 VSS.n831 VSS.t1781 548.331
R5097 VSS.n832 VSS.t1723 548.331
R5098 VSS.n837 VSS.t2518 548.331
R5099 VSS.n842 VSS.t2192 548.331
R5100 VSS.n847 VSS.t1765 548.331
R5101 VSS.n848 VSS.t1673 548.331
R5102 VSS.n853 VSS.t2484 548.331
R5103 VSS.t1807 VSS.n2698 548.331
R5104 VSS.n774 VSS.t1364 548.331
R5105 VSS.n775 VSS.t2309 548.331
R5106 VSS.n776 VSS.t2506 548.331
R5107 VSS.n1871 VSS.t2319 548.331
R5108 VSS.n1876 VSS.t2320 548.331
R5109 VSS.n1877 VSS.t1392 548.331
R5110 VSS.n1882 VSS.t1748 548.331
R5111 VSS.n1844 VSS.t2513 548.331
R5112 VSS.n1843 VSS.t660 548.331
R5113 VSS.t1353 VSS.n1490 548.331
R5114 VSS.n1837 VSS.t644 548.331
R5115 VSS.t877 VSS.n1955 548.331
R5116 VSS.n1118 VSS.t2466 548.331
R5117 VSS.n1119 VSS.t156 548.331
R5118 VSS.n1120 VSS.t2457 548.331
R5119 VSS.t2248 VSS.n1440 548.331
R5120 VSS.n1354 VSS.t1763 548.331
R5121 VSS.n1355 VSS.t1520 548.331
R5122 VSS.n1356 VSS.t2489 548.331
R5123 VSS.t2001 VSS.n2226 548.331
R5124 VSS.t1264 VSS.n2228 548.331
R5125 VSS.t2005 VSS.n2230 548.331
R5126 VSS.n2238 VSS.t984 548.331
R5127 VSS.t1152 VSS.n1111 548.331
R5128 VSS.t2185 VSS.n1113 548.331
R5129 VSS.t1964 VSS.n1115 548.331
R5130 VSS.n1962 VSS.t1837 548.331
R5131 VSS.n2331 VSS.t2276 548.331
R5132 VSS.n2330 VSS.t118 548.331
R5133 VSS.n2329 VSS.t943 548.331
R5134 VSS.n1384 VSS.t1158 548.331
R5135 VSS.n1383 VSS.t19 548.331
R5136 VSS.n1382 VSS.t427 548.331
R5137 VSS.n1381 VSS.t535 548.331
R5138 VSS.n1095 VSS.t859 548.331
R5139 VSS.n1096 VSS.t909 548.331
R5140 VSS.n1101 VSS.t1716 548.331
R5141 VSS.n1102 VSS.t2119 548.331
R5142 VSS.n2296 VSS.t366 548.331
R5143 VSS.n2297 VSS.t1839 548.331
R5144 VSS.n2300 VSS.t307 548.331
R5145 VSS.n2304 VSS.t684 548.331
R5146 VSS.t1131 VSS.n2058 548.331
R5147 VSS.t1774 VSS.n2057 548.331
R5148 VSS.n2050 VSS.t66 548.331
R5149 VSS.n2051 VSS.t2112 548.331
R5150 VSS.n2390 VSS.t2122 548.331
R5151 VSS.n2391 VSS.t813 548.331
R5152 VSS.n2394 VSS.t789 548.331
R5153 VSS.n2399 VSS.t2536 548.331
R5154 VSS.t1556 VSS.n2008 548.331
R5155 VSS.t635 VSS.n2010 548.331
R5156 VSS.t1960 VSS.n2012 548.331
R5157 VSS.n2015 VSS.t816 548.331
R5158 VSS.n2070 VSS.t2205 548.331
R5159 VSS.t1387 VSS.n2074 548.331
R5160 VSS.n2075 VSS.t613 548.331
R5161 VSS.t1309 VSS.n2079 548.331
R5162 VSS.n2098 VSS.t1228 548.331
R5163 VSS.n2097 VSS.t1545 548.331
R5164 VSS.n2096 VSS.t1138 548.331
R5165 VSS.n2095 VSS.t569 548.331
R5166 VSS.n2143 VSS.t2212 548.331
R5167 VSS.n2142 VSS.t2328 548.331
R5168 VSS.n2141 VSS.t331 548.331
R5169 VSS.n2140 VSS.t1071 548.331
R5170 VSS.t1890 VSS.n1660 548.331
R5171 VSS.t831 VSS.n1659 548.331
R5172 VSS.t1575 VSS.n1658 548.331
R5173 VSS.t872 VSS.n1657 548.331
R5174 VSS.t894 VSS.n1653 548.331
R5175 VSS.t396 VSS.n1652 548.331
R5176 VSS.t1996 VSS.n1651 548.331
R5177 VSS.t1320 VSS.n1650 548.331
R5178 VSS.n2632 VSS.t1317 548.331
R5179 VSS.n2633 VSS.t544 548.331
R5180 VSS.n2638 VSS.t1827 548.331
R5181 VSS.n2639 VSS.t542 548.331
R5182 VSS.n881 VSS.t964 548.331
R5183 VSS.n882 VSS.t1547 548.331
R5184 VSS.n887 VSS.t837 548.331
R5185 VSS.n888 VSS.t2480 548.331
R5186 VSS.n1826 VSS.t2232 548.331
R5187 VSS.n1825 VSS.t927 548.331
R5188 VSS.t362 VSS.n1511 548.331
R5189 VSS.n1819 VSS.t738 548.331
R5190 VSS.n1815 VSS.t2241 548.331
R5191 VSS.n1814 VSS.t1511 548.331
R5192 VSS.n1813 VSS.t351 548.331
R5193 VSS.n1812 VSS.t991 548.331
R5194 VSS.n921 VSS.t750 548.331
R5195 VSS.n922 VSS.t704 548.331
R5196 VSS.n925 VSS.t160 548.331
R5197 VSS.n930 VSS.t696 548.331
R5198 VSS.t561 VSS.n944 548.331
R5199 VSS.t2093 VSS.n943 548.331
R5200 VSS.t188 VSS.n942 548.331
R5201 VSS.t699 VSS.n941 548.331
R5202 VSS.n428 VSS.t2534 548.331
R5203 VSS.t1930 VSS.n432 548.331
R5204 VSS.n433 VSS.t1640 548.331
R5205 VSS.t2346 VSS.n437 548.331
R5206 VSS.t2519 VSS.n448 548.331
R5207 VSS.n452 VSS.t328 548.331
R5208 VSS.t2370 VSS.n456 548.331
R5209 VSS.n462 VSS.t1119 548.331
R5210 VSS.t893 VSS.n466 548.331
R5211 VSS.n467 VSS.t281 548.331
R5212 VSS.t1408 VSS.n471 548.331
R5213 VSS.n491 VSS.t1117 548.331
R5214 VSS.n490 VSS.t990 548.331
R5215 VSS.n489 VSS.t1638 548.331
R5216 VSS.n488 VSS.t2383 548.331
R5217 VSS.n2511 VSS.t2549 546.41
R5218 VSS.n2578 VSS.t284 546.41
R5219 VSS.n1911 VSS.t502 546.41
R5220 VSS.n1528 VSS.t1189 546.41
R5221 VSS.n502 VSS.n501 545.501
R5222 VSS.n2621 VSS.n2620 545.501
R5223 VSS.t2242 VSS.n1506 522.021
R5224 VSS.t1210 VSS.t276 518.962
R5225 VSS.t1206 VSS.t275 518.962
R5226 VSS.t1208 VSS.t278 518.962
R5227 VSS.n1466 VSS.t2034 513.159
R5228 VSS.n1960 VSS.n1958 508.851
R5229 VSS.n2063 VSS.n2061 508.851
R5230 VSS.n1061 VSS.n1060 508.697
R5231 VSS.n397 VSS.t2500 507.317
R5232 VSS.n643 VSS.t1120 507.317
R5233 VSS.n688 VSS.t987 503.682
R5234 VSS.n2522 VSS.t1329 496.815
R5235 VSS.n2526 VSS.t2027 496.815
R5236 VSS.n2527 VSS.t445 496.815
R5237 VSS.t2550 VSS.n2541 496.815
R5238 VSS.t1052 VSS.n2540 496.815
R5239 VSS.n2533 VSS.t2071 496.815
R5240 VSS.n2534 VSS.t443 496.815
R5241 VSS.n3135 VSS.t669 485.95
R5242 VSS.n298 VSS.n296 484.921
R5243 VSS.t939 VSS.t2269 480.776
R5244 VSS.t1024 VSS.t1354 480.074
R5245 VSS.t430 VSS.n1979 479.959
R5246 VSS.n1277 VSS.t460 479.959
R5247 VSS.n2418 VSS.t2009 479.959
R5248 VSS.n1417 VSS.t370 479.959
R5249 VSS.n2177 VSS.t1499 479.959
R5250 VSS.n1597 VSS.t1772 479.959
R5251 VSS.n1835 VSS.n1834 479.789
R5252 VSS.t440 VSS.t760 470.442
R5253 VSS.t1829 VSS.t428 470.442
R5254 VSS.n2700 VSS.t1806 470.426
R5255 VSS.t1015 VSS.n1575 470.426
R5256 VSS.n3084 VSS.n3083 468.62
R5257 VSS.n1222 VSS.n1221 459.906
R5258 VSS.t2395 VSS.n1242 458.837
R5259 VSS.t136 VSS.t552 457.144
R5260 VSS.n300 VSS.n293 455
R5261 VSS.n576 VSS.n575 453.219
R5262 VSS.n2618 VSS.n2617 453.219
R5263 VSS.n1662 VSS.n1661 451.231
R5264 VSS.n3091 VSS.n306 448.392
R5265 VSS.t1318 VSS.n814 445.519
R5266 VSS.n1923 VSS.n914 444.738
R5267 VSS.n23 VSS.n22 443.99
R5268 VSS.n1783 VSS.t507 442.755
R5269 VSS.t1285 VSS.n1760 442.75
R5270 VSS.t921 VSS.t503 441.493
R5271 VSS.n788 VSS.n787 440.476
R5272 VSS.n673 VSS.n672 439.236
R5273 VSS.t98 VSS.t626 438.545
R5274 VSS.t1833 VSS.t944 438.545
R5275 VSS.t166 VSS.t1283 438.106
R5276 VSS.t1034 VSS.t1751 438.106
R5277 VSS.t2429 VSS.t2136 434.212
R5278 VSS.t1846 VSS.t2368 434.212
R5279 VSS.n55 VSS.n52 434.096
R5280 VSS.t2013 VSS.t2435 433.334
R5281 VSS.t682 VSS.t2274 433.334
R5282 VSS.t2120 VSS.t1083 433.334
R5283 VSS.t1588 VSS.t218 432.336
R5284 VSS.n208 VSS.n207 431.777
R5285 VSS.n209 VSS.n208 431.777
R5286 VSS.n210 VSS.n209 431.777
R5287 VSS.n211 VSS.n210 431.777
R5288 VSS.n212 VSS.n211 431.777
R5289 VSS.n213 VSS.n212 431.777
R5290 VSS.n214 VSS.n213 431.777
R5291 VSS.n215 VSS.n214 431.777
R5292 VSS.n216 VSS.n215 431.777
R5293 VSS.n217 VSS.n216 431.777
R5294 VSS.n218 VSS.n217 431.777
R5295 VSS.n302 VSS.n301 430.197
R5296 VSS.n3099 VSS.n301 426.837
R5297 VSS.n539 VSS.n538 426.769
R5298 VSS.n824 VSS.n823 426.769
R5299 VSS.n857 VSS.t913 426.396
R5300 VSS.n617 VSS.t1579 426.396
R5301 VSS.t247 VSS.n947 425.094
R5302 VSS.n221 VSS.n220 425.05
R5303 VSS.n947 VSS.t287 424.089
R5304 VSS.t361 VSS.t663 422.866
R5305 VSS.t119 VSS.t2219 422.866
R5306 VSS.n2444 VSS.t916 422.671
R5307 VSS.n1327 VSS.n1326 418.692
R5308 VSS.t298 VSS.t2250 416.635
R5309 VSS.t1567 VSS.t1232 414.719
R5310 VSS.n2412 VSS.n222 412.745
R5311 VSS.n3261 VSS.n3226 412.745
R5312 VSS.t2497 VSS.t753 412.045
R5313 VSS.t2068 VSS.t1530 412.045
R5314 VSS.t1077 VSS.t2479 412.045
R5315 VSS.t2069 VSS.t1434 412.045
R5316 VSS.t1181 VSS.t1240 412.045
R5317 VSS.t2079 VSS.t1875 412.045
R5318 VSS.t2387 VSS.t1239 412.045
R5319 VSS.t2037 VSS.t1313 412.045
R5320 VSS.t705 VSS.t1961 406
R5321 VSS.t2092 VSS.t380 406
R5322 VSS.t397 VSS.t340 405.356
R5323 VSS.t1671 VSS.t1999 405.356
R5324 VSS.t871 VSS.t765 405.356
R5325 VSS.t1749 VSS.n1238 400.906
R5326 VSS.n3420 VSS.n68 399.878
R5327 VSS.t1081 VSS.t1767 398.623
R5328 VSS.t492 VSS.t724 398.623
R5329 VSS.t1322 VSS.t1503 398.623
R5330 VSS.t806 VSS.t456 398.241
R5331 VSS.n12 VSS.t1132 396.058
R5332 VSS.t1734 VSS.n1717 396.058
R5333 VSS.n1463 VSS.t1035 394.728
R5334 VSS.n2510 VSS.n2509 390.582
R5335 VSS.t523 VSS.n1784 386.233
R5336 VSS.n1587 VSS.n1579 383.952
R5337 VSS.t1327 VSS.t871 381.512
R5338 VSS.t543 VSS.t1321 380.952
R5339 VSS.t557 VSS.t1376 380.952
R5340 VSS.t679 VSS.t706 379.551
R5341 VSS.n1572 VSS.t1892 373.81
R5342 VSS.t2515 VSS.n3012 372.873
R5343 VSS.t2049 VSS.t1935 370.132
R5344 VSS.t2471 VSS.t2108 370.132
R5345 VSS.t2017 VSS.t2018 367.89
R5346 VSS.t191 VSS.t452 367.142
R5347 VSS.n2981 VSS.t2344 366.197
R5348 VSS.t1230 VSS.n2986 366.197
R5349 VSS.t253 VSS.n2991 366.197
R5350 VSS.n1481 VSS.t1661 365.555
R5351 VSS.t1055 VSS.n1471 365.555
R5352 VSS.t1049 VSS.n1472 365.555
R5353 VSS.n1473 VSS.t521 365.555
R5354 VSS.t1190 VSS.n1832 365.555
R5355 VSS.t1492 VSS.n1831 365.555
R5356 VSS.t1901 VSS.n1830 365.555
R5357 VSS.t1953 VSS.n1829 365.555
R5358 VSS.n1983 VSS.t2114 365.555
R5359 VSS.t2014 VSS.n1985 365.555
R5360 VSS.n1987 VSS.t680 365.555
R5361 VSS.n1258 VSS.t2459 365.555
R5362 VSS.t1037 VSS.n1260 365.555
R5363 VSS.n1262 VSS.t878 365.555
R5364 VSS.t2193 VSS.n1295 365.555
R5365 VSS.n1296 VSS.t228 365.555
R5366 VSS.t850 VSS.n1301 365.555
R5367 VSS.n1302 VSS.t848 365.555
R5368 VSS.t1867 VSS.n1312 365.555
R5369 VSS.n1313 VSS.t432 365.555
R5370 VSS.n1316 VSS.t946 365.555
R5371 VSS.t2413 VSS.n1320 365.555
R5372 VSS.n3279 VSS.t744 365.555
R5373 VSS.n3283 VSS.t302 365.555
R5374 VSS.n3284 VSS.t1531 365.555
R5375 VSS.n3288 VSS.t818 365.555
R5376 VSS.t754 VSS.n3348 365.555
R5377 VSS.n3295 VSS.t1788 365.555
R5378 VSS.n3297 VSS.t1435 365.555
R5379 VSS.n3340 VSS.t762 365.555
R5380 VSS.n980 VSS.t1466 365.555
R5381 VSS.n982 VSS.t325 365.555
R5382 VSS.n984 VSS.t1551 365.555
R5383 VSS.n988 VSS.t337 365.555
R5384 VSS.t1482 VSS.n276 365.555
R5385 VSS.t1277 VSS.n275 365.555
R5386 VSS.n267 VSS.t1870 365.555
R5387 VSS.n269 VSS.t1686 365.555
R5388 VSS.t661 VSS.n58 365.555
R5389 VSS.n59 VSS.t1968 365.555
R5390 VSS.t22 VSS.n64 365.555
R5391 VSS.n65 VSS.t1478 365.555
R5392 VSS.n2488 VSS.t387 365.555
R5393 VSS.n2487 VSS.t948 365.555
R5394 VSS.n2486 VSS.t975 365.555
R5395 VSS.n2485 VSS.t204 365.555
R5396 VSS.t300 VSS.n2448 365.555
R5397 VSS.n2449 VSS.t197 365.555
R5398 VSS.t240 VSS.n2454 365.555
R5399 VSS.n2455 VSS.t216 365.555
R5400 VSS.t88 VSS.n2467 365.555
R5401 VSS.n2468 VSS.t1416 365.555
R5402 VSS.n2471 VSS.t1268 365.555
R5403 VSS.t1160 VSS.n2476 365.555
R5404 VSS.n2430 VSS.t1627 365.555
R5405 VSS.t1338 VSS.n2433 365.555
R5406 VSS.n2435 VSS.t2257 365.555
R5407 VSS.n1005 VSS.t1992 365.555
R5408 VSS.t474 VSS.n1010 365.555
R5409 VSS.n1011 VSS.t2541 365.555
R5410 VSS.t2539 VSS.n1016 365.555
R5411 VSS.n1029 VSS.t10 365.555
R5412 VSS.n1028 VSS.t1611 365.555
R5413 VSS.n1022 VSS.t1457 365.555
R5414 VSS.n1056 VSS.t1331 365.555
R5415 VSS.n1055 VSS.t1878 365.555
R5416 VSS.n1054 VSS.t639 365.555
R5417 VSS.n1049 VSS.t2546 365.555
R5418 VSS.n1046 VSS.t1400 365.555
R5419 VSS.n1045 VSS.t174 365.555
R5420 VSS.t354 VSS.n1038 365.555
R5421 VSS.n1039 VSS.t2203 365.555
R5422 VSS.t263 VSS.n3007 365.555
R5423 VSS.t1527 VSS.n3006 365.555
R5424 VSS.n2998 VSS.t1705 365.555
R5425 VSS.n3000 VSS.t1711 365.555
R5426 VSS.n3464 VSS.t711 365.555
R5427 VSS.t709 VSS.n26 365.555
R5428 VSS.n27 VSS.t1663 365.555
R5429 VSS.t266 VSS.n28 365.555
R5430 VSS.n526 VSS.t1586 365.555
R5431 VSS.t2544 VSS.n531 365.555
R5432 VSS.n532 VSS.t2170 365.555
R5433 VSS.t2166 VSS.n537 365.555
R5434 VSS.n541 VSS.t1333 365.555
R5435 VSS.t2100 VSS.n547 365.555
R5436 VSS.n548 VSS.t1432 365.555
R5437 VSS.n551 VSS.t2123 365.555
R5438 VSS.n3056 VSS.t40 365.555
R5439 VSS.t1370 VSS.n3017 365.555
R5440 VSS.t258 VSS.n3018 365.555
R5441 VSS.n559 VSS.t602 365.555
R5442 VSS.t2139 VSS.n565 365.555
R5443 VSS.n566 VSS.t2321 365.555
R5444 VSS.n569 VSS.t2366 365.555
R5445 VSS.n577 VSS.t1990 365.555
R5446 VSS.t1857 VSS.n582 365.555
R5447 VSS.n583 VSS.t130 365.555
R5448 VSS.t181 VSS.n587 365.555
R5449 VSS.n2551 VSS.t2154 365.555
R5450 VSS.t2143 VSS.n2543 365.555
R5451 VSS.n2544 VSS.t1695 365.555
R5452 VSS.t1462 VSS.n3154 365.555
R5453 VSS.n826 VSS.t466 365.555
R5454 VSS.t829 VSS.n831 365.555
R5455 VSS.n832 VSS.t2086 365.555
R5456 VSS.t1409 VSS.n837 365.555
R5457 VSS.n842 VSS.t2090 365.555
R5458 VSS.t1675 VSS.n847 365.555
R5459 VSS.n848 VSS.t1709 365.555
R5460 VSS.t2307 VSS.n853 365.555
R5461 VSS.n2698 VSS.t901 365.555
R5462 VSS.t1786 VSS.n774 365.555
R5463 VSS.t1988 VSS.n775 365.555
R5464 VSS.t1682 VSS.n776 365.555
R5465 VSS.n1871 VSS.t1294 365.555
R5466 VSS.t1394 VSS.n1876 365.555
R5467 VSS.n1877 VSS.t981 365.555
R5468 VSS.t517 VSS.n1882 365.555
R5469 VSS.t2264 VSS.n1844 365.555
R5470 VSS.t645 VSS.n1843 365.555
R5471 VSS.n1490 VSS.t653 365.555
R5472 VSS.n1837 VSS.t799 365.555
R5473 VSS.n1955 VSS.t1495 365.555
R5474 VSS.t841 VSS.n1118 365.555
R5475 VSS.t476 VSS.n1119 365.555
R5476 VSS.t1174 VSS.n1120 365.555
R5477 VSS.n1440 VSS.t373 365.555
R5478 VSS.t1799 VSS.n1354 365.555
R5479 VSS.t1873 VSS.n1355 365.555
R5480 VSS.t2391 VSS.n1356 365.555
R5481 VSS.n2226 VSS.t2407 365.555
R5482 VSS.n2228 VSS.t37 365.555
R5483 VSS.n2230 VSS.t599 365.555
R5484 VSS.n2238 VSS.t1881 365.555
R5485 VSS.n1111 VSS.t532 365.555
R5486 VSS.n1113 VSS.t1916 365.555
R5487 VSS.n1115 VSS.t929 365.555
R5488 VSS.n1962 VSS.t1965 365.555
R5489 VSS.t2397 VSS.n2331 365.555
R5490 VSS.t546 VSS.n2330 365.555
R5491 VSS.t1720 VSS.n2329 365.555
R5492 VSS.t2127 VSS.n2328 365.555
R5493 VSS.t69 VSS.n1384 365.555
R5494 VSS.t72 VSS.n1383 365.555
R5495 VSS.t1850 VSS.n1382 365.555
R5496 VSS.t1905 VSS.n1381 365.555
R5497 VSS.t1608 VSS.n1095 365.555
R5498 VSS.n1096 VSS.t1835 365.555
R5499 VSS.t1548 VSS.n1101 365.555
R5500 VSS.n1102 VSS.t60 365.555
R5501 VSS.t179 VSS.n2296 365.555
R5502 VSS.n2297 VSS.t623 365.555
R5503 VSS.n2300 VSS.t2084 365.555
R5504 VSS.t1102 VSS.n2304 365.555
R5505 VSS.n2058 VSS.t86 365.555
R5506 VSS.n2057 VSS.t839 365.555
R5507 VSS.t844 VSS.n2050 365.555
R5508 VSS.n2051 VSS.t860 365.555
R5509 VSS.t814 VSS.n2390 365.555
R5510 VSS.n2391 VSS.t1455 365.555
R5511 VSS.n2394 VSS.t1742 365.555
R5512 VSS.t1087 VSS.n2399 365.555
R5513 VSS.n2008 VSS.t1112 365.555
R5514 VSS.n2010 VSS.t1861 365.555
R5515 VSS.n2012 VSS.t1426 365.555
R5516 VSS.n2015 VSS.t1429 365.555
R5517 VSS.n2070 VSS.t1068 365.555
R5518 VSS.n2074 VSS.t1449 365.555
R5519 VSS.n2075 VSS.t1591 365.555
R5520 VSS.n2079 VSS.t1594 365.555
R5521 VSS.t1099 VSS.n2098 365.555
R5522 VSS.t774 VSS.n2097 365.555
R5523 VSS.t1538 VSS.n2096 365.555
R5524 VSS.t185 VSS.n2095 365.555
R5525 VSS.t777 VSS.n2143 365.555
R5526 VSS.t780 VSS.n2142 365.555
R5527 VSS.t321 VSS.n2141 365.555
R5528 VSS.t332 VSS.n2140 365.555
R5529 VSS.n1660 VSS.t833 365.555
R5530 VSS.n1659 VSS.t666 365.555
R5531 VSS.n1658 VSS.t413 365.555
R5532 VSS.n1657 VSS.t1007 365.555
R5533 VSS.n1653 VSS.t619 365.555
R5534 VSS.n1652 VSS.t1997 365.555
R5535 VSS.n1651 VSS.t641 365.555
R5536 VSS.n1650 VSS.t1246 365.555
R5537 VSS.t1351 VSS.n2632 365.555
R5538 VSS.n2633 VSS.t2162 365.555
R5539 VSS.t148 VSS.n2638 365.555
R5540 VSS.n2639 VSS.t1011 365.555
R5541 VSS.t481 VSS.n881 365.555
R5542 VSS.n882 VSS.t478 365.555
R5543 VSS.t967 VSS.n887 365.555
R5544 VSS.n888 VSS.t1374 365.555
R5545 VSS.t993 VSS.n1826 365.555
R5546 VSS.t572 VSS.n1825 365.555
R5547 VSS.n1511 VSS.t1288 365.555
R5548 VSS.n1819 VSS.t363 365.555
R5549 VSS.t504 VSS.n1815 365.555
R5550 VSS.t1485 VSS.n1814 365.555
R5551 VSS.t1489 VSS.n1813 365.555
R5552 VSS.t1913 VSS.n1812 365.555
R5553 VSS.t633 VSS.n921 365.555
R5554 VSS.n922 VSS.t158 365.555
R5555 VSS.n925 VSS.t1569 365.555
R5556 VSS.t285 VSS.n930 365.555
R5557 VSS.n944 VSS.t2094 365.555
R5558 VSS.n943 VSS.t1045 365.555
R5559 VSS.n942 VSS.t50 365.555
R5560 VSS.n941 VSS.t748 365.555
R5561 VSS.n428 VSS.t2371 365.555
R5562 VSS.n432 VSS.t2294 365.555
R5563 VSS.n433 VSS.t1270 365.555
R5564 VSS.n437 VSS.t1642 365.555
R5565 VSS.n448 VSS.t854 365.555
R5566 VSS.n449 VSS.t2195 365.555
R5567 VSS.n452 VSS.t1793 365.555
R5568 VSS.n456 VSS.t1563 365.555
R5569 VSS.n462 VSS.t2380 365.555
R5570 VSS.n467 VSS.t935 365.555
R5571 VSS.n471 VSS.t729 365.555
R5572 VSS.t2356 VSS.n491 365.555
R5573 VSS.t1599 VSS.n490 365.555
R5574 VSS.t1813 VSS.n489 365.555
R5575 VSS.t1817 VSS.n488 365.555
R5576 VSS.n2511 VSS.t441 364.274
R5577 VSS.n2578 VSS.t694 364.274
R5578 VSS.n1911 VSS.t2238 364.274
R5579 VSS.n1528 VSS.t2491 364.274
R5580 VSS.t692 VSS.n324 363.014
R5581 VSS.t1000 VSS.t2157 357.092
R5582 VSS.t1944 VSS.n918 354.747
R5583 VSS.t2543 VSS.t2028 351.351
R5584 VSS.t2512 VSS.t1076 350.877
R5585 VSS.t1165 VSS.t2339 350.877
R5586 VSS.t2036 VSS.t1792 350.877
R5587 VSS.t2138 VSS.t2026 350.877
R5588 VSS.t2078 VSS.t1856 350.404
R5589 VSS.t1123 VSS.t2374 350.404
R5590 VSS.t1982 VSS.t1171 350.404
R5591 VSS.n1131 VSS.n1130 349.661
R5592 VSS.n1187 VSS.n1186 349.661
R5593 VSS.n1160 VSS.n1159 349.661
R5594 VSS.n1169 VSS.n1139 349.661
R5595 VSS.t122 VSS.n2966 348.531
R5596 VSS.n1444 VSS.n1443 347.502
R5597 VSS.n317 VSS.n316 347.168
R5598 VSS.n1152 VSS.n1151 345.981
R5599 VSS.n1723 VSS.n1722 345.394
R5600 VSS.n505 VSS.n504 345.394
R5601 VSS.t2146 VSS.t1092 343.717
R5602 VSS.t2415 VSS.t579 343.717
R5603 VSS.t1094 VSS.t1602 343.717
R5604 VSS.t1776 VSS.t2388 343.717
R5605 VSS.t2323 VSS.t1110 343.717
R5606 VSS.t2400 VSS.t1142 343.717
R5607 VSS.n1466 VSS.t1938 342.106
R5608 VSS.n1217 VSS.n1216 338.957
R5609 VSS.t998 VSS.t0 337.038
R5610 VSS.t125 VSS.t141 337.038
R5611 VSS.t1665 VSS.t985 335.264
R5612 VSS.t143 VSS.t1509 335.264
R5613 VSS.t1115 VSS.t2 331.341
R5614 VSS.t1554 VSS.n2521 331.211
R5615 VSS.n2522 VSS.t1296 331.211
R5616 VSS.t1584 VSS.n2526 331.211
R5617 VSS.n2527 VSS.t1480 331.211
R5618 VSS.n2541 VSS.t1053 331.211
R5619 VSS.n2540 VSS.t176 331.211
R5620 VSS.t961 VSS.n2533 331.211
R5621 VSS.n2534 VSS.t1471 331.211
R5622 VSS.t411 VSS.t577 330.394
R5623 VSS.t1507 VSS.t1726 330.394
R5624 VSS.t450 VSS.t2302 329.37
R5625 VSS.t314 VSS.t234 329.37
R5626 VSS.t399 VSS.t409 329.029
R5627 VSS.t1576 VSS.t391 329.029
R5628 VSS.t1183 VSS.t81 327.675
R5629 VSS.t758 VSS.t595 327.675
R5630 VSS.t497 VSS.t52 327.675
R5631 VSS.t828 VSS.t668 326.19
R5632 VSS.t398 VSS.t1894 326.19
R5633 VSS.n685 VSS.t1349 319.466
R5634 VSS.t1647 VSS.n3142 313.253
R5635 VSS.t2527 VSS.t1583 311.825
R5636 VSS.t1249 VSS.t853 311.825
R5637 VSS.n440 VSS.t2099 311.404
R5638 VSS.n3238 VSS.t1210 311.377
R5639 VSS.n3246 VSS.t1206 311.377
R5640 VSS.n3254 VSS.t1208 311.377
R5641 VSS.t2035 VSS.t1057 310.634
R5642 VSS.t1184 VSS.t2312 310.634
R5643 VSS.t2130 VSS.n2969 306.305
R5644 VSS.t2032 VSS.n347 306.084
R5645 VSS.t1185 VSS.n1847 305.685
R5646 VSS.n3013 VSS.t2515 300.704
R5647 VSS.n1144 VSS.t1355 298.279
R5648 VSS.t1345 VSS.n1197 298.279
R5649 VSS.n507 VSS.n506 297.363
R5650 VSS.n1725 VSS.n1724 297.363
R5651 VSS.t2099 VSS.n439 296.053
R5652 VSS.t277 VSS.t1199 294.406
R5653 VSS.t356 VSS.t1215 291.519
R5654 VSS.n3274 VSS.n3273 290.997
R5655 VSS.n2625 VSS.n2624 287.072
R5656 VSS.n1700 VSS.t1497 281.091
R5657 VSS.n3488 VSS.t2297 281.091
R5658 VSS.n221 VSS.n218 280.072
R5659 VSS.n519 VSS.n518 278.426
R5660 VSS.n1835 VSS.n1493 275.082
R5661 VSS.n1860 VSS.n1859 273.747
R5662 VSS.n3334 VSS.n3333 270.834
R5663 VSS.n3316 VSS.n3315 270.834
R5664 VSS.n1899 VSS.n1898 270.834
R5665 VSS.n2827 VSS.n2826 269.966
R5666 VSS.n856 VSS.t2363 269.688
R5667 VSS.n614 VSS.t1194 269.688
R5668 VSS.t1656 VSS.t1187 265.683
R5669 VSS.n3441 VSS.n33 265.515
R5670 VSS.n2699 VSS.n773 263.781
R5671 VSS.t283 VSS.t288 263.497
R5672 VSS.n871 VSS.t555 255.748
R5673 VSS.n601 VSS.t1977 255.748
R5674 VSS.n3451 VSS.n3450 253.648
R5675 VSS.n1326 VSS.t2403 253.143
R5676 VSS.n3334 VSS.n3318 251.548
R5677 VSS.n3316 VSS.n3300 251.548
R5678 VSS.n1899 VSS.n1233 251.548
R5679 VSS.n248 VSS.n247 251.368
R5680 VSS.n525 VSS.n524 249.748
R5681 VSS.n2591 VSS.n2590 249.748
R5682 VSS.n140 VSS.t2497 247.227
R5683 VSS.n139 VSS.t2068 247.227
R5684 VSS.n135 VSS.t48 247.227
R5685 VSS.n3352 VSS.t757 247.227
R5686 VSS.t2479 VSS.n3359 247.227
R5687 VSS.n3360 VSS.t2069 247.227
R5688 VSS.n3363 VSS.t56 247.227
R5689 VSS.t1078 VSS.n3367 247.227
R5690 VSS.t1240 VSS.n3369 247.227
R5691 VSS.n3371 VSS.t2079 247.227
R5692 VSS.n3373 VSS.t393 247.227
R5693 VSS.n3392 VSS.t1182 247.227
R5694 VSS.t1239 VSS.n3399 247.227
R5695 VSS.n3400 VSS.t2037 247.227
R5696 VSS.t652 VSS.n3404 247.227
R5697 VSS.n3406 VSS.t2386 247.227
R5698 VSS.n2951 VSS.n2950 247.184
R5699 VSS.n2782 VSS.n2781 242.537
R5700 VSS.t1459 VSS.t132 239.969
R5701 VSS.t2270 VSS.n1762 239.774
R5702 VSS.n2703 VSS.n2702 238.584
R5703 VSS.n3471 VSS.n3470 237.565
R5704 VSS.n2964 VSS.n324 237.444
R5705 VSS.t1779 VSS.n1129 235.561
R5706 VSS.t575 VSS.n1131 235.561
R5707 VSS.n1188 VSS.t2290 235.561
R5708 VSS.n1186 VSS.t1343 235.561
R5709 VSS.n1134 VSS.t2288 235.561
R5710 VSS.t1975 VSS.n1150 235.561
R5711 VSS.n1152 VSS.t24 235.561
R5712 VSS.t2180 VSS.n1158 235.561
R5713 VSS.n1160 VSS.t621 235.561
R5714 VSS.n1165 VSS.t751 235.561
R5715 VSS.t1274 VSS.n1169 235.561
R5716 VSS.n1179 VSS.t2378 235.561
R5717 VSS.n1322 VSS.n1117 234.184
R5718 VSS.t1740 VSS.t260 234.03
R5719 VSS.t2088 VSS.t42 234.03
R5720 VSS.t906 VSS.t1464 234.03
R5721 VSS.n1363 VSS.t1081 231.852
R5722 VSS.n2123 VSS.t492 231.852
R5723 VSS.n1589 VSS.t1322 231.852
R5724 VSS.n3272 VSS.n3271 230.413
R5725 VSS.n792 VSS.t2190 228.907
R5726 VSS.n798 VSS.t397 228.907
R5727 VSS.n797 VSS.t1766 228.907
R5728 VSS.n802 VSS.t2030 228.907
R5729 VSS.n807 VSS.t2472 228.907
R5730 VSS.t1892 VSS.n1571 228.571
R5731 VSS.n1566 VSS.t832 228.571
R5732 VSS.n783 VSS.t2080 228.571
R5733 VSS.n1629 VSS.t875 228.571
R5734 VSS.t552 VSS.n810 228.571
R5735 VSS.n815 VSS.t545 228.571
R5736 VSS.n811 VSS.t1546 228.571
R5737 VSS.n2642 VSS.t2045 228.571
R5738 VSS.n813 VSS.t2081 228.571
R5739 VSS.n2645 VSS.t543 228.571
R5740 VSS.t2216 VSS.t1560 225.695
R5741 VSS.t2024 VSS.t1425 225.695
R5742 VSS.t1227 VSS.t2206 225.695
R5743 VSS.t2059 VSS.t1590 225.695
R5744 VSS.t491 VSS.t1229 225.695
R5745 VSS.t2042 VSS.t1541 225.695
R5746 VSS.t1824 VSS.t2211 225.695
R5747 VSS.t2082 VSS.t324 225.695
R5748 VSS.t62 VSS.t2426 223.987
R5749 VSS.t1841 VSS.t2168 223.987
R5750 VSS.n968 VSS.t2159 222.76
R5751 VSS.n1222 VSS.n1203 220
R5752 VSS.n1557 VSS.t2105 217.304
R5753 VSS.t1936 VSS.n1559 217.304
R5754 VSS.n1564 VSS.t2075 217.304
R5755 VSS.n1675 VSS.t1328 217.304
R5756 VSS.n2412 VSS.t277 216.475
R5757 VSS.n3261 VSS.t356 216.475
R5758 VSS.t2350 VSS.t329 214.912
R5759 VSS.t55 VSS.t1075 214.912
R5760 VSS.t1082 VSS.t163 211.208
R5761 VSS.t488 VSS.t1653 211.208
R5762 VSS.t868 VSS.t1636 211.208
R5763 VSS.t1581 VSS.n337 210.811
R5764 VSS.n750 VSS.t1369 210.811
R5765 VSS.t2028 VSS.n749 210.811
R5766 VSS.n748 VSS.t2527 210.811
R5767 VSS.n343 VSS.t1249 210.811
R5768 VSS.n348 VSS.t2032 210.811
R5769 VSS.t1641 VSS.n351 210.526
R5770 VSS.n352 VSS.t2334 210.526
R5771 VSS.t852 VSS.n354 210.526
R5772 VSS.n355 VSS.t1397 210.526
R5773 VSS.t2065 VSS.n358 210.526
R5774 VSS.n359 VSS.t2512 210.526
R5775 VSS.n361 VSS.t1165 210.526
R5776 VSS.n362 VSS.t2036 210.526
R5777 VSS.t329 VSS.n365 210.526
R5778 VSS.n366 VSS.t2350 210.526
R5779 VSS.t1075 VSS.n368 210.526
R5780 VSS.n369 VSS.t55 210.526
R5781 VSS.t2026 VSS.n371 210.526
R5782 VSS.n373 VSS.t1118 210.526
R5783 VSS.n374 VSS.t1250 210.526
R5784 VSS.t2052 VSS.n376 210.526
R5785 VSS.n495 VSS.t2078 210.244
R5786 VSS.n594 VSS.t1123 210.244
R5787 VSS.t1171 VSS.n593 210.244
R5788 VSS.n3238 VSS.t1203 207.585
R5789 VSS.n3246 VSS.t783 207.585
R5790 VSS.n3254 VSS.t358 207.585
R5791 VSS.n1664 VSS.n1587 206.661
R5792 VSS.n2625 VSS.t2305 202.679
R5793 VSS.n3026 VSS.t2421 202.078
R5794 VSS.n3441 VSS.n34 200.053
R5795 VSS.t1255 VSS.t2062 198.954
R5796 VSS.n1144 VSS.t1536 198.853
R5797 VSS.n1197 VSS.t795 198.853
R5798 VSS.n2254 VSS.t911 196.276
R5799 VSS.n295 VSS.t998 196.032
R5800 VSS.n3114 VSS.t125 196.032
R5801 VSS.t311 VSS.t631 195.589
R5802 VSS.t2249 VSS.t154 195.589
R5803 VSS.t1618 VSS.t319 195.589
R5804 VSS.t1521 VSS.t145 195.589
R5805 VSS.n1408 VSS.n1407 195.244
R5806 VSS.n2168 VSS.n2167 195.244
R5807 VSS.n1620 VSS.n1588 195.244
R5808 VSS.n292 VSS.t1665 195
R5809 VSS.n3106 VSS.t143 195
R5810 VSS.n2987 VSS.n18 194.542
R5811 VSS.t965 VSS.n856 192.633
R5812 VSS.n614 VSS.t971 192.633
R5813 VSS.t206 VSS.t417 192.316
R5814 VSS.n3085 VSS.t411 192.168
R5815 VSS.n3090 VSS.t1507 192.168
R5816 VSS.n303 VSS.t450 191.572
R5817 VSS.n3098 VSS.t314 191.572
R5818 VSS.n858 VSS.t399 191.375
R5819 VSS.n620 VSS.t1576 191.375
R5820 VSS.n3332 VSS.t1183 190.587
R5821 VSS.n3314 VSS.t758 190.587
R5822 VSS.n1897 VSS.t497 190.587
R5823 VSS.t2269 VSS.t2514 190.406
R5824 VSS.n1907 VSS.t494 190.095
R5825 VSS.n1863 VSS.t2317 186.715
R5826 VSS.n11 VSS.t1582 186.381
R5827 VSS.t1801 VSS.n1718 186.381
R5828 VSS.n1851 VSS.t1562 186.381
R5829 VSS.n1854 VSS.t2035 186.381
R5830 VSS.n1858 VSS.t2312 186.381
R5831 VSS.t2050 VSS.t1610 186.314
R5832 VSS.t2156 VSS.t440 186.314
R5833 VSS.t1346 VSS.t2377 183.456
R5834 VSS.t244 VSS.n667 180.292
R5835 VSS.n1850 VSS.t1185 180.036
R5836 VSS.n10 VSS.t1254 176.673
R5837 VSS.t2481 VSS.n1719 176.673
R5838 VSS.n3441 VSS.t1001 176.633
R5839 VSS.t1674 VSS.t2033 176.45
R5840 VSS.t2187 VSS.t1327 176.45
R5841 VSS.t2432 VSS.t242 175.202
R5842 VSS.n2978 VSS.n2977 174.951
R5843 VSS.t503 VSS.t2237 174.85
R5844 VSS.t2072 VSS.t1291 174.85
R5845 VSS.n3334 VSS.t721 174.407
R5846 VSS.n3316 VSS.t1079 174.407
R5847 VSS.n1899 VSS.t8 174.407
R5848 VSS.t1888 VSS.n779 173.81
R5849 VSS.t2046 VSS.t230 173.681
R5850 VSS.t2455 VSS.t1833 173.681
R5851 VSS.t2070 VSS.t434 173.507
R5852 VSS.t884 VSS.t1034 173.507
R5853 VSS.n3269 VSS.n222 173.179
R5854 VSS.n3269 VSS.n3226 173.179
R5855 VSS.n3212 VSS.n234 171.989
R5856 VSS.t650 VSS.n18 171.655
R5857 VSS.n962 VSS.t2145 171.576
R5858 VSS.n2959 VSS.t1042 170.512
R5859 VSS.t2023 VSS.t196 169.216
R5860 VSS.t2219 VSS.t2236 167.472
R5861 VSS.t2058 VSS.t1488 167.472
R5862 VSS.t1326 VSS.n2623 166.667
R5863 VSS.t1985 VSS.t2551 166.059
R5864 VSS.t2114 VSS.n1090 165.642
R5865 VSS.t2459 VSS.n1248 165.642
R5866 VSS.t211 VSS.n140 164.819
R5867 VSS.t958 VSS.n139 164.819
R5868 VSS.n135 VSS.t484 164.819
R5869 VSS.n3352 VSS.t1303 164.819
R5870 VSS.n3359 VSS.t225 164.819
R5871 VSS.n3360 VSS.t590 164.819
R5872 VSS.n3363 VSS.t1439 164.819
R5873 VSS.n3367 VSS.t587 164.819
R5874 VSS.n3369 VSS.t208 164.819
R5875 VSS.n3371 VSS.t1864 164.819
R5876 VSS.n3373 VSS.t342 164.819
R5877 VSS.n3392 VSS.t345 164.819
R5878 VSS.n3399 VSS.t220 164.819
R5879 VSS.n3400 VSS.t614 164.819
R5880 VSS.n3404 VSS.t1310 164.819
R5881 VSS.n3406 VSS.t1736 164.819
R5882 VSS.n1573 VSS.n1572 164.286
R5883 VSS.t1232 VSS.t2055 164.245
R5884 VSS.n874 VSS.t407 163.793
R5885 VSS.n639 VSS.t2337 163.793
R5886 VSS.n1325 VSS.n1117 162.359
R5887 VSS.n2597 VSS.t78 161.192
R5888 VSS.t2060 VSS.t157 160.792
R5889 VSS.t697 VSS.t1944 160.792
R5890 VSS.n380 VSS.n379 159.873
R5891 VSS.n383 VSS.n382 159.873
R5892 VSS.n393 VSS.t2138 157.895
R5893 VSS.t1006 VSS.t126 157.72
R5894 VSS.t2053 VSS.t1923 157.72
R5895 VSS.n658 VSS.t1346 154.988
R5896 VSS.n3081 VSS.n3080 154.197
R5897 VSS.n793 VSS.t1634 152.606
R5898 VSS.t340 VSS.n792 152.606
R5899 VSS.n798 VSS.t1994 152.606
R5900 VSS.n797 VSS.t1671 152.606
R5901 VSS.n803 VSS.t977 152.606
R5902 VSS.t765 VSS.n802 152.606
R5903 VSS.n1641 VSS.t1017 152.606
R5904 VSS.t2305 VSS.n807 152.606
R5905 VSS.t1783 VSS.n779 152.381
R5906 VSS.n780 VSS.t1724 152.381
R5907 VSS.t1361 VSS.n782 152.381
R5908 VSS.n789 VSS.t1411 152.381
R5909 VSS.n820 VSS.t136 152.381
R5910 VSS.t2292 VSS.n810 152.381
R5911 VSS.n815 VSS.t1825 152.381
R5912 VSS.n811 VSS.t835 152.381
R5913 VSS.n2642 VSS.t375 152.381
R5914 VSS.t570 VSS.n813 152.381
R5915 VSS.n2645 VSS.t1009 152.381
R5916 VSS.t1616 VSS.n1427 151.915
R5917 VSS.t843 VSS.t2074 151.915
R5918 VSS.t2025 VSS.t1030 151.915
R5919 VSS.t883 VSS.t2462 151.915
R5920 VSS.t308 VSS.t496 151.915
R5921 VSS.t2051 VSS.t1798 151.915
R5922 VSS.t2043 VSS.t463 151.915
R5923 VSS.t2520 VSS.t2458 151.915
R5924 VSS.n675 VSS.t1981 151.826
R5925 VSS.t862 VSS.n1980 150.845
R5926 VSS.t1597 VSS.n1981 150.845
R5927 VSS.n1276 VSS.t458 150.845
R5928 VSS.n1275 VSS.t866 150.845
R5929 VSS.n2421 VSS.t236 150.845
R5930 VSS.t384 VSS.n2426 150.845
R5931 VSS.n1409 VSS.t1605 150.845
R5932 VSS.n1415 VSS.t2132 150.845
R5933 VSS.n2169 VSS.t604 150.845
R5934 VSS.n2175 VSS.t607 150.845
R5935 VSS.t1770 VSS.n1602 150.845
R5936 VSS.n1603 VSS.t1359 150.845
R5937 VSS.n3277 VSS.n3276 147.727
R5938 VSS.t452 VSS.t1173 143.173
R5939 VSS.n1664 VSS.n1662 142.794
R5940 VSS.n1592 VSS.t826 140.889
R5941 VSS.n1560 VSS.t2310 140.889
R5942 VSS.t1684 VSS.n1674 140.889
R5943 VSS.n1576 VSS.t1680 140.889
R5944 VSS.t727 VSS.n337 140.542
R5945 VSS.n750 VSS.t1378 140.542
R5946 VSS.n749 VSS.t62 140.542
R5947 VSS.t2426 VSS.n748 140.542
R5948 VSS.t2168 VSS.n343 140.542
R5949 VSS.n348 VSS.t1841 140.542
R5950 VSS.n351 VSS.t1927 140.351
R5951 VSS.n352 VSS.t1398 140.351
R5952 VSS.n354 VSS.t1931 140.351
R5953 VSS.t2102 VSS.n355 140.351
R5954 VSS.n365 VSS.t1147 140.351
R5955 VSS.n366 VSS.t1884 140.351
R5956 VSS.n368 VSS.t127 140.351
R5957 VSS.n369 VSS.t1280 140.351
R5958 VSS.t2136 VSS.n371 140.351
R5959 VSS.n373 VSS.t2429 140.351
R5960 VSS.t2368 VSS.n374 140.351
R5961 VSS.n376 VSS.t1846 140.351
R5962 VSS.t242 VSS.n495 140.162
R5963 VSS.n594 VSS.t2432 140.162
R5964 VSS.n593 VSS.t183 140.162
R5965 VSS.n597 VSS.t675 140.162
R5966 VSS.t1560 VSS.n2025 135.417
R5967 VSS.n2027 VSS.t2024 135.417
R5968 VSS.t1959 VSS.n2029 135.417
R5969 VSS.t2210 VSS.n2031 135.417
R5970 VSS.t2206 VSS.n2039 135.417
R5971 VSS.n2041 VSS.t2059 135.417
R5972 VSS.t612 VSS.n2043 135.417
R5973 VSS.t1226 VSS.n2045 135.417
R5974 VSS.t1229 VSS.n2102 135.417
R5975 VSS.n2104 VSS.t2042 135.417
R5976 VSS.t1137 VSS.n2106 135.417
R5977 VSS.t487 VSS.n2108 135.417
R5978 VSS.t2211 VSS.n2111 135.417
R5979 VSS.n2113 VSS.t2082 135.417
R5980 VSS.t330 VSS.n2115 135.417
R5981 VSS.n2117 VSS.t1820 135.417
R5982 VSS.n3448 VSS.t2449 135.018
R5983 VSS.t1582 VSS.n10 133.962
R5984 VSS.n1719 VSS.t1801 133.962
R5985 VSS.t2067 VSS.t997 133.862
R5986 VSS.t2029 VSS.t1067 133.862
R5987 VSS.n2494 VSS.t1630 131.371
R5988 VSS.n2251 VSS.t2002 126.761
R5989 VSS.t2473 VSS.n1846 126.603
R5990 VSS.n998 VSS.t2485 125.201
R5991 VSS.t111 VSS.n251 125.201
R5992 VSS.n1000 VSS.t2038 125.201
R5993 VSS.t2063 VSS.n252 125.201
R5994 VSS.n1002 VSS.t335 125.201
R5995 VSS.t1633 VSS.n253 125.201
R5996 VSS.n2498 VSS.t2283 125.201
R5997 VSS.n1863 VSS.t1388 124.477
R5998 VSS.t2342 VSS.n9 124.254
R5999 VSS.t1132 VSS.n11 124.254
R6000 VSS.n1720 VSS.t403 124.254
R6001 VSS.n1718 VSS.t1734 124.254
R6002 VSS.n1851 VSS.t1059 124.254
R6003 VSS.n1854 VSS.t152 124.254
R6004 VSS.t515 VSS.n1858 124.254
R6005 VSS.t545 VSS.t2292 123.811
R6006 VSS.t835 VSS.t2161 123.811
R6007 VSS.t1321 VSS.t570 123.811
R6008 VSS.n1406 VSS.t1082 122.846
R6009 VSS.n2166 VSS.t488 122.846
R6010 VSS.n1618 VSS.t868 122.846
R6011 VSS.n686 VSS.t1639 120.883
R6012 VSS.t296 VSS.n1850 120.023
R6013 VSS.n1308 VSS.n1307 119.948
R6014 VSS.n2463 VSS.n2462 119.948
R6015 VSS.t1622 VSS.n1061 119.948
R6016 VSS.n1048 VSS.n1047 119.948
R6017 VSS.n1442 VSS.n1353 119.948
R6018 VSS.n2292 VSS.n2291 119.948
R6019 VSS.n2305 VSS.n1084 119.948
R6020 VSS.n2386 VSS.n2385 119.948
R6021 VSS.n1656 VSS.n1655 119.948
R6022 VSS.n946 VSS.n932 119.948
R6023 VSS.n3422 VSS.t1063 118.447
R6024 VSS.t2514 VSS.n1753 114.245
R6025 VSS.n1755 VSS.t2066 114.245
R6026 VSS.n3350 VSS.n3349 114.236
R6027 VSS.n2236 VSS.n2234 114.236
R6028 VSS.n2332 VSS.n1083 114.236
R6029 VSS.n1386 VSS.n1385 114.236
R6030 VSS.n2037 VSS.n2036 114.236
R6031 VSS.n2100 VSS.n2099 114.236
R6032 VSS.n2145 VSS.n2144 114.236
R6033 VSS.n1817 VSS.n1816 114.236
R6034 VSS.n444 VSS.n441 114.236
R6035 VSS.n493 VSS.n492 114.236
R6036 VSS.t1951 VSS.n1759 113.953
R6037 VSS.n1763 VSS.t2270 113.953
R6038 VSS.t109 VSS.t1324 113.144
R6039 VSS.n959 VSS.t446 111.788
R6040 VSS.n960 VSS.t1829 111.788
R6041 VSS.n961 VSS.t2050 111.788
R6042 VSS.n964 VSS.t2156 111.788
R6043 VSS.t790 VSS.n658 110.707
R6044 VSS.n1058 VSS.n1017 108.103
R6045 VSS.n3390 VSS.n3389 106.921
R6046 VSS.n1906 VSS.n1231 106.921
R6047 VSS.n2967 VSS.t122 106.558
R6048 VSS.n2878 VSS.n2877 105.492
R6049 VSS.t1187 VSS.t2490 105.222
R6050 VSS.t2054 VSS.t656 105.222
R6051 VSS.t2299 VSS.t1023 105.201
R6052 VSS.n1775 VSS.t2072 104.909
R6053 VSS.t698 VSS.t283 104.356
R6054 VSS.n1282 VSS.t1830 104.209
R6055 VSS.n1283 VSS.t98 104.209
R6056 VSS.n1287 VSS.t2046 104.209
R6057 VSS.n1288 VSS.t2455 104.209
R6058 VSS.n2783 VSS.n2782 104.126
R6059 VSS.t1035 VSS.n1462 104.105
R6060 VSS.t1283 VSS.n1461 104.105
R6061 VSS.n1245 VSS.t2070 104.105
R6062 VSS.n1246 VSS.t884 104.105
R6063 VSS.n499 VSS.t938 103.785
R6064 VSS.t1639 VSS.n685 103.255
R6065 VSS.n246 VSS.t298 101.529
R6066 VSS.n668 VSS.t244 101.218
R6067 VSS.n675 VSS.t2335 101.218
R6068 VSS.t1118 VSS.t2354 100.877
R6069 VSS.t1250 VSS.t2359 100.877
R6070 VSS.n1778 VSS.t361 100.484
R6071 VSS.t507 VSS.n1782 100.484
R6072 VSS.t2236 VSS.n1785 100.484
R6073 VSS.n1787 VSS.t2058 100.484
R6074 VSS.n1789 VSS.t350 100.484
R6075 VSS.n2969 VSS.t382 100.43
R6076 VSS.n311 VSS.n310 100.334
R6077 VSS.t1134 VSS.n503 99.0148
R6078 VSS.t1733 VSS.n1721 99.0148
R6079 VSS.n499 VSS.t2052 99.0121
R6080 VSS.n2971 VSS.t2130 98.5476
R6081 VSS.n2417 VSS.t1809 97.7946
R6082 VSS.n1571 VSS.t400 97.6195
R6083 VSS.n1566 VSS.t1782 97.6195
R6084 VSS.n783 VSS.t2044 97.6195
R6085 VSS.n1629 VSS.t2496 97.6195
R6086 VSS.n915 VSS.t1940 96.4755
R6087 VSS.n916 VSS.t705 96.4755
R6088 VSS.n917 VSS.t2060 96.4755
R6089 VSS.n948 VSS.t697 96.4755
R6090 VSS.n2925 VSS.t287 96.4755
R6091 VSS.n2926 VSS.t2092 96.4755
R6092 VSS.n245 VSS.t1337 95.7942
R6093 VSS.n2974 VSS.t1006 94.632
R6094 VSS.t1005 VSS.n3469 94.632
R6095 VSS.t456 VSS.n3468 94.632
R6096 VSS.n3023 VSS.t2053 94.632
R6097 VSS.n3029 VSS.t449 94.632
R6098 VSS.t913 VSS.t2252 94.0088
R6099 VSS.t1579 VSS.t1518 94.0088
R6100 VSS.t721 VSS.t316 93.9117
R6101 VSS.t1079 VSS.t170 93.9117
R6102 VSS.t8 VSS.t1744 93.9117
R6103 VSS.n3033 VSS.n3032 92.9707
R6104 VSS.n1328 VSS.t885 91.1486
R6105 VSS.n1332 VSS.t311 91.1486
R6106 VSS.n1333 VSS.t2465 91.1486
R6107 VSS.n1334 VSS.t2249 91.1486
R6108 VSS.n1337 VSS.t2025 91.1486
R6109 VSS.n1446 VSS.t2462 91.1486
R6110 VSS.t496 VSS.n1445 91.1486
R6111 VSS.t2456 VSS.n1122 91.1486
R6112 VSS.n1939 VSS.t1618 91.1486
R6113 VSS.n1940 VSS.t1764 91.1486
R6114 VSS.n1425 VSS.t2051 91.1486
R6115 VSS.n1426 VSS.t2043 91.1486
R6116 VSS.n1428 VSS.t2520 91.1486
R6117 VSS.n3036 VSS.t2076 90.4091
R6118 VSS.n2025 VSS.t1089 90.2783
R6119 VSS.n2027 VSS.t1442 90.2783
R6120 VSS.n2029 VSS.t636 90.2783
R6121 VSS.n2031 VSS.t628 90.2783
R6122 VSS.n2039 VSS.t1107 90.2783
R6123 VSS.n2041 VSS.t1702 90.2783
R6124 VSS.n2043 VSS.t1384 90.2783
R6125 VSS.n2045 VSS.t1356 90.2783
R6126 VSS.n2102 VSS.t1104 90.2783
R6127 VSS.n2104 VSS.t1422 90.2783
R6128 VSS.n2106 VSS.t1542 90.2783
R6129 VSS.n2108 VSS.t1139 90.2783
R6130 VSS.t1096 VSS.n2111 90.2783
R6131 VSS.n2113 VSS.t887 90.2783
R6132 VSS.n2115 VSS.t2329 90.2783
R6133 VSS.n2117 VSS.t2096 90.2783
R6134 VSS.t1980 VSS.t890 89.7916
R6135 VSS.t1525 VSS.t282 89.7916
R6136 VSS.t1524 VSS.t1404 89.7916
R6137 VSS.t1853 VSS.t2355 89.7916
R6138 VSS.n3195 VSS.t2023 89.278
R6139 VSS.t1354 VSS.n1744 87.9347
R6140 VSS.t1667 VSS.t2423 87.7198
R6141 VSS.t2125 VSS.t1515 87.7198
R6142 VSS.n3143 VSS.t1647 87.4199
R6143 VSS.n3430 VSS.t2017 87.4199
R6144 VSS.n3444 VSS.t2385 87.4199
R6145 VSS.n503 VSS.n9 87.3661
R6146 VSS.n1721 VSS.n1720 87.3661
R6147 VSS.n1171 VSS.t138 87.1833
R6148 VSS.n3223 VSS.t2285 86.8686
R6149 VSS.t1004 VSS.t1690 84.6881
R6150 VSS.n998 VSS.t1459 83.4676
R6151 VSS.n253 VSS.t214 83.4676
R6152 VSS.n2498 VSS.t955 83.4676
R6153 VSS.n3136 VSS.t1701 81.0184
R6154 VSS.n2740 VSS.n2739 80.5908
R6155 VSS.n3222 VSS.n3221 79.6296
R6156 VSS.n511 VSS.t2047 78.9188
R6157 VSS.n3223 VSS.n223 78.6854
R6158 VSS.t2485 VSS.t111 78.2509
R6159 VSS.t2284 VSS.t1420 78.2509
R6160 VSS.t1418 VSS.t823 78.2509
R6161 VSS.t2038 VSS.t2063 78.2509
R6162 VSS.t1550 VSS.t713 78.2509
R6163 VSS.t2263 VSS.t952 78.2509
R6164 VSS.t335 VSS.t1633 78.2509
R6165 VSS.n2601 VSS.n2600 77.2216
R6166 VSS.n634 VSS.n633 77.2216
R6167 VSS.t2237 VSS.n1774 76.4968
R6168 VSS.t375 VSS.t480 76.191
R6169 VSS.t1009 VSS.t557 76.191
R6170 VSS.n1753 VSS.t508 76.1631
R6171 VSS.n1755 VSS.t939 76.1631
R6172 VSS.n1746 VSS.t1024 76.0517
R6173 VSS.n1759 VSS.t1897 75.9684
R6174 VSS.n1763 VSS.t1285 75.9684
R6175 VSS.t1970 VSS.n49 75.5819
R6176 VSS.n3144 VSS.t1172 75.5819
R6177 VSS.n3428 VSS.t1694 75.5819
R6178 VSS.t905 VSS.n3427 75.5819
R6179 VSS.n1058 VSS.n1057 75.1074
R6180 VSS.n310 VSS.t12 74.768
R6181 VSS.t428 VSS.n959 74.5258
R6182 VSS.n960 VSS.t1614 74.5258
R6183 VSS.t760 VSS.n961 74.5258
R6184 VSS.t5 VSS.n3079 72.8445
R6185 VSS.n2259 VSS.t2410 72.6008
R6186 VSS.n2258 VSS.t1717 72.6008
R6187 VSS.n2267 VSS.t1144 72.6008
R6188 VSS.n2268 VSS.t1445 72.6008
R6189 VSS.n2263 VSS.t1265 72.6008
R6190 VSS.t1092 VSS.n2272 72.6008
R6191 VSS.n2273 VSS.t2146 72.6008
R6192 VSS.t579 VSS.n1106 72.6008
R6193 VSS.n2277 VSS.t2415 72.6008
R6194 VSS.n1107 VSS.t305 72.6008
R6195 VSS.n2281 VSS.t1760 72.6008
R6196 VSS.n2282 VSS.t105 72.6008
R6197 VSS.n2312 VSS.t2182 72.6008
R6198 VSS.n2311 VSS.t1094 72.6008
R6199 VSS.n2339 VSS.t1602 72.6008
R6200 VSS.n2342 VSS.t1776 72.6008
R6201 VSS.n2347 VSS.t2388 72.6008
R6202 VSS.n2346 VSS.t67 72.6008
R6203 VSS.n2355 VSS.t672 72.6008
R6204 VSS.n2356 VSS.t979 72.6008
R6205 VSS.n2351 VSS.t115 72.6008
R6206 VSS.t1110 VSS.n2360 72.6008
R6207 VSS.n2361 VSS.t2323 72.6008
R6208 VSS.t1142 VSS.n1074 72.6008
R6209 VSS.n2365 VSS.t2400 72.6008
R6210 VSS.n1075 VSS.t787 72.6008
R6211 VSS.n2375 VSS.t26 72.6008
R6212 VSS.n2376 VSS.t846 72.6008
R6213 VSS.n2369 VSS.t16 72.6008
R6214 VSS.n2404 VSS.t1115 72.6008
R6215 VSS.n3042 VSS.n3041 72.5157
R6216 VSS.t2061 VSS.n3124 71.4189
R6217 VSS.n3125 VSS.t2530 71.4189
R6218 VSS.n3130 VSS.t1693 71.4189
R6219 VSS.t2040 VSS.n3129 71.4189
R6220 VSS.t382 VSS.n2967 71.0388
R6221 VSS.n1771 VSS.t529 69.94
R6222 VSS.n1775 VSS.t921 69.94
R6223 VSS.t626 VSS.n1282 69.4728
R6224 VSS.n1283 VSS.t232 69.4728
R6225 VSS.t944 VSS.n1287 69.4728
R6226 VSS.n1288 VSS.t2395 69.4728
R6227 VSS.n1462 VSS.t166 69.4032
R6228 VSS.n1461 VSS.t90 69.4032
R6229 VSS.t1751 VSS.n1245 69.4032
R6230 VSS.t2403 VSS.n1246 69.4032
R6231 VSS.t501 VSS.n1124 69.0271
R6232 VSS.t1811 VSS.n240 68.5066
R6233 VSS.n3195 VSS.t1588 68.4891
R6234 VSS.t1173 VSS.n3035 68.0071
R6235 VSS.n246 VSS.t194 67.6868
R6236 VSS.n1778 VSS.t924 66.9892
R6237 VSS.n1782 VSS.t663 66.9892
R6238 VSS.n1785 VSS.t523 66.9892
R6239 VSS.n1787 VSS.t119 66.9892
R6240 VSS.n1789 VSS.t1512 66.9892
R6241 VSS.t78 VSS.n2596 66.9892
R6242 VSS.t910 VSS.t2000 66.9289
R6243 VSS.t1717 VSS.t1261 66.9289
R6244 VSS.t1144 VSS.t1834 66.9289
R6245 VSS.t2031 VSS.t2041 66.9289
R6246 VSS.t1445 VSS.t598 66.9289
R6247 VSS.t1265 VSS.t1948 66.9289
R6248 VSS.t2111 VSS.t2006 66.9289
R6249 VSS.t1840 VSS.t1151 66.9289
R6250 VSS.t305 VSS.t2273 66.9289
R6251 VSS.t1760 VSS.t625 66.9289
R6252 VSS.t2077 VSS.t2022 66.9289
R6253 VSS.t105 VSS.t928 66.9289
R6254 VSS.t2182 VSS.t2016 66.9289
R6255 VSS.t688 VSS.t1963 66.9289
R6256 VSS.t1775 VSS.t2275 66.9289
R6257 VSS.t67 VSS.t1084 66.9289
R6258 VSS.t672 VSS.t838 66.9289
R6259 VSS.t2064 VSS.t2073 66.9289
R6260 VSS.t979 VSS.t1719 66.9289
R6261 VSS.t115 VSS.t683 66.9289
R6262 VSS.t2113 VSS.t942 66.9289
R6263 VSS.t812 VSS.t2200 66.9289
R6264 VSS.t787 VSS.t1908 66.9289
R6265 VSS.t26 VSS.t1454 66.9289
R6266 VSS.t2057 VSS.t2048 66.9289
R6267 VSS.t846 VSS.t1849 66.9289
R6268 VSS.t16 VSS.t2116 66.9289
R6269 VSS.t2528 VSS.t426 66.9289
R6270 VSS.n2708 VSS.n2707 66.6913
R6271 VSS.n2589 VSS.n2588 66.5534
R6272 VSS.t1062 VSS.n3419 66.4117
R6273 VSS.n2971 VSS.t1567 65.6985
R6274 VSS.t2 VSS.n2403 64.7577
R6275 VSS.t1961 VSS.n915 64.3171
R6276 VSS.n916 VSS.t161 64.3171
R6277 VSS.t1299 VSS.n917 64.3171
R6278 VSS.n948 VSS.t247 64.3171
R6279 VSS.t380 VSS.n2925 64.3171
R6280 VSS.n2926 VSS.t189 64.3171
R6281 VSS.n239 VSS.t470 64.0579
R6282 VSS.t2250 VSS.n245 63.8629
R6283 VSS.n2273 VSS.n1091 63.5258
R6284 VSS.n2340 VSS.n2339 63.5258
R6285 VSS.n2361 VSS.n1071 63.5258
R6286 VSS.t706 VSS.n3033 63.2993
R6287 VSS.t2490 VSS.n1738 63.1328
R6288 VSS.n1739 VSS.t2054 63.1328
R6289 VSS.n2974 VSS.t273 63.0882
R6290 VSS.n3469 VSS.t806 63.0882
R6291 VSS.n3468 VSS.t1924 63.0882
R6292 VSS.n3023 VSS.t1306 63.0882
R6293 VSS.n3029 VSS.t271 63.0882
R6294 VSS.n1463 VSS.n1242 62.8967
R6295 VSS.n2930 VSS.t2047 62.6134
R6296 VSS.n2933 VSS.t698 62.6134
R6297 VSS.n2235 VSS.n1106 62.3914
R6298 VSS.n2342 VSS.n2341 62.3914
R6299 VSS.n1365 VSS.n1074 62.3914
R6300 VSS.n2623 VSS.n820 61.9053
R6301 VSS.t631 VSS.n1328 60.7659
R6302 VSS.t735 VSS.n1332 60.7659
R6303 VSS.t154 VSS.n1333 60.7659
R6304 VSS.n1334 VSS.t1505 60.7659
R6305 VSS.t368 VSS.n1329 60.7659
R6306 VSS.n1337 VSS.t1659 60.7659
R6307 VSS.n1446 VSS.t2393 60.7659
R6308 VSS.n1445 VSS.t519 60.7659
R6309 VSS.t319 VSS.n1122 60.7659
R6310 VSS.t797 VSS.n1939 60.7659
R6311 VSS.n1940 VSS.t1521 60.7659
R6312 VSS.t464 VSS.n1123 60.7659
R6313 VSS.t1886 VSS.n1425 60.7659
R6314 VSS.t821 VSS.n1426 60.7659
R6315 VSS.n1428 VSS.t2405 60.7659
R6316 VSS.n3042 VSS.t549 60.2729
R6317 VSS.n3036 VSS.t191 60.2729
R6318 VSS.n2402 VSS.t1909 59.8291
R6319 VSS.n3124 VSS.t255 59.3612
R6320 VSS.n3125 VSS.t29 59.3612
R6321 VSS.n3130 VSS.t1413 59.3612
R6322 VSS.n3129 VSS.t1469 59.3612
R6323 VSS.n2976 VSS.n311 59.271
R6324 VSS.t112 VSS.t1241 58.5375
R6325 VSS.t146 VSS.t499 58.5375
R6326 VSS.n3140 VSS.t669 58.2801
R6327 VSS.t1648 VSS.n3141 58.2801
R6328 VSS.n3143 VSS.t1740 58.2801
R6329 VSS.n3144 VSS.t2088 58.2801
R6330 VSS.n3428 VSS.t42 58.2801
R6331 VSS.n3430 VSS.t906 58.2801
R6332 VSS.n3444 VSS.t2018 58.2801
R6333 VSS.n3452 VSS.t251 57.2692
R6334 VSS.n1574 VSS.n1573 57.1434
R6335 VSS.n687 VSS.n686 56.6646
R6336 VSS.n2815 VSS.n2814 56.0488
R6337 VSS.t218 VSS.t132 55.8599
R6338 VSS.n3034 VSS.t708 55.5641
R6339 VSS.n1784 VSS.n1783 55.4755
R6340 VSS.t271 VSS.n19 55.2022
R6341 VSS.n1017 VSS.t223 55.1368
R6342 VSS.n439 VSS.t2065 54.8251
R6343 VSS.t400 VSS.t1888 54.7624
R6344 VSS.t1782 VSS.t1573 54.7624
R6345 VSS.t2080 VSS.t828 54.7624
R6346 VSS.t2044 VSS.t1341 54.7624
R6347 VSS.t875 VSS.t398 54.7624
R6348 VSS.t2496 VSS.t1013 54.7624
R6349 VSS.n3142 VSS.t1648 54.6377
R6350 VSS.n544 VSS.n363 54.1355
R6351 VSS.t519 VSS.n1444 54.1197
R6352 VSS.n3136 VSS.t292 54.0124
R6353 VSS.n1443 VSS.t2456 53.1702
R6354 VSS.n500 VSS.n499 52.8093
R6355 VSS.t2423 VSS.n358 52.6321
R6356 VSS.n359 VSS.t1667 52.6321
R6357 VSS.t1515 VSS.n361 52.6321
R6358 VSS.n362 VSS.t2125 52.6321
R6359 VSS.t1812 VSS.n236 52.6004
R6360 VSS.n803 VSS.t1674 52.4583
R6361 VSS.n1641 VSS.t2187 52.4583
R6362 VSS.n2978 VSS.n2966 52.1692
R6363 VSS.n918 VSS.t1299 51.2528
R6364 VSS.n379 VSS.t1980 50.3711
R6365 VSS.t282 VSS.n380 50.3711
R6366 VSS.n382 VSS.t1524 50.3711
R6367 VSS.t2355 VSS.n383 50.3711
R6368 VSS.n2944 VSS.n2943 50.3016
R6369 VSS.t1856 VSS.n494 48.1811
R6370 VSS.t1626 VSS.t1811 47.865
R6371 VSS.t422 VSS.n13 47.8266
R6372 VSS.n3474 VSS.t2351 47.8266
R6373 VSS.t348 VSS.n1710 47.8266
R6374 VSS.n1711 VSS.t2188 47.8266
R6375 VSS.n1542 VSS.t732 47.5615
R6376 VSS.n971 VSS.t424 47.5615
R6377 VSS.t1381 VSS.n410 47.5615
R6378 VSS.t1956 VSS.n671 47.5615
R6379 VSS.t1372 VSS.n2586 47.5615
R6380 VSS.n1925 VSS.t31 47.5615
R6381 VSS.n2235 VSS.t2013 46.5101
R6382 VSS.n2341 VSS.t682 46.5101
R6383 VSS.n1365 VSS.t2120 46.5101
R6384 VSS.t513 VSS.n1124 46.0182
R6385 VSS.t2435 VSS.n1091 45.3757
R6386 VSS.t2274 VSS.n2340 45.3757
R6387 VSS.t1083 VSS.n1071 45.3757
R6388 VSS.t2062 VSS.n588 45.3318
R6389 VSS.t2066 VSS.n1754 45.222
R6390 VSS.n3174 VSS.t1475 44.2747
R6391 VSS.n256 VSS.t792 44.2747
R6392 VSS.n3178 VSS.t1753 44.2747
R6393 VSS.n3179 VSS.t1032 44.2747
R6394 VSS.n3415 VSS.t1757 44.2747
R6395 VSS.n3414 VSS.t206 44.2747
R6396 VSS.n3419 VSS.t417 44.2747
R6397 VSS.t1030 VSS.t368 43.6756
R6398 VSS.t2393 VSS.t308 43.6756
R6399 VSS.t463 VSS.t1886 43.6756
R6400 VSS.t2405 VSS.t1616 43.6756
R6401 VSS.n2731 VSS.n2730 43.2086
R6402 VSS.n3174 VSS.t2255 42.8911
R6403 VSS.t1220 VSS.n256 42.8911
R6404 VSS.t2056 VSS.n3178 42.8911
R6405 VSS.n3179 VSS.t2039 42.8911
R6406 VSS.n3415 VSS.t96 42.8911
R6407 VSS.t1534 VSS.n3414 42.8911
R6408 VSS.n1738 VSS.t526 42.0887
R6409 VSS.n1739 VSS.t1656 42.0887
R6410 VSS.n1743 VSS.t657 42.0887
R6411 VSS.n2259 VSS.t910 41.9726
R6412 VSS.t2000 VSS.n2258 41.9726
R6413 VSS.t2041 VSS.n2267 41.9726
R6414 VSS.n2268 VSS.t2031 41.9726
R6415 VSS.n2263 VSS.t2111 41.9726
R6416 VSS.n2272 VSS.t2006 41.9726
R6417 VSS.n2277 VSS.t1840 41.9726
R6418 VSS.t1151 VSS.n1107 41.9726
R6419 VSS.t2022 VSS.n2281 41.9726
R6420 VSS.n2282 VSS.t2077 41.9726
R6421 VSS.n2312 VSS.t688 41.9726
R6422 VSS.t1963 VSS.n2311 41.9726
R6423 VSS.n2347 VSS.t1775 41.9726
R6424 VSS.t2275 VSS.n2346 41.9726
R6425 VSS.t2073 VSS.n2355 41.9726
R6426 VSS.n2356 VSS.t2064 41.9726
R6427 VSS.n2351 VSS.t2113 41.9726
R6428 VSS.n2360 VSS.t942 41.9726
R6429 VSS.n2365 VSS.t812 41.9726
R6430 VSS.t2200 VSS.n1075 41.9726
R6431 VSS.t2048 VSS.n2375 41.9726
R6432 VSS.n2376 VSS.t2057 41.9726
R6433 VSS.n2369 VSS.t2528 41.9726
R6434 VSS.n2404 VSS.t426 41.9726
R6435 VSS.t288 VSS.n2930 41.7424
R6436 VSS.n2933 VSS.t249 41.7424
R6437 VSS.n3164 VSS.n3163 41.0359
R6438 VSS.n3156 VSS.n3155 41.0359
R6439 VSS.n538 VSS.n509 41.0359
R6440 VSS.n2400 VSS.n1070 41.0359
R6441 VSS.n823 VSS.n822 41.0359
R6442 VSS.n347 VSS.t1273 40.4928
R6443 VSS.t1924 VSS.n3467 40.416
R6444 VSS.n1665 VSS.t689 40.409
R6445 VSS.t2283 VSS.n2497 39.2057
R6446 VSS.n511 VSS.t1044 39.1934
R6447 VSS.n3440 VSS.t268 39.1167
R6448 VSS.n2403 VSS.n2402 37.2714
R6449 VSS.n3020 VSS.n3019 37.1859
R6450 VSS.n2651 VSS.n2650 37.1434
R6451 VSS.n1760 VSS.t1951 36.7974
R6452 VSS.t2465 VSS.t735 36.08
R6453 VSS.t1505 VSS.t843 36.08
R6454 VSS.t1659 VSS.t883 36.08
R6455 VSS.t1764 VSS.t797 36.08
R6456 VSS.t1798 VSS.t464 36.08
R6457 VSS.t2458 VSS.t821 36.08
R6458 VSS.n1861 VSS.t1393 36.0732
R6459 VSS.n3236 VSS.n3232 35.7094
R6460 VSS.n183 VSS.n141 34.5908
R6461 VSS.n3058 VSS.t2418 34.3315
R6462 VSS.n242 VSS.n241 34.2979
R6463 VSS.n1982 VSS.t394 34.2711
R6464 VSS.n1986 VSS.t101 34.2711
R6465 VSS.t864 VSS.n1274 34.2711
R6466 VSS.n1261 VSS.t1040 34.2711
R6467 VSS.n1307 VSS.t2463 34.2711
R6468 VSS.n3349 VSS.t2503 34.2711
R6469 VSS.t1236 VSS.n3383 34.2711
R6470 VSS.t93 VSS.n74 34.2711
R6471 VSS.n2462 VSS.t2260 34.2711
R6472 VSS.t1630 VSS.n2493 34.2711
R6473 VSS.n2427 VSS.t352 34.2711
R6474 VSS.t916 VSS.n2443 34.2711
R6475 VSS.n2434 VSS.t2175 34.2711
R6476 VSS.n1063 VSS.t1622 34.2711
R6477 VSS.t2159 VSS.n967 34.2711
R6478 VSS.t436 VSS.n1048 34.2711
R6479 VSS.n1834 VSS.t2521 34.2711
R6480 VSS.n1322 VSS.t881 34.2711
R6481 VSS.n1353 VSS.t2453 34.2711
R6482 VSS.n2234 VSS.t1155 34.2711
R6483 VSS.n2332 VSS.t2277 34.2711
R6484 VSS.n1385 VSS.t1258 34.2711
R6485 VSS.n2291 VSS.t2109 34.2711
R6486 VSS.n2305 VSS.t686 34.2711
R6487 VSS.n2385 VSS.t2117 34.2711
R6488 VSS.n2036 VSS.t2213 34.2711
R6489 VSS.n2099 VSS.t1221 34.2711
R6490 VSS.n2144 VSS.t2207 34.2711
R6491 VSS.t869 VSS.n1656 34.2711
R6492 VSS.n1645 VSS.t1318 34.2711
R6493 VSS.n1816 VSS.t2233 34.2711
R6494 VSS.n932 VSS.t702 34.2711
R6495 VSS.t2476 VSS.n427 34.2711
R6496 VSS.t2468 VSS.n444 34.2711
R6497 VSS.t1127 VSS.n461 34.2711
R6498 VSS.n492 VSS.t1124 34.2711
R6499 VSS.n974 VSS.t389 34.1511
R6500 VSS.n2575 VSS.t771 34.1511
R6501 VSS.t2229 VSS.n1918 34.1511
R6502 VSS.t802 VSS.n1535 34.1511
R6503 VSS.n3278 VSS.n3277 32.8288
R6504 VSS.n2221 VSS.n2220 32.8288
R6505 VSS.n3169 VSS.n3168 32.7461
R6506 VSS.n2542 VSS.t1480 32.6553
R6507 VSS.n2797 VSS.n2796 31.6277
R6508 VSS.t449 VSS.n3028 31.5443
R6509 VSS.n2596 VSS.n2595 31.4015
R6510 VSS.n2654 VSS.n2653 30.9563
R6511 VSS.n524 VSS.n522 30.0931
R6512 VSS.n2592 VSS.n2591 30.0931
R6513 VSS.n2590 VSS.n2589 30.0931
R6514 VSS.n3019 VSS.n25 29.7488
R6515 VSS.n1774 VSS.n1771 28.4134
R6516 VSS.n2803 VSS.t312 28.0246
R6517 VSS.t223 VSS.n242 27.7857
R6518 VSS.n562 VSS.n377 27.068
R6519 VSS.n1984 VSS.n1090 27.0388
R6520 VSS.n1259 VSS.n1248 27.0388
R6521 VSS.t218 VSS.n248 26.7539
R6522 VSS.n2624 VSS.t1326 25.9531
R6523 VSS.t2055 VSS.n2970 25.6638
R6524 VSS.n2815 VSS.t405 25.6226
R6525 VSS.t689 VSS.t109 25.4001
R6526 VSS.n2951 VSS.t583 25.1766
R6527 VSS.t1042 VSS.n2958 25.1766
R6528 VSS.t810 VSS.n2964 25.1147
R6529 VSS.n2965 VSS.t808 25.1147
R6530 VSS.n2939 VSS.t1983 25.0286
R6531 VSS.n237 VSS.t1812 24.9985
R6532 VSS.t1023 VSS.n3208 24.9985
R6533 VSS.n2593 VSS.n2592 24.7283
R6534 VSS.t268 VSS.t720 24.5878
R6535 VSS.n2811 VSS.t556 24.4215
R6536 VSS.t987 VSS.n687 23.9253
R6537 VSS.n557 VSS.n556 23.5512
R6538 VSS.n840 VSS.n839 23.5512
R6539 VSS.t2255 VSS.t1220 23.5211
R6540 VSS.t792 VSS.t1065 23.5211
R6541 VSS.t1753 VSS.t950 23.5211
R6542 VSS.t2039 VSS.t2056 23.5211
R6543 VSS.t1032 VSS.t1869 23.5211
R6544 VSS.t1757 VSS.t1632 23.5211
R6545 VSS.t96 VSS.t1534 23.5211
R6546 VSS.t2537 VSS.t513 23.0094
R6547 VSS.n522 VSS.n514 22.8611
R6548 VSS.t1166 VSS.n502 22.8476
R6549 VSS.n2620 VSS.t2486 22.8476
R6550 VSS.n1172 VSS.t700 22.8476
R6551 VSS.n1869 VSS.n1868 22.5699
R6552 VSS.n2811 VSS.n2810 22.0195
R6553 VSS.n1407 VSS.n1364 21.6311
R6554 VSS.n2167 VSS.n2147 21.6311
R6555 VSS.n1620 VSS.n1619 21.6311
R6556 VSS.n693 VSS.n692 21.6005
R6557 VSS.n3388 VSS.t1178 20.9066
R6558 VSS.n1905 VSS.t493 20.9066
R6559 VSS.n2808 VSS.n2807 20.8184
R6560 VSS.n692 VSS.n691 20.6105
R6561 VSS.n300 VSS.n299 20.5268
R6562 VSS.n2802 VSS.t896 20.4181
R6563 VSS.t555 VSS.t1802 20.1154
R6564 VSS.t407 VSS.t401 20.1154
R6565 VSS.t1977 VSS.t1578 20.1154
R6566 VSS.t2337 VSS.t2340 20.1154
R6567 VSS.n2803 VSS.n2802 18.8167
R6568 VSS.n3041 VSS.t679 17.8939
R6569 VSS.n1861 VSS.t1390 17.8773
R6570 VSS.t292 VSS.n3133 17.7232
R6571 VSS.t2145 VSS.t255 17.6232
R6572 VSS.t2530 VSS.t2061 17.6232
R6573 VSS.t29 VSS.t1000 17.6232
R6574 VSS.t2157 VSS.t1413 17.6232
R6575 VSS.t1693 VSS.t2040 17.6232
R6576 VSS.t1469 VSS.t1708 17.6232
R6577 VSS.t558 VSS.n909 17.2419
R6578 VSS.n636 VSS.t2245 17.2419
R6579 VSS.n3083 VSS.n306 16.8573
R6580 VSS.n1827 VSS.n1506 16.8399
R6581 VSS.n3333 VSS.n3332 16.7186
R6582 VSS.n3315 VSS.n3314 16.7186
R6583 VSS.n1898 VSS.n1897 16.7186
R6584 VSS.n3208 VSS.t470 16.6658
R6585 VSS.n3465 VSS.n25 16.6063
R6586 VSS.t1844 VSS.n2614 16.5119
R6587 VSS.n610 VSS.t973 16.5119
R6588 VSS.n1575 VSS.n1574 16.3322
R6589 VSS.n1407 VSS.n1363 16.2708
R6590 VSS.n2167 VSS.n2123 16.2708
R6591 VSS.n1620 VSS.n1589 16.2708
R6592 VSS.t885 VSS.n1327 16.1413
R6593 VSS.n1745 VSS.t508 15.4501
R6594 VSS.n964 VSS.n963 15.1384
R6595 VSS.n3209 VSS.t2299 15.1035
R6596 VSS.n1744 VSS.n1743 14.4683
R6597 VSS.n3211 VSS.n235 13.8894
R6598 VSS.n2945 VSS.n2944 13.8389
R6599 VSS.n2950 VSS.n2949 13.7329
R6600 VSS.n1870 VSS.n1869 13.5422
R6601 VSS.n691 VSS.n497 13.2511
R6602 VSS.n899 VSS.n898 13.1576
R6603 VSS.t1178 VSS.t112 13.1415
R6604 VSS.t493 VSS.t146 13.1415
R6605 VSS.n2944 VSS.t84 12.5802
R6606 VSS.n694 VSS.t243 11.9903
R6607 VSS.t2105 VSS.t1806 11.9402
R6608 VSS.t826 VSS.t1292 11.9402
R6609 VSS.t1363 VSS.t1936 11.9402
R6610 VSS.t2310 VSS.t107 11.9402
R6611 VSS.t1935 VSS.t1785 11.9402
R6612 VSS.t2075 VSS.t2049 11.9402
R6613 VSS.t617 VSS.t1684 11.9402
R6614 VSS.t2108 VSS.t1803 11.9402
R6615 VSS.t1328 VSS.t2471 11.9402
R6616 VSS.t1680 VSS.t1015 11.9402
R6617 VSS.t997 VSS.t1970 11.8385
R6618 VSS.t1172 VSS.t2067 11.8385
R6619 VSS.t1694 VSS.t2029 11.8385
R6620 VSS.t1067 VSS.t905 11.8385
R6621 VSS.t692 VSS.n2959 11.6322
R6622 VSS.n2950 VSS.t585 11.4343
R6623 VSS.n574 VSS.n502 11.424
R6624 VSS.n2620 VSS.n2619 11.424
R6625 VSS.n1174 VSS.n1172 11.424
R6626 VSS.n1202 VSS.n1200 11.2384
R6627 VSS.n298 VSS.n297 10.318
R6628 VSS.n233 VSS.t2552 10.2719
R6629 VSS.n660 VSS.t151 10.2623
R6630 VSS.n2806 VSS.t1302 10.2623
R6631 VSS.n2509 VSS.n977 10.1567
R6632 VSS.n3012 VSS.n3009 9.623
R6633 VSS.n667 VSS.t1349 9.48955
R6634 VSS.n659 VSS.t150 9.48955
R6635 VSS VSS.t124 9.43705
R6636 VSS.n558 VSS.n557 9.42079
R6637 VSS.n841 VSS.n840 9.42079
R6638 VSS VSS.t1200 9.40995
R6639 VSS VSS.t1216 9.40995
R6640 VSS.n3475 VSS.t2352 9.40866
R6641 VSS.n1712 VSS.t2189 9.40866
R6642 VSS.n2003 VSS.t431 9.37686
R6643 VSS.n1253 VSS.t461 9.37686
R6644 VSS.n2420 VSS.t2010 9.37686
R6645 VSS.n1413 VSS.n1412 9.37686
R6646 VSS.n2173 VSS.n2172 9.37686
R6647 VSS.n1599 VSS.t1773 9.37686
R6648 VSS.n1867 VSS.t2314 9.3736
R6649 VSS.n1239 VSS.t1747 9.3736
R6650 VSS.n821 VSS.t2483 9.3736
R6651 VSS.n838 VSS.t2495 9.3736
R6652 VSS.n1232 VSS.t500 9.3736
R6653 VSS.n2290 VSS.t2110 9.3736
R6654 VSS.n2306 VSS.t687 9.3736
R6655 VSS.n2384 VSS.t2118 9.3736
R6656 VSS.n1323 VSS.t882 9.3736
R6657 VSS.n1306 VSS.t2464 9.3736
R6658 VSS.n1352 VSS.t2454 9.3736
R6659 VSS.n3059 VSS.t2419 9.3736
R6660 VSS.n3021 VSS.t455 9.3736
R6661 VSS.n1062 VSS.t1623 9.3736
R6662 VSS.n2461 VSS.t2261 9.3736
R6663 VSS.n2477 VSS.t1631 9.3736
R6664 VSS.n3423 VSS.t1064 9.3736
R6665 VSS.n1035 VSS.t437 9.3736
R6666 VSS.n3162 VSS.t439 9.3736
R6667 VSS.n931 VSS.t703 9.3736
R6668 VSS.n1173 VSS.t701 9.3736
R6669 VSS.n966 VSS.t2160 9.3736
R6670 VSS.n508 VSS.t1169 9.3736
R6671 VSS.n555 VSS.t1252 9.3736
R6672 VSS.n573 VSS.t1167 9.3736
R6673 VSS.n689 VSS.t1256 9.3736
R6674 VSS.n854 VSS.t2487 9.3736
R6675 VSS.n895 VSS.t2499 9.3736
R6676 VSS.n2649 VSS.t541 9.3736
R6677 VSS.n1646 VSS.t1319 9.3736
R6678 VSS.n1634 VSS.t870 9.3736
R6679 VSS.n1666 VSS.t1325 9.3736
R6680 VSS.n1495 VSS.n1494 9.37275
R6681 VSS.n3386 VSS.n3385 9.37275
R6682 VSS.n3382 VSS.n105 9.37275
R6683 VSS.n3291 VSS.n3290 9.37275
R6684 VSS.n123 VSS.n122 9.37275
R6685 VSS.n2508 VSS.n978 9.37275
R6686 VSS.n3011 VSS.n3010 9.37275
R6687 VSS.n3439 VSS.n35 9.37275
R6688 VSS.n460 VSS.n459 9.37275
R6689 VSS.n474 VSS.n473 9.37275
R6690 VSS.n443 VSS.n442 9.37275
R6691 VSS.n426 VSS.n421 9.37275
R6692 VSS.n1367 VSS.n1366 9.37275
R6693 VSS.n2333 VSS.n2317 9.37275
R6694 VSS.n2233 VSS.n2232 9.37275
R6695 VSS.n2250 VSS.n2224 9.37275
R6696 VSS.n2126 VSS.n2125 9.37275
R6697 VSS.n2082 VSS.n2081 9.37275
R6698 VSS.n2035 VSS.n2034 9.37275
R6699 VSS.n2219 VSS.n2006 9.37275
R6700 VSS.n1523 VSS.n1522 9.37275
R6701 VSS.n1514 VSS.n1513 9.37275
R6702 VSS.n521 VSS.n520 9.36649
R6703 VSS.n2848 VSS.n2847 9.36649
R6704 VSS.n976 VSS.t390 9.36521
R6705 VSS.n2577 VSS.t772 9.36521
R6706 VSS.n2607 VSS.t2253 9.3645
R6707 VSS.n619 VSS.t1519 9.3645
R6708 VSS.n1895 VSS.t53 9.364
R6709 VSS.n3086 VSS.t578 9.3533
R6710 VSS.n291 VSS.t986 9.3533
R6711 VSS.n3105 VSS.t1510 9.3533
R6712 VSS.n294 VSS.t1 9.35181
R6713 VSS.n3113 VSS.t142 9.35181
R6714 VSS.n262 VSS.n261 9.3508
R6715 VSS.n1183 VSS.t2440 9.34566
R6716 VSS.n3267 VSS.t386 9.34566
R6717 VSS.n3252 VSS.t280 9.34566
R6718 VSS.n3244 VSS.t1061 9.34566
R6719 VSS.n3237 VSS.t611 9.34566
R6720 VSS.n3234 VSS.t1021 9.34566
R6721 VSS.n3233 VSS.t2438 9.34566
R6722 VSS.n3242 VSS.t649 9.34566
R6723 VSS.n3250 VSS.t1340 9.34566
R6724 VSS.n3259 VSS.t100 9.34566
R6725 VSS.n1147 VSS.t1202 9.34566
R6726 VSS.n1155 VSS.t1214 9.34566
R6727 VSS.n1162 VSS.t2446 9.34566
R6728 VSS.n1137 VSS.t2444 9.34566
R6729 VSS.n1190 VSS.t2448 9.34566
R6730 VSS.n1194 VSS.t1212 9.34566
R6731 VSS.n226 VSS.n225 9.33837
R6732 VSS.n2611 VSS.n855 9.3221
R6733 VSS.n2609 VSS.t966 9.3221
R6734 VSS.n2605 VSS.n861 9.3221
R6735 VSS.n868 VSS.t1805 9.3221
R6736 VSS.n3326 VSS.t2422 9.3221
R6737 VSS.n3328 VSS.n3322 9.3221
R6738 VSS.n3308 VSS.t1080 9.3221
R6739 VSS.n3310 VSS.n3304 9.3221
R6740 VSS.n2516 VSS.n972 9.3221
R6741 VSS.n2514 VSS.t1797 9.3221
R6742 VSS.n2583 VSS.n2573 9.3221
R6743 VSS.n2581 VSS.t770 9.3221
R6744 VSS.n653 VSS.t2376 9.3221
R6745 VSS.n646 VSS.n645 9.3221
R6746 VSS.n407 VSS.t1074 9.3221
R6747 VSS.n400 VSS.n399 9.3221
R6748 VSS.n624 VSS.n608 9.3221
R6749 VSS.n628 VSS.t1580 9.3221
R6750 VSS.n613 VSS.n609 9.3221
R6751 VSS.n616 VSS.t972 9.3221
R6752 VSS.n3214 VSS.n232 9.3221
R6753 VSS.n1914 VSS.n1913 9.3221
R6754 VSS.n1921 VSS.t2221 9.3221
R6755 VSS.n1893 VSS.t9 9.3221
R6756 VSS.n1891 VSS.n1235 9.3221
R6757 VSS.n1531 VSS.n1530 9.3221
R6758 VSS.n1538 VSS.t2272 9.3221
R6759 VSS.n3089 VSS.t1727 9.31766
R6760 VSS.n304 VSS.t2303 9.31744
R6761 VSS.n3097 VSS.t235 9.31744
R6762 VSS.n907 VSS.t559 9.30652
R6763 VSS.n891 VSS.t1920 9.30652
R6764 VSS.n2612 VSS.t1845 9.30652
R6765 VSS.n860 VSS.t410 9.30652
R6766 VSS.n1732 VSS.n1731 9.30652
R6767 VSS.n1687 VSS.t1448 9.30652
R6768 VSS.n1707 VSS.t716 9.30652
R6769 VSS.n1997 VSS.t395 9.30652
R6770 VSS.n1993 VSS.t59 9.30652
R6771 VSS.n1989 VSS.t102 9.30652
R6772 VSS.n2181 VSS.t2509 9.30652
R6773 VSS.n1272 VSS.t865 9.30652
R6774 VSS.n1268 VSS.t291 9.30652
R6775 VSS.n1264 VSS.t1041 9.30652
R6776 VSS.n307 VSS.t1729 9.30652
R6777 VSS.n638 VSS.t2246 9.30652
R6778 VSS.n2429 VSS.t353 9.30652
R6779 VSS.n2441 VSS.t917 9.30652
R6780 VSS.n2437 VSS.t2176 9.30652
R6781 VSS.n3409 VSS.t94 9.30652
R6782 VSS.n3330 VSS.n3319 9.30652
R6783 VSS.n3325 VSS.n3323 9.30652
R6784 VSS.n3307 VSS.n3305 9.30652
R6785 VSS.n3312 VSS.n3301 9.30652
R6786 VSS.n3158 VSS.t1692 9.30652
R6787 VSS.n2517 VSS.t425 9.30652
R6788 VSS.n1389 VSS.n1388 9.30652
R6789 VSS.n1397 VSS.n1395 9.30652
R6790 VSS.n1402 VSS.n1394 9.30652
R6791 VSS.n2584 VSS.t1373 9.30652
R6792 VSS.n3446 VSS.t2450 9.30652
R6793 VSS.n654 VSS.n640 9.30652
R6794 VSS.n648 VSS.n641 9.30652
R6795 VSS.n402 VSS.n395 9.30652
R6796 VSS.n408 VSS.n394 9.30652
R6797 VSS.n682 VSS.t104 9.30652
R6798 VSS.n622 VSS.t392 9.30652
R6799 VSS.n612 VSS.t974 9.30652
R6800 VSS.n3486 VSS.t768 9.30652
R6801 VSS.n3482 VSS.t1136 9.30652
R6802 VSS.n322 VSS.n321 9.30652
R6803 VSS.n320 VSS.n312 9.30652
R6804 VSS.n318 VSS.n313 9.30652
R6805 VSS.n1421 VSS.t2538 9.30652
R6806 VSS.n2149 VSS.n2148 9.30652
R6807 VSS.n2162 VSS.n2154 9.30652
R6808 VSS.n2158 VSS.n2156 9.30652
R6809 VSS.n1922 VSS.n1908 9.30652
R6810 VSS.n1916 VSS.n1909 9.30652
R6811 VSS.n1890 VSS.t1745 9.30652
R6812 VSS.n1928 VSS.t495 9.30652
R6813 VSS.n1702 VSS.t919 9.30652
R6814 VSS.n1616 VSS.t1637 9.30652
R6815 VSS.n1611 VSS.t582 9.30652
R6816 VSS.n1607 VSS.t1504 9.30652
R6817 VSS.n1533 VSS.n1526 9.30652
R6818 VSS.n1539 VSS.n1525 9.30652
R6819 VSS.n332 VSS.t1974 9.30652
R6820 VSS.n2001 VSS.t863 9.30518
R6821 VSS.n1255 VSS.t459 9.30518
R6822 VSS.n2423 VSS.t237 9.30518
R6823 VSS.n1411 VSS.n1360 9.30518
R6824 VSS.n2941 VSS.t1984 9.30518
R6825 VSS.n2946 VSS.t85 9.30518
R6826 VSS.n2947 VSS.t586 9.30518
R6827 VSS.n2953 VSS.t584 9.30518
R6828 VSS.n2956 VSS.t1043 9.30518
R6829 VSS.n2962 VSS.t693 9.30518
R6830 VSS.n323 VSS.t811 9.30518
R6831 VSS.n3074 VSS.t809 9.30518
R6832 VSS.n7 VSS.t805 9.30518
R6833 VSS.n3484 VSS.t2298 9.30518
R6834 VSS.n2171 VSS.n2120 9.30518
R6835 VSS.n1704 VSS.t1498 9.30518
R6836 VSS.n1695 VSS.t920 9.30518
R6837 VSS.n1600 VSS.t1771 9.30518
R6838 VSS.n1692 VSS.t469 9.30323
R6839 VSS.n3491 VSS.t1972 9.30323
R6840 VSS.n665 VSS.t1350 9.30204
R6841 VSS.n877 VSS.t900 9.30204
R6842 VSS.n3476 VSS.t423 9.29981
R6843 VSS.n1713 VSS.t349 9.29981
R6844 VSS.n663 VSS.n657 9.29009
R6845 VSS.n661 VSS.t791 9.29009
R6846 VSS.n759 VSS.n758 9.29009
R6847 VSS.n2805 VSS.t313 9.29009
R6848 VSS.n3217 VSS.n3216 9.28776
R6849 VSS.n315 VSS.n314 9.26757
R6850 VSS.n3219 VSS.n228 9.26488
R6851 VSS.n227 VSS.n224 9.26488
R6852 VSS.n1999 VSS.t1598 9.25414
R6853 VSS.n1257 VSS.t867 9.25414
R6854 VSS.n2424 VSS.t385 9.25414
R6855 VSS.n1362 VSS.n1361 9.25414
R6856 VSS.n2122 VSS.n2121 9.25414
R6857 VSS.n1605 VSS.t1360 9.25414
R6858 VSS.n3159 VSS.n3158 9.19275
R6859 VSS.n1862 VSS.n1861 8.85568
R6860 VSS.t2374 VSS.t1982 8.76061
R6861 VSS.n3248 VSS.t784 8.70232
R6862 VSS.n3248 VSS.t785 8.70232
R6863 VSS.n1407 VSS.n1406 8.62119
R6864 VSS.n2167 VSS.n2166 8.62119
R6865 VSS.n1620 VSS.n1618 8.62119
R6866 VSS.n869 VSS.n866 7.39136
R6867 VSS.n626 VSS.n607 7.39136
R6868 VSS.n3409 VSS.n3408 7.3796
R6869 VSS.n1151 VSS.t15 7.36177
R6870 VSS VSS.n1527 7.30633
R6871 VSS VSS.t681 7.30633
R6872 VSS VSS.t879 7.30633
R6873 VSS VSS.n3320 7.30633
R6874 VSS VSS.n3302 7.30633
R6875 VSS VSS.t442 7.30633
R6876 VSS VSS.t2258 7.30633
R6877 VSS VSS.n1391 7.30633
R6878 VSS VSS.t695 7.30633
R6879 VSS VSS.n396 7.30633
R6880 VSS VSS.n642 7.30633
R6881 VSS VSS.n2151 7.30633
R6882 VSS VSS.n1910 7.30633
R6883 VSS VSS.t498 7.30633
R6884 VSS VSS.t873 7.30633
R6885 VSS.n867 VSS.t1804 7.19156
R6886 VSS.n1488 VSS.n1487 7.19156
R6887 VSS.n1841 VSS.n1489 7.19156
R6888 VSS.n1839 VSS.n1491 7.19156
R6889 VSS.n1741 VSS.n1726 7.19156
R6890 VSS.n1552 VSS.n1551 7.19156
R6891 VSS.n1757 VSS.n1546 7.19156
R6892 VSS.n1545 VSS.n1544 7.19156
R6893 VSS.n1479 VSS.t1662 7.19156
R6894 VSS.n1477 VSS.t1056 7.19156
R6895 VSS.n1475 VSS.t1050 7.19156
R6896 VSS.n1498 VSS.n1497 7.19156
R6897 VSS.n1501 VSS.n1500 7.19156
R6898 VSS.n1504 VSS.n1503 7.19156
R6899 VSS.n1935 VSS.t465 7.19156
R6900 VSS.n1937 VSS.t798 7.19156
R6901 VSS.n1225 VSS.t2135 7.19156
R6902 VSS.n1227 VSS.t462 7.19156
R6903 VSS.n1229 VSS.t147 7.19156
R6904 VSS.n2256 VSS.t912 7.19156
R6905 VSS.n1974 VSS.t1718 7.19156
R6906 VSS.n1093 VSS.t1609 7.19156
R6907 VSS.n1098 VSS.t1836 7.19156
R6908 VSS.n1099 VSS.t1549 7.19156
R6909 VSS.n2286 VSS.t580 7.19156
R6910 VSS.n2284 VSS.t306 7.19156
R6911 VSS.n2294 VSS.t180 7.19156
R6912 VSS.n2299 VSS.t624 7.19156
R6913 VSS.n2302 VSS.t2085 7.19156
R6914 VSS.n2344 VSS.t1777 7.19156
R6915 VSS.n1081 VSS.t68 7.19156
R6916 VSS.n2049 VSS.t87 7.19156
R6917 VSS.n2055 VSS.t840 7.19156
R6918 VSS.n2053 VSS.t845 7.19156
R6919 VSS.n2380 VSS.t1143 7.19156
R6920 VSS.n2378 VSS.t788 7.19156
R6921 VSS.n1438 VSS.t374 7.19156
R6922 VSS.n1436 VSS.t1800 7.19156
R6923 VSS.n1434 VSS.t1874 7.19156
R6924 VSS.n1280 VSS.t627 7.19156
R6925 VSS.n1285 VSS.t233 7.19156
R6926 VSS.n1244 VSS.t167 7.19156
R6927 VSS.n1459 VSS.t91 7.19156
R6928 VSS.n1293 VSS.t2194 7.19156
R6929 VSS.n1298 VSS.t229 7.19156
R6930 VSS.n1299 VSS.t851 7.19156
R6931 VSS.n1310 VSS.t1868 7.19156
R6932 VSS.n1315 VSS.t433 7.19156
R6933 VSS.n1318 VSS.t947 7.19156
R6934 VSS.n1452 VSS.t632 7.19156
R6935 VSS.n1450 VSS.t155 7.19156
R6936 VSS.n1953 VSS.t1496 7.19156
R6937 VSS.n1951 VSS.t842 7.19156
R6938 VSS.n1949 VSS.t477 7.19156
R6939 VSS.n1943 VSS.t320 7.19156
R6940 VSS.n1941 VSS.t1522 7.19156
R6941 VSS.n3069 VSS.t383 7.19156
R6942 VSS.n3067 VSS.t1568 7.19156
R6943 VSS.n16 VSS.t807 7.19156
R6944 VSS.n3022 VSS.t1925 7.19156
R6945 VSS.n3016 VSS.t41 7.19156
R6946 VSS.n3053 VSS.t1922 7.19156
R6947 VSS.n3051 VSS.t1371 7.19156
R6948 VSS.n2409 VSS.t2300 7.19156
R6949 VSS.n3206 VSS.t471 7.19156
R6950 VSS.n1007 VSS.t1993 7.19156
R6951 VSS.n1008 VSS.t475 7.19156
R6952 VSS.n1013 VSS.t2542 7.19156
R6953 VSS.n3199 VSS.t2251 7.19156
R6954 VSS.n3197 VSS.t195 7.19156
R6955 VSS.n2446 VSS.t301 7.19156
R6956 VSS.n2451 VSS.t198 7.19156
R6957 VSS.n2452 VSS.t241 7.19156
R6958 VSS.n3192 VSS.t133 7.19156
R6959 VSS.n3190 VSS.t1421 7.19156
R6960 VSS.n2465 VSS.t89 7.19156
R6961 VSS.n2470 VSS.t1417 7.19156
R6962 VSS.n2473 VSS.t1269 7.19156
R6963 VSS.n3183 VSS.t2256 7.19156
R6964 VSS.n3181 VSS.t793 7.19156
R6965 VSS.n76 VSS.n75 7.19156
R6966 VSS.n3402 VSS.n77 7.19156
R6967 VSS.n102 VSS.n101 7.19156
R6968 VSS.n99 VSS.n98 7.19156
R6969 VSS.n96 VSS.n95 7.19156
R6970 VSS.n81 VSS.n80 7.19156
R6971 VSS.n3375 VSS.n3372 7.19156
R6972 VSS.n90 VSS.n89 7.19156
R6973 VSS.n87 VSS.n86 7.19156
R6974 VSS.n84 VSS.n83 7.19156
R6975 VSS.n3365 VSS.n110 7.19156
R6976 VSS.n3362 VSS.n111 7.19156
R6977 VSS.n3342 VSS.n3298 7.19156
R6978 VSS.n3344 VSS.n3296 7.19156
R6979 VSS.n3346 VSS.n3294 7.19156
R6980 VSS.n115 VSS.n114 7.19156
R6981 VSS.n137 VSS.n134 7.19156
R6982 VSS.n3286 VSS.n118 7.19156
R6983 VSS.n120 VSS.n119 7.19156
R6984 VSS.n3281 VSS.n121 7.19156
R6985 VSS.n56 VSS.t662 7.19156
R6986 VSS.n61 VSS.t1969 7.19156
R6987 VSS.n62 VSS.t23 7.19156
R6988 VSS.n3148 VSS.t1649 7.19156
R6989 VSS.n3146 VSS.t1741 7.19156
R6990 VSS.n271 VSS.n268 7.19156
R6991 VSS.n273 VSS.n266 7.19156
R6992 VSS.n265 VSS.n264 7.19156
R6993 VSS.n2519 VSS.t1555 7.19156
R6994 VSS.n2524 VSS.t1297 7.19156
R6995 VSS.n1032 VSS.t1332 7.19156
R6996 VSS.n1034 VSS.t1879 7.19156
R6997 VSS.n1052 VSS.t640 7.19156
R6998 VSS.n2532 VSS.t1054 7.19156
R6999 VSS.n2538 VSS.t177 7.19156
R7000 VSS.n1037 VSS.t1401 7.19156
R7001 VSS.n1043 VSS.t175 7.19156
R7002 VSS.n1041 VSS.t355 7.19156
R7003 VSS.n990 VSS.n985 7.19156
R7004 VSS.n992 VSS.n983 7.19156
R7005 VSS.n994 VSS.n981 7.19156
R7006 VSS.n2479 VSS.t388 7.19156
R7007 VSS.n2481 VSS.t949 7.19156
R7008 VSS.n2483 VSS.t976 7.19156
R7009 VSS.n954 VSS.t1962 7.19156
R7010 VSS.n952 VSS.t162 7.19156
R7011 VSS.n919 VSS.t634 7.19156
R7012 VSS.n924 VSS.t159 7.19156
R7013 VSS.n927 VSS.t1570 7.19156
R7014 VSS.n2923 VSS.t381 7.19156
R7015 VSS.n2928 VSS.t190 7.19156
R7016 VSS.n934 VSS.t2095 7.19156
R7017 VSS.n936 VSS.t1046 7.19156
R7018 VSS.n938 VSS.t51 7.19156
R7019 VSS.n1019 VSS.t11 7.19156
R7020 VSS.n1021 VSS.t1612 7.19156
R7021 VSS.n1025 VSS.t594 7.19156
R7022 VSS.n3138 VSS.n283 7.19156
R7023 VSS.n3132 VSS.n284 7.19156
R7024 VSS.n3002 VSS.n2999 7.19156
R7025 VSS.n3004 VSS.n2997 7.19156
R7026 VSS.n2996 VSS.n2995 7.19156
R7027 VSS.n41 VSS.n39 7.19156
R7028 VSS.n43 VSS.n38 7.19156
R7029 VSS.n45 VSS.n37 7.19156
R7030 VSS.n31 VSS.n30 7.19156
R7031 VSS.n3432 VSS.n3429 7.19156
R7032 VSS.n3462 VSS.t712 7.19156
R7033 VSS.n3460 VSS.t710 7.19156
R7034 VSS.n3458 VSS.t1664 7.19156
R7035 VSS.n700 VSS.n381 7.19156
R7036 VSS.n704 VSS.n378 7.19156
R7037 VSS.n469 VSS.n387 7.19156
R7038 VSS.n389 VSS.n388 7.19156
R7039 VSS.n464 VSS.n390 7.19156
R7040 VSS.n656 VSS.n655 7.19156
R7041 VSS.n599 VSS.n589 7.19156
R7042 VSS.n486 VSS.n485 7.19156
R7043 VSS.n483 VSS.n482 7.19156
R7044 VSS.n480 VSS.n479 7.19156
R7045 VSS.n720 VSS.n367 7.19156
R7046 VSS.n723 VSS.n364 7.19156
R7047 VSS.n454 VSS.n412 7.19156
R7048 VSS.n451 VSS.n413 7.19156
R7049 VSS.n415 VSS.n414 7.19156
R7050 VSS.n737 VSS.n353 7.19156
R7051 VSS.n741 VSS.n350 7.19156
R7052 VSS.n435 VSS.n417 7.19156
R7053 VSS.n419 VSS.n418 7.19156
R7054 VSS.n430 VSS.n420 7.19156
R7055 VSS.n629 VSS.t1577 7.19156
R7056 VSS.n2983 VSS.t2345 7.19156
R7057 VSS.n2984 VSS.t1231 7.19156
R7058 VSS.n2989 VSS.t651 7.19156
R7059 VSS.n2549 VSS.t2155 7.19156
R7060 VSS.n2547 VSS.t2144 7.19156
R7061 VSS.n2545 VSS.t1696 7.19156
R7062 VSS.n2371 VSS.n2370 7.19156
R7063 VSS.n2373 VSS.n2368 7.19156
R7064 VSS.n1378 VSS.n1377 7.19156
R7065 VSS.n1375 VSS.n1374 7.19156
R7066 VSS.n1372 VSS.n1371 7.19156
R7067 VSS.n1080 VSS.n1079 7.19156
R7068 VSS.n2353 VSS.n2350 7.19156
R7069 VSS.n2326 VSS.n2325 7.19156
R7070 VSS.n2323 VSS.n2322 7.19156
R7071 VSS.n2320 VSS.n2319 7.19156
R7072 VSS.n2314 VSS.n1085 7.19156
R7073 VSS.n1087 VSS.n1086 7.19156
R7074 VSS.n1964 VSS.n1116 7.19156
R7075 VSS.n1966 VSS.n1114 7.19156
R7076 VSS.n1968 VSS.n1112 7.19156
R7077 VSS.n1973 VSS.n1972 7.19156
R7078 VSS.n2265 VSS.n2262 7.19156
R7079 VSS.n2240 VSS.n2231 7.19156
R7080 VSS.n2242 VSS.n2229 7.19156
R7081 VSS.n2244 VSS.n2227 7.19156
R7082 VSS.n2184 VSS.n2116 7.19156
R7083 VSS.n2186 VSS.n2114 7.19156
R7084 VSS.n2137 VSS.n2136 7.19156
R7085 VSS.n2134 VSS.n2133 7.19156
R7086 VSS.n2131 VSS.n2130 7.19156
R7087 VSS.n2193 VSS.n2107 7.19156
R7088 VSS.n2195 VSS.n2105 7.19156
R7089 VSS.n2093 VSS.n2092 7.19156
R7090 VSS.n2090 VSS.n2089 7.19156
R7091 VSS.n2087 VSS.n2086 7.19156
R7092 VSS.n2202 VSS.n2044 7.19156
R7093 VSS.n2204 VSS.n2042 7.19156
R7094 VSS.n2077 VSS.n2064 7.19156
R7095 VSS.n2066 VSS.n2065 7.19156
R7096 VSS.n2072 VSS.n2067 7.19156
R7097 VSS.n2211 VSS.n2030 7.19156
R7098 VSS.n2213 VSS.n2028 7.19156
R7099 VSS.n2017 VSS.n2013 7.19156
R7100 VSS.n2019 VSS.n2011 7.19156
R7101 VSS.n2021 VSS.n2009 7.19156
R7102 VSS.n2388 VSS.t815 7.19156
R7103 VSS.n2393 VSS.t1456 7.19156
R7104 VSS.n2396 VSS.t1743 7.19156
R7105 VSS.n1145 VSS.t2172 7.19156
R7106 VSS.n1145 VSS.t1537 7.19156
R7107 VSS.n1148 VSS.t1976 7.19156
R7108 VSS.n1153 VSS.t25 7.19156
R7109 VSS.n1153 VSS.t1502 7.19156
R7110 VSS.n1156 VSS.t2181 7.19156
R7111 VSS.n1161 VSS.t1791 7.19156
R7112 VSS.n1161 VSS.t622 7.19156
R7113 VSS.n1167 VSS.t752 7.19156
R7114 VSS.n1168 VSS.t1645 7.19156
R7115 VSS.n1168 VSS.t1275 7.19156
R7116 VSS.n1181 VSS.t2379 7.19156
R7117 VSS.n1182 VSS.t2289 7.19156
R7118 VSS.n1136 VSS.t2021 7.19156
R7119 VSS.n1136 VSS.t1344 7.19156
R7120 VSS.n1133 VSS.t2291 7.19156
R7121 VSS.n1192 VSS.t576 7.19156
R7122 VSS.n1192 VSS.t1778 7.19156
R7123 VSS.n1193 VSS.t1780 7.19156
R7124 VSS.n1128 VSS.t796 7.19156
R7125 VSS.n1128 VSS.t1750 7.19156
R7126 VSS.n1345 VSS.t2083 7.19156
R7127 VSS.n1343 VSS.t1029 7.19156
R7128 VSS.n1341 VSS.t1031 7.19156
R7129 VSS.n1336 VSS.t1506 7.19156
R7130 VSS.n1330 VSS.t736 7.19156
R7131 VSS.n1509 VSS.n1508 7.19156
R7132 VSS.n1823 VSS.n1510 7.19156
R7133 VSS.n1821 VSS.n1512 7.19156
R7134 VSS.n1777 VSS.n1518 7.19156
R7135 VSS.n1780 VSS.n1517 7.19156
R7136 VSS.n1803 VSS.n1802 7.19156
R7137 VSS.n1806 VSS.n1805 7.19156
R7138 VSS.n1809 VSS.n1808 7.19156
R7139 VSS.n1793 VSS.n1788 7.19156
R7140 VSS.n1791 VSS.n1790 7.19156
R7141 VSS.n2636 VSS.t149 7.19156
R7142 VSS.n2635 VSS.t2163 7.19156
R7143 VSS.n2630 VSS.t1352 7.19156
R7144 VSS.n816 VSS.t1826 7.19156
R7145 VSS.n818 VSS.t137 7.19156
R7146 VSS.n1640 VSS.t642 7.19156
R7147 VSS.n1638 VSS.t1998 7.19156
R7148 VSS.n1636 VSS.t620 7.19156
R7149 VSS.n800 VSS.t1995 7.19156
R7150 VSS.n795 VSS.t1635 7.19156
R7151 VSS.n1626 VSS.t414 7.19156
R7152 VSS.n1624 VSS.t667 7.19156
R7153 VSS.n1622 VSS.t834 7.19156
R7154 VSS.n1567 VSS.t1574 7.19156
R7155 VSS.n1569 VSS.t1889 7.19156
R7156 VSS.n1585 VSS.t691 7.19156
R7157 VSS.n1583 VSS.t1934 7.19156
R7158 VSS.n1581 VSS.t1937 7.19156
R7159 VSS.n1562 VSS.t108 7.19156
R7160 VSS.n1593 VSS.t1293 7.19156
R7161 VSS.n1873 VSS.t1295 7.19156
R7162 VSS.n1874 VSS.t1395 7.19156
R7163 VSS.n1879 VSS.t982 7.19156
R7164 VSS.n3044 VSS.t707 7.17823
R7165 VSS.n3040 VSS.t550 7.17823
R7166 VSS.n2685 VSS.t1784 7.17323
R7167 VSS.n2683 VSS.t1725 7.17323
R7168 VSS.n738 VSS.t1399 7.17323
R7169 VSS.n734 VSS.t2103 7.17323
R7170 VSS.n701 VSS.t1526 7.17323
R7171 VSS.n697 VSS.t1854 7.17323
R7172 VSS.n2660 VSS.t2293 7.17323
R7173 VSS.n2657 VSS.t836 7.17323
R7174 VSS.n3480 VSS.t2343 7.17156
R7175 VSS.n1709 VSS.t404 7.17156
R7176 VSS.n347 VSS.n346 7.17112
R7177 VSS.n719 VSS.t1885 7.16989
R7178 VSS.n715 VSS.t1281 7.16989
R7179 VSS.n2672 VSS.t341 7.16989
R7180 VSS.n2670 VSS.t1672 7.16989
R7181 VSS.n1684 VSS.t827 7.16656
R7182 VSS.n1681 VSS.t2311 7.16656
R7183 VSS.n752 VSS.t728 7.16656
R7184 VSS.n338 VSS.t1379 7.16656
R7185 VSS.n904 VSS.t402 7.16085
R7186 VSS.n678 VSS.t2341 7.16085
R7187 VSS.n677 VSS.t2336 7.15156
R7188 VSS.n902 VSS.t406 7.15156
R7189 VSS.n3417 VSS.n69 7.14989
R7190 VSS.n71 VSS.n70 7.14989
R7191 VSS.n3117 VSS.t999 7.14823
R7192 VSS.n3118 VSS.t996 7.14823
R7193 VSS.n2500 VSS.n1003 7.14489
R7194 VSS.n2502 VSS.n1001 7.14489
R7195 VSS.n3093 VSS.t412 7.13989
R7196 VSS.n3109 VSS.t1666 7.13989
R7197 VSS.n3110 VSS.t144 7.13989
R7198 VSS.n3094 VSS.t1508 7.13989
R7199 VSS.n1848 VSS.t297 7.13823
R7200 VSS.n1853 VSS.t1060 7.13823
R7201 VSS.n543 VSS.t1334 7.13489
R7202 VSS.n545 VSS.t2101 7.13489
R7203 VSS.n550 VSS.t1433 7.13489
R7204 VSS.n828 VSS.t467 7.13489
R7205 VSS.n829 VSS.t830 7.13489
R7206 VSS.n834 VSS.t2087 7.13489
R7207 VSS.n1470 VSS.t1389 7.13323
R7208 VSS.n1468 VSS.t1391 7.13323
R7209 VSS.n579 VSS.t1991 7.13323
R7210 VSS.n580 VSS.t1858 7.13323
R7211 VSS.n585 VSS.t131 7.13323
R7212 VSS.n879 VSS.t482 7.13323
R7213 VSS.n884 VSS.t479 7.13323
R7214 VSS.n885 VSS.t968 7.13323
R7215 VSS.n561 VSS.t603 7.13156
R7216 VSS.n563 VSS.t2140 7.13156
R7217 VSS.n568 VSS.t2322 7.13156
R7218 VSS.n844 VSS.t2091 7.13156
R7219 VSS.n845 VSS.t1676 7.13156
R7220 VSS.n850 VSS.t1710 7.13156
R7221 VSS.n1699 VSS.n1693 7.1285
R7222 VSS.n528 VSS.t1587 7.12823
R7223 VSS.n529 VSS.t2545 7.12823
R7224 VSS.n534 VSS.t2171 7.12823
R7225 VSS.n2696 VSS.t902 7.12823
R7226 VSS.n2694 VSS.t1787 7.12823
R7227 VSS.n2692 VSS.t1989 7.12823
R7228 VSS.n3101 VSS.t2301 7.12156
R7229 VSS.n3102 VSS.t315 7.12156
R7230 VSS.n2567 VSS.t429 7.11489
R7231 VSS.n2565 VSS.t1615 7.11489
R7232 VSS.n2558 VSS.t1699 7.11489
R7233 VSS.n285 VSS.t2142 7.11489
R7234 VSS.t138 VSS.n223 6.92477
R7235 VSS.t2285 VSS.n3222 6.92477
R7236 VSS.n1995 VSS.t2115 6.88656
R7237 VSS.n1991 VSS.t2015 6.88656
R7238 VSS.n2160 VSS.n2155 6.88656
R7239 VSS.n2164 VSS.n2150 6.88656
R7240 VSS.n1270 VSS.t2460 6.88656
R7241 VSS.n1266 VSS.t1038 6.88656
R7242 VSS.n2432 VSS.t1628 6.88656
R7243 VSS.n2439 VSS.t1339 6.88656
R7244 VSS.n1404 VSS.n1390 6.88656
R7245 VSS.n1400 VSS.n1399 6.88656
R7246 VSS.n1609 VSS.t1323 6.88656
R7247 VSS.n1612 VSS.t1893 6.88656
R7248 VSS.n1746 VSS.n1745 6.53419
R7249 VSS.n678 VSS.n677 6.41993
R7250 VSS.n3077 VSS.n3076 6.06679
R7251 VSS VSS.t408 6.02876
R7252 VSS VSS.t2338 6.02876
R7253 VSS.n1977 VSS.n1976 6.01414
R7254 VSS.n1977 VSS.t1950 6.01414
R7255 VSS.n1251 VSS.n1250 6.01414
R7256 VSS.n1251 VSS.t1832 6.01414
R7257 VSS.n1066 VSS.n1065 6.01414
R7258 VSS.n1066 VSS.t1810 6.01414
R7259 VSS.n1359 VSS.n1358 6.01414
R7260 VSS.n1359 VSS.t1896 6.01414
R7261 VSS.n2119 VSS.n2118 6.01414
R7262 VSS.n2119 VSS.t2199 6.01414
R7263 VSS.n1556 VSS.n1555 6.01414
R7264 VSS.n1556 VSS.t554 6.01414
R7265 VSS.n1591 VSS.n1590 6.01414
R7266 VSS.n1591 VSS.t2107 6.01414
R7267 VSS.n334 VSS.n333 6.01414
R7268 VSS.n334 VSS.t1979 6.01414
R7269 VSS.n3470 VSS.t1005 5.91497
R7270 VSS.n1729 VSS.n1728 5.91399
R7271 VSS.n1734 VSS.n1727 5.91399
R7272 VSS.n1736 VSS.n1735 5.91399
R7273 VSS.n1749 VSS.n1547 5.91399
R7274 VSS.n1751 VSS.n1750 5.91399
R7275 VSS.n1464 VSS.t522 5.91399
R7276 VSS.n1549 VSS.n1548 5.91399
R7277 VSS.n1931 VSS.t514 5.91399
R7278 VSS.n1933 VSS.t822 5.91399
R7279 VSS.n1125 VSS.t1235 5.91399
R7280 VSS.n2270 VSS.t1446 5.91399
R7281 VSS.n1105 VSS.t1093 5.91399
R7282 VSS.n1104 VSS.t61 5.91399
R7283 VSS.n1088 VSS.t106 5.91399
R7284 VSS.n2309 VSS.t1095 5.91399
R7285 VSS.n1089 VSS.t1103 5.91399
R7286 VSS.n2358 VSS.t980 5.91399
R7287 VSS.n1073 VSS.t1111 5.91399
R7288 VSS.n1072 VSS.t861 5.91399
R7289 VSS.n1068 VSS.t847 5.91399
R7290 VSS.n2406 VSS.t1116 5.91399
R7291 VSS.n1432 VSS.t2392 5.91399
R7292 VSS.n1249 VSS.t945 5.91399
R7293 VSS.n1290 VSS.t2396 5.91399
R7294 VSS.n1457 VSS.t1752 5.91399
R7295 VSS.n1455 VSS.t2404 5.91399
R7296 VSS.n1304 VSS.t849 5.91399
R7297 VSS.n1247 VSS.t2414 5.91399
R7298 VSS.n1448 VSS.t369 5.91399
R7299 VSS.n1121 VSS.t2394 5.91399
R7300 VSS.n1947 VSS.t1175 5.91399
R7301 VSS.n3064 VSS.t2165 5.91399
R7302 VSS.n3062 VSS.t274 5.91399
R7303 VSS.n3025 VSS.t1307 5.91399
R7304 VSS.n3031 VSS.t272 5.91399
R7305 VSS.n3049 VSS.t259 5.91399
R7306 VSS.n3204 VSS.t773 5.91399
R7307 VSS.n3202 VSS.t224 5.91399
R7308 VSS.n1014 VSS.t2540 5.91399
R7309 VSS.n249 VSS.t1589 5.91399
R7310 VSS.n2458 VSS.t219 5.91399
R7311 VSS.n2457 VSS.t217 5.91399
R7312 VSS.n3188 VSS.t714 5.91399
R7313 VSS.n3186 VSS.t215 5.91399
R7314 VSS.n2474 VSS.t1161 5.91399
R7315 VSS.n72 VSS.t1033 5.91399
R7316 VSS.n3412 VSS.t207 5.91399
R7317 VSS.n3397 VSS.n3396 5.91399
R7318 VSS.n3395 VSS.n78 5.91399
R7319 VSS.n93 VSS.n92 5.91399
R7320 VSS.n3377 VSS.n3370 5.91399
R7321 VSS.n3379 VSS.n109 5.91399
R7322 VSS.n107 VSS.n106 5.91399
R7323 VSS.n3357 VSS.n3356 5.91399
R7324 VSS.n3355 VSS.n112 5.91399
R7325 VSS.n3293 VSS.n3292 5.91399
R7326 VSS.n133 VSS.n132 5.91399
R7327 VSS.n130 VSS.n126 5.91399
R7328 VSS.n128 VSS.n127 5.91399
R7329 VSS.n67 VSS.t1479 5.91399
R7330 VSS.n51 VSS.t2089 5.91399
R7331 VSS.n3425 VSS.t1465 5.91399
R7332 VSS.n260 VSS.n259 5.91399
R7333 VSS.n970 VSS.t1585 5.91399
R7334 VSS.n2529 VSS.t1481 5.91399
R7335 VSS.n1050 VSS.t2547 5.91399
R7336 VSS.n2536 VSS.t962 5.91399
R7337 VSS.n279 VSS.t1472 5.91399
R7338 VSS.n278 VSS.t2204 5.91399
R7339 VSS.n996 VSS.n979 5.91399
R7340 VSS.n73 VSS.t205 5.91399
R7341 VSS.n3240 VSS.t1205 5.91399
R7342 VSS.n3240 VSS.t1204 5.91399
R7343 VSS.n3256 VSS.t359 5.91399
R7344 VSS.n3256 VSS.t360 5.91399
R7345 VSS.n3264 VSS.t357 5.91399
R7346 VSS.n3264 VSS.t786 5.91399
R7347 VSS.n950 VSS.t1300 5.91399
R7348 VSS.n328 VSS.t248 5.91399
R7349 VSS.n928 VSS.t286 5.91399
R7350 VSS.n326 VSS.t289 5.91399
R7351 VSS.n2935 VSS.t250 5.91399
R7352 VSS.n939 VSS.t749 5.91399
R7353 VSS.n1023 VSS.t1458 5.91399
R7354 VSS.n3122 VSS.n3121 5.91399
R7355 VSS.n3120 VSS.n286 5.91399
R7356 VSS.n2993 VSS.n2992 5.91399
R7357 VSS.n47 VSS.n36 5.91399
R7358 VSS.n3434 VSS.n50 5.91399
R7359 VSS.n3436 VSS.n48 5.91399
R7360 VSS.n3456 VSS.t267 5.91399
R7361 VSS.n707 VSS.n375 5.91399
R7362 VSS.n711 VSS.n372 5.91399
R7363 VSS.n392 VSS.n391 5.91399
R7364 VSS.n596 VSS.n590 5.91399
R7365 VSS.n592 VSS.n591 5.91399
R7366 VSS.n477 VSS.n475 5.91399
R7367 VSS.n728 VSS.n360 5.91399
R7368 VSS.n732 VSS.n357 5.91399
R7369 VSS.n446 VSS.n445 5.91399
R7370 VSS.n745 VSS.n344 5.91399
R7371 VSS.n341 VSS.n340 5.91399
R7372 VSS.n423 VSS.n422 5.91399
R7373 VSS.n2975 VSS.t254 5.91399
R7374 VSS.n3152 VSS.t1463 5.91399
R7375 VSS.n1423 VSS.t1887 5.91399
R7376 VSS.n1430 VSS.t2406 5.91399
R7377 VSS.n2367 VSS.n1076 5.91399
R7378 VSS.n2364 VSS.n1077 5.91399
R7379 VSS.n1369 VSS.n1368 5.91399
R7380 VSS.n2349 VSS.n1082 5.91399
R7381 VSS.n2336 VSS.n2335 5.91399
R7382 VSS.n2316 VSS.n2315 5.91399
R7383 VSS.n2279 VSS.n1108 5.91399
R7384 VSS.n2276 VSS.n1109 5.91399
R7385 VSS.n1970 VSS.n1110 5.91399
R7386 VSS.n2261 VSS.n1975 5.91399
R7387 VSS.n2248 VSS.n2247 5.91399
R7388 VSS.n2246 VSS.n2225 5.91399
R7389 VSS.n2188 VSS.n2112 5.91399
R7390 VSS.n2190 VSS.n2110 5.91399
R7391 VSS.n2128 VSS.n2127 5.91399
R7392 VSS.n2197 VSS.n2103 5.91399
R7393 VSS.n2199 VSS.n2047 5.91399
R7394 VSS.n2084 VSS.n2083 5.91399
R7395 VSS.n2206 VSS.n2040 5.91399
R7396 VSS.n2208 VSS.n2033 5.91399
R7397 VSS.n2069 VSS.n2068 5.91399
R7398 VSS.n2215 VSS.n2026 5.91399
R7399 VSS.n2217 VSS.n2024 5.91399
R7400 VSS.n2023 VSS.n2007 5.91399
R7401 VSS.n2397 VSS.t1088 5.91399
R7402 VSS.n1347 VSS.t1617 5.91399
R7403 VSS.n1350 VSS.t520 5.91399
R7404 VSS.n1339 VSS.t1660 5.91399
R7405 VSS.n1521 VSS.n1520 5.91399
R7406 VSS.n1767 VSS.n1519 5.91399
R7407 VSS.n1769 VSS.n1768 5.91399
R7408 VSS.n1800 VSS.n1515 5.91399
R7409 VSS.n1797 VSS.n1516 5.91399
R7410 VSS.n1795 VSS.n1786 5.91399
R7411 VSS.n2641 VSS.t1012 5.91399
R7412 VSS.n2647 VSS.t1010 5.91399
R7413 VSS.n2644 VSS.t376 5.91399
R7414 VSS.n1648 VSS.t1247 5.91399
R7415 VSS.n1643 VSS.t1018 5.91399
R7416 VSS.n805 VSS.t978 5.91399
R7417 VSS.n1628 VSS.t1008 5.91399
R7418 VSS.n1631 VSS.t1014 5.91399
R7419 VSS.n785 VSS.t1342 5.91399
R7420 VSS.n1577 VSS.t690 5.91399
R7421 VSS.n1669 VSS.t1016 5.91399
R7422 VSS.n1672 VSS.t618 5.91399
R7423 VSS.n1880 VSS.t518 5.91399
R7424 VSS.n3037 VSS.t192 5.90065
R7425 VSS.n3454 VSS.t252 5.90065
R7426 VSS.n3478 VSS.t1133 5.89898
R7427 VSS.n1715 VSS.t1735 5.89898
R7428 VSS.n2680 VSS.t1362 5.89565
R7429 VSS.n2677 VSS.t1412 5.89565
R7430 VSS.n692 VSS.t184 5.89565
R7431 VSS.n729 VSS.t1668 5.89565
R7432 VSS.n725 VSS.t2126 5.89565
R7433 VSS.n2655 VSS.t571 5.89565
R7434 VSS.n897 VSS.t1377 5.89565
R7435 VSS.n712 VSS.t2137 5.89232
R7436 VSS.n708 VSS.t2369 5.89232
R7437 VSS.n2667 VSS.t766 5.89232
R7438 VSS.n2664 VSS.t2306 5.89232
R7439 VSS.n1678 VSS.t1685 5.88898
R7440 VSS.n777 VSS.t1681 5.88898
R7441 VSS.n342 VSS.t63 5.88898
R7442 VSS.n744 VSS.t2169 5.88898
R7443 VSS.n3176 VSS.n257 5.87232
R7444 VSS.n3173 VSS.n258 5.87232
R7445 VSS.n2504 VSS.n999 5.86732
R7446 VSS.n2506 VSS.n997 5.86732
R7447 VSS.n1856 VSS.t153 5.86065
R7448 VSS.n1465 VSS.t516 5.86065
R7449 VSS.n553 VSS.t2124 5.85732
R7450 VSS.n835 VSS.t1410 5.85732
R7451 VSS.n1237 VSS.t1939 5.85565
R7452 VSS.n1886 VSS.t512 5.85565
R7453 VSS.n498 VSS.t182 5.85565
R7454 VSS.n890 VSS.t1375 5.85565
R7455 VSS.n571 VSS.t2367 5.85398
R7456 VSS.n851 VSS.t2308 5.85398
R7457 VSS.n535 VSS.t2167 5.85065
R7458 VSS.n2690 VSS.t1683 5.85065
R7459 VSS.n2563 VSS.t761 5.83732
R7460 VSS.n2561 VSS.t1474 5.83732
R7461 VSS.n3127 VSS.t30 5.83732
R7462 VSS.n282 VSS.t1470 5.83732
R7463 VSS.n3079 VSS.n3078 5.82215
R7464 VSS.n2849 VSS.n2848 5.68397
R7465 VSS.n904 VSS.n903 5.43892
R7466 VSS.n6 VSS.n4 5.4332
R7467 VSS.n2569 VSS 5.34271
R7468 VSS.n2940 VSS.n2939 5.27581
R7469 VSS.n251 VSS.t2284 5.21719
R7470 VSS.n1000 VSS.t1418 5.21719
R7471 VSS.n252 VSS.t1550 5.21719
R7472 VSS.n1002 VSS.t2263 5.21719
R7473 VSS VSS.n659 5.20234
R7474 VSS.n2807 VSS 5.20234
R7475 VSS.n574 VSS 5.20137
R7476 VSS.n2619 VSS 5.20137
R7477 VSS.t610 VSS 5.20126
R7478 VSS.n872 VSS.n871 5.2005
R7479 VSS.n905 VSS.n874 5.2005
R7480 VSS.n909 VSS.n908 5.2005
R7481 VSS.n864 VSS.n863 5.2005
R7482 VSS.n859 VSS.n858 5.2005
R7483 VSS.n2608 VSS.n857 5.2005
R7484 VSS.n2614 VSS.n2613 5.2005
R7485 VSS.n2610 VSS.n856 5.2005
R7486 VSS.n1481 VSS.n1480 5.2005
R7487 VSS.n1478 VSS.n1471 5.2005
R7488 VSS.n1476 VSS.n1472 5.2005
R7489 VSS.n1474 VSS.n1473 5.2005
R7490 VSS.n1832 VSS.n1496 5.2005
R7491 VSS.n1831 VSS.n1499 5.2005
R7492 VSS.n1830 VSS.n1502 5.2005
R7493 VSS.n1829 VSS.n1505 5.2005
R7494 VSS.n1988 VSS.n1987 5.2005
R7495 VSS.n1990 VSS.n1986 5.2005
R7496 VSS.n1992 VSS.n1985 5.2005
R7497 VSS.n1994 VSS.n1984 5.2005
R7498 VSS.n1996 VSS.n1983 5.2005
R7499 VSS.n1998 VSS.n1982 5.2005
R7500 VSS.n2000 VSS.n1981 5.2005
R7501 VSS.n2002 VSS.n1980 5.2005
R7502 VSS.n2004 VSS.n1979 5.2005
R7503 VSS.n1278 VSS.n1277 5.2005
R7504 VSS.n1276 VSS.n1254 5.2005
R7505 VSS.n1275 VSS.n1256 5.2005
R7506 VSS.n1274 VSS.n1273 5.2005
R7507 VSS.n1271 VSS.n1258 5.2005
R7508 VSS.n1265 VSS.n1261 5.2005
R7509 VSS.n1263 VSS.n1262 5.2005
R7510 VSS.n1267 VSS.n1260 5.2005
R7511 VSS.n1269 VSS.n1259 5.2005
R7512 VSS.n1295 VSS.n1294 5.2005
R7513 VSS.n1297 VSS.n1296 5.2005
R7514 VSS.n1301 VSS.n1300 5.2005
R7515 VSS.n1303 VSS.n1302 5.2005
R7516 VSS.n1307 VSS.n1306 5.2005
R7517 VSS.n1312 VSS.n1311 5.2005
R7518 VSS.n1314 VSS.n1313 5.2005
R7519 VSS.n1317 VSS.n1316 5.2005
R7520 VSS.n1320 VSS.n1319 5.2005
R7521 VSS.n1282 VSS.n1281 5.2005
R7522 VSS.n1284 VSS.n1283 5.2005
R7523 VSS.n1287 VSS.n1286 5.2005
R7524 VSS.n1289 VSS.n1288 5.2005
R7525 VSS.n3332 VSS.n3331 5.2005
R7526 VSS.n3324 VSS.n3318 5.2005
R7527 VSS.n3306 VSS.n3300 5.2005
R7528 VSS.n3314 VSS.n3313 5.2005
R7529 VSS.n3383 VSS.n3382 5.2005
R7530 VSS.n3341 VSS.n3340 5.2005
R7531 VSS.n3343 VSS.n3297 5.2005
R7532 VSS.n3345 VSS.n3295 5.2005
R7533 VSS.n3348 VSS.n3347 5.2005
R7534 VSS.n3349 VSS.n3291 5.2005
R7535 VSS.n3288 VSS.n3287 5.2005
R7536 VSS.n3285 VSS.n3284 5.2005
R7537 VSS.n3283 VSS.n3282 5.2005
R7538 VSS.n3280 VSS.n3279 5.2005
R7539 VSS.n3277 VSS.n123 5.2005
R7540 VSS.n140 VSS.n131 5.2005
R7541 VSS.n139 VSS.n138 5.2005
R7542 VSS.n136 VSS.n135 5.2005
R7543 VSS.n3353 VSS.n3352 5.2005
R7544 VSS.n3359 VSS.n3358 5.2005
R7545 VSS.n3361 VSS.n3360 5.2005
R7546 VSS.n3364 VSS.n3363 5.2005
R7547 VSS.n3367 VSS.n3366 5.2005
R7548 VSS.n3378 VSS.n3369 5.2005
R7549 VSS.n3376 VSS.n3371 5.2005
R7550 VSS.n3374 VSS.n3373 5.2005
R7551 VSS.n3393 VSS.n3392 5.2005
R7552 VSS.n3399 VSS.n3398 5.2005
R7553 VSS.n3401 VSS.n3400 5.2005
R7554 VSS.n3404 VSS.n3403 5.2005
R7555 VSS.n3407 VSS.n3406 5.2005
R7556 VSS.n3390 VSS.n103 5.2005
R7557 VSS.n3390 VSS.n100 5.2005
R7558 VSS.n3390 VSS.n97 5.2005
R7559 VSS.n3390 VSS.n94 5.2005
R7560 VSS.n3388 VSS.n3386 5.2005
R7561 VSS.n3390 VSS.n91 5.2005
R7562 VSS.n3390 VSS.n88 5.2005
R7563 VSS.n3390 VSS.n85 5.2005
R7564 VSS.n3390 VSS.n82 5.2005
R7565 VSS.n2528 VSS.n2527 5.2005
R7566 VSS.n2526 VSS.n2525 5.2005
R7567 VSS.n2523 VSS.n2522 5.2005
R7568 VSS.n2521 VSS.n2520 5.2005
R7569 VSS.n989 VSS.n988 5.2005
R7570 VSS.n991 VSS.n984 5.2005
R7571 VSS.n993 VSS.n982 5.2005
R7572 VSS.n995 VSS.n980 5.2005
R7573 VSS.n2505 VSS.n998 5.2005
R7574 VSS.n2503 VSS.n1000 5.2005
R7575 VSS.n2501 VSS.n1002 5.2005
R7576 VSS.n2499 VSS.n2498 5.2005
R7577 VSS.n3175 VSS.n3174 5.2005
R7578 VSS.n3178 VSS.n3177 5.2005
R7579 VSS.n3416 VSS.n3415 5.2005
R7580 VSS.n3419 VSS.n3418 5.2005
R7581 VSS.n276 VSS.n263 5.2005
R7582 VSS.n275 VSS.n274 5.2005
R7583 VSS.n272 VSS.n267 5.2005
R7584 VSS.n270 VSS.n269 5.2005
R7585 VSS.n3423 VSS.n3422 5.2005
R7586 VSS.n58 VSS.n57 5.2005
R7587 VSS.n60 VSS.n59 5.2005
R7588 VSS.n64 VSS.n63 5.2005
R7589 VSS.n66 VSS.n65 5.2005
R7590 VSS.n3170 VSS.n3169 5.2005
R7591 VSS.n3410 VSS.n74 5.2005
R7592 VSS.n2485 VSS.n2484 5.2005
R7593 VSS.n2486 VSS.n2482 5.2005
R7594 VSS.n2487 VSS.n2480 5.2005
R7595 VSS.n2488 VSS.n2478 5.2005
R7596 VSS.n3414 VSS.n3413 5.2005
R7597 VSS.n3180 VSS.n3179 5.2005
R7598 VSS.n3182 VSS.n256 5.2005
R7599 VSS.n3184 VSS.n255 5.2005
R7600 VSS.n3187 VSS.n253 5.2005
R7601 VSS.n3189 VSS.n252 5.2005
R7602 VSS.n3191 VSS.n251 5.2005
R7603 VSS.n3208 VSS.n3207 5.2005
R7604 VSS.n2410 VSS.n237 5.2005
R7605 VSS.n3196 VSS.n3195 5.2005
R7606 VSS.n3198 VSS.n246 5.2005
R7607 VSS.n3200 VSS.n245 5.2005
R7608 VSS.n2515 VSS.n973 5.2005
R7609 VSS.n2518 VSS.n971 5.2005
R7610 VSS.n2512 VSS.n2511 5.2005
R7611 VSS.n975 VSS.n974 5.2005
R7612 VSS.n3194 VSS.n3193 5.2005
R7613 VSS.n3194 VSS.n250 5.2005
R7614 VSS.n2509 VSS.n2508 5.2005
R7615 VSS.n2448 VSS.n2447 5.2005
R7616 VSS.n2450 VSS.n2449 5.2005
R7617 VSS.n2454 VSS.n2453 5.2005
R7618 VSS.n2456 VSS.n2455 5.2005
R7619 VSS.n2462 VSS.n2461 5.2005
R7620 VSS.n2467 VSS.n2466 5.2005
R7621 VSS.n2469 VSS.n2468 5.2005
R7622 VSS.n2472 VSS.n2471 5.2005
R7623 VSS.n2476 VSS.n2475 5.2005
R7624 VSS.n2493 VSS.n2477 5.2005
R7625 VSS.n2436 VSS.n2435 5.2005
R7626 VSS.n2438 VSS.n2434 5.2005
R7627 VSS.n2440 VSS.n2433 5.2005
R7628 VSS.n2443 VSS.n2442 5.2005
R7629 VSS.n2431 VSS.n2430 5.2005
R7630 VSS.n2428 VSS.n2427 5.2005
R7631 VSS.n2426 VSS.n2425 5.2005
R7632 VSS.n2422 VSS.n2421 5.2005
R7633 VSS.n2419 VSS.n2418 5.2005
R7634 VSS.n3262 VSS.n3261 5.2005
R7635 VSS.n2413 VSS.n2412 5.2005
R7636 VSS.t99 VSS.n3268 5.2005
R7637 VSS.t99 VSS.n3258 5.2005
R7638 VSS.t648 VSS.n3245 5.2005
R7639 VSS.t279 VSS.n3253 5.2005
R7640 VSS.t648 VSS.n3243 5.2005
R7641 VSS.t279 VSS.n3251 5.2005
R7642 VSS.n1393 VSS.n1392 5.2005
R7643 VSS.n1406 VSS.n1405 5.2005
R7644 VSS.n1403 VSS.n1393 5.2005
R7645 VSS.n1396 VSS.n1363 5.2005
R7646 VSS.n1418 VSS.n1417 5.2005
R7647 VSS.n1415 VSS.n1414 5.2005
R7648 VSS.n1410 VSS.n1409 5.2005
R7649 VSS.n2961 VSS.n2960 5.2005
R7650 VSS.n2955 VSS.n2954 5.2005
R7651 VSS.n2958 VSS.n2957 5.2005
R7652 VSS.n2952 VSS.n2951 5.2005
R7653 VSS.n2949 VSS.n2948 5.2005
R7654 VSS.n2943 VSS.n2942 5.2005
R7655 VSS.n1006 VSS.n1005 5.2005
R7656 VSS.n1010 VSS.n1009 5.2005
R7657 VSS.n1012 VSS.n1011 5.2005
R7658 VSS.n1016 VSS.n1015 5.2005
R7659 VSS.n1063 VSS.n1062 5.2005
R7660 VSS.n1029 VSS.n1018 5.2005
R7661 VSS.n1028 VSS.n1020 5.2005
R7662 VSS.n1027 VSS.n1026 5.2005
R7663 VSS.n1024 VSS.n1022 5.2005
R7664 VSS.n967 VSS.n966 5.2005
R7665 VSS.n3203 VSS.n242 5.2005
R7666 VSS.n1046 VSS.n1036 5.2005
R7667 VSS.n1045 VSS.n1044 5.2005
R7668 VSS.n1042 VSS.n1038 5.2005
R7669 VSS.n1040 VSS.n1039 5.2005
R7670 VSS.n1056 VSS.n1031 5.2005
R7671 VSS.n1055 VSS.n1033 5.2005
R7672 VSS.n1054 VSS.n1053 5.2005
R7673 VSS.n1051 VSS.n1049 5.2005
R7674 VSS.n1048 VSS.n1035 5.2005
R7675 VSS.n2535 VSS.n2534 5.2005
R7676 VSS.n2537 VSS.n2533 5.2005
R7677 VSS.n2540 VSS.n2539 5.2005
R7678 VSS.n2541 VSS.n2531 5.2005
R7679 VSS.n3163 VSS.n3162 5.2005
R7680 VSS.n3157 VSS.n3156 5.2005
R7681 VSS.n3001 VSS.n3000 5.2005
R7682 VSS.n3003 VSS.n2998 5.2005
R7683 VSS.n3006 VSS.n3005 5.2005
R7684 VSS.n3007 VSS.n2994 5.2005
R7685 VSS.n3124 VSS.n3123 5.2005
R7686 VSS.n3131 VSS.n3130 5.2005
R7687 VSS.n3137 VSS.n3136 5.2005
R7688 VSS.n3464 VSS.n3463 5.2005
R7689 VSS.n3461 VSS.n26 5.2005
R7690 VSS.n3459 VSS.n27 5.2005
R7691 VSS.n3457 VSS.n28 5.2005
R7692 VSS.n3043 VSS.n3042 5.2005
R7693 VSS.n3038 VSS.n3036 5.2005
R7694 VSS.n3039 VSS.n3034 5.2005
R7695 VSS.n3045 VSS.n3033 5.2005
R7696 VSS.n3046 VSS.n3032 5.2005
R7697 VSS.n40 VSS.n34 5.2005
R7698 VSS.n42 VSS.n34 5.2005
R7699 VSS.n44 VSS.n34 5.2005
R7700 VSS.n46 VSS.n34 5.2005
R7701 VSS.n3440 VSS.n3439 5.2005
R7702 VSS.n3427 VSS.n3426 5.2005
R7703 VSS.n3145 VSS.n3144 5.2005
R7704 VSS.n3147 VSS.n3143 5.2005
R7705 VSS.n3149 VSS.n3141 5.2005
R7706 VSS.n3140 VSS.n3139 5.2005
R7707 VSS.n3435 VSS.n49 5.2005
R7708 VSS.n3433 VSS.n3428 5.2005
R7709 VSS.n3431 VSS.n3430 5.2005
R7710 VSS.n3445 VSS.n3444 5.2005
R7711 VSS.n3448 VSS.n3447 5.2005
R7712 VSS.n3453 VSS.n3452 5.2005
R7713 VSS.n3035 VSS.n29 5.2005
R7714 VSS.n509 VSS.n508 5.2005
R7715 VSS.n751 VSS.n750 5.2005
R7716 VSS.n753 VSS.n337 5.2005
R7717 VSS.n527 VSS.n526 5.2005
R7718 VSS.n531 VSS.n530 5.2005
R7719 VSS.n533 VSS.n532 5.2005
R7720 VSS.n537 VSS.n536 5.2005
R7721 VSS.n542 VSS.n541 5.2005
R7722 VSS.n547 VSS.n546 5.2005
R7723 VSS.n549 VSS.n548 5.2005
R7724 VSS.n552 VSS.n551 5.2005
R7725 VSS.n652 VSS.n651 5.2005
R7726 VSS.n644 VSS.n643 5.2005
R7727 VSS.n671 VSS.n670 5.2005
R7728 VSS.n650 VSS.n649 5.2005
R7729 VSS.n398 VSS.n397 5.2005
R7730 VSS.n404 VSS.n403 5.2005
R7731 VSS.n406 VSS.n405 5.2005
R7732 VSS.n410 VSS.n409 5.2005
R7733 VSS.n746 VSS.n343 5.2005
R7734 VSS.n749 VSS.n339 5.2005
R7735 VSS.n743 VSS.n348 5.2005
R7736 VSS.n748 VSS.n747 5.2005
R7737 VSS.n689 VSS.n688 5.2005
R7738 VSS.n686 VSS.n600 5.2005
R7739 VSS.n676 VSS.n675 5.2005
R7740 VSS.n662 VSS.n658 5.2005
R7741 VSS.n667 VSS.n666 5.2005
R7742 VSS.n669 VSS.n668 5.2005
R7743 VSS.n602 VSS.n601 5.2005
R7744 VSS.n679 VSS.n639 5.2005
R7745 VSS.n637 VSS.n636 5.2005
R7746 VSS.n611 VSS.n610 5.2005
R7747 VSS.n615 VSS.n614 5.2005
R7748 VSS.n684 VSS.n683 5.2005
R7749 VSS.n605 VSS.n604 5.2005
R7750 VSS.n621 VSS.n620 5.2005
R7751 VSS.n618 VSS.n617 5.2005
R7752 VSS.n3021 VSS.n3020 5.2005
R7753 VSS.n3056 VSS.n3015 5.2005
R7754 VSS.n3055 VSS.n3054 5.2005
R7755 VSS.n3052 VSS.n3017 5.2005
R7756 VSS.n3050 VSS.n3018 5.2005
R7757 VSS.n3075 VSS.n2965 5.2005
R7758 VSS.n2964 VSS.n2963 5.2005
R7759 VSS.n3 VSS.n2 5.2005
R7760 VSS.n3488 VSS.n3487 5.2005
R7761 VSS.n3485 VSS.n5 5.2005
R7762 VSS.n3483 VSS.n8 5.2005
R7763 VSS.n3475 VSS.n3474 5.2005
R7764 VSS.n3477 VSS.n13 5.2005
R7765 VSS.n3479 VSS.n11 5.2005
R7766 VSS.n3481 VSS.n9 5.2005
R7767 VSS.n556 VSS.n555 5.2005
R7768 VSS.n560 VSS.n559 5.2005
R7769 VSS.n565 VSS.n564 5.2005
R7770 VSS.n567 VSS.n566 5.2005
R7771 VSS.n570 VSS.n569 5.2005
R7772 VSS.n593 VSS.n496 5.2005
R7773 VSS.n695 VSS.n495 5.2005
R7774 VSS.n698 VSS.n383 5.2005
R7775 VSS.n702 VSS.n380 5.2005
R7776 VSS.n598 VSS.n597 5.2005
R7777 VSS.n595 VSS.n594 5.2005
R7778 VSS.n699 VSS.n382 5.2005
R7779 VSS.n703 VSS.n379 5.2005
R7780 VSS.n578 VSS.n577 5.2005
R7781 VSS.n582 VSS.n581 5.2005
R7782 VSS.n584 VSS.n583 5.2005
R7783 VSS.n587 VSS.n586 5.2005
R7784 VSS.n3469 VSS.n15 5.2005
R7785 VSS.n3468 VSS.n17 5.2005
R7786 VSS.n3024 VSS.n3023 5.2005
R7787 VSS.n3030 VSS.n3029 5.2005
R7788 VSS.n3027 VSS.n3026 5.2005
R7789 VSS.n3470 VSS.n14 5.2005
R7790 VSS.n3059 VSS.n3058 5.2005
R7791 VSS.n2982 VSS.n2981 5.2005
R7792 VSS.n2986 VSS.n2985 5.2005
R7793 VSS.n2988 VSS.n2987 5.2005
R7794 VSS.n2991 VSS.n2990 5.2005
R7795 VSS.n3070 VSS.n2967 5.2005
R7796 VSS.n3068 VSS.n2971 5.2005
R7797 VSS.n3065 VSS.n2973 5.2005
R7798 VSS.n3063 VSS.n2974 5.2005
R7799 VSS.n3071 VSS.n2966 5.2005
R7800 VSS.n3066 VSS.n2972 5.2005
R7801 VSS.n319 VSS.n309 5.2005
R7802 VSS.n226 VSS.n223 5.2005
R7803 VSS.n3222 VSS.n3220 5.2005
R7804 VSS.n3213 VSS.n3212 5.2005
R7805 VSS.n234 VSS.n233 5.2005
R7806 VSS.n231 VSS.n230 5.2005
R7807 VSS.n3205 VSS.n238 5.2005
R7808 VSS.n3082 VSS.n308 5.2005
R7809 VSS.n3086 VSS.n3085 5.2005
R7810 VSS.n3090 VSS.n3089 5.2005
R7811 VSS.n3092 VSS.n3091 5.2005
R7812 VSS.n304 VSS.n303 5.2005
R7813 VSS.n3100 VSS.n3099 5.2005
R7814 VSS.n3098 VSS.n3097 5.2005
R7815 VSS.n293 VSS.n289 5.2005
R7816 VSS.n292 VSS.n291 5.2005
R7817 VSS.n3108 VSS.n3107 5.2005
R7818 VSS.n3106 VSS.n3105 5.2005
R7819 VSS.n296 VSS.n288 5.2005
R7820 VSS.n295 VSS.n294 5.2005
R7821 VSS.n3116 VSS.n3115 5.2005
R7822 VSS.n3114 VSS.n3113 5.2005
R7823 VSS.n3012 VSS.n3011 5.2005
R7824 VSS.n2551 VSS.n2550 5.2005
R7825 VSS.n2548 VSS.n2543 5.2005
R7826 VSS.n2546 VSS.n2544 5.2005
R7827 VSS.n3154 VSS.n3153 5.2005
R7828 VSS.n3129 VSS.n3128 5.2005
R7829 VSS.n3126 VSS.n3125 5.2005
R7830 VSS.n2557 VSS.n2556 5.2005
R7831 VSS.n2559 VSS.n2556 5.2005
R7832 VSS.n2562 VSS.n964 5.2005
R7833 VSS.n2564 VSS.n961 5.2005
R7834 VSS.n2566 VSS.n960 5.2005
R7835 VSS.n2568 VSS.n959 5.2005
R7836 VSS.n2403 VSS.n1069 5.2005
R7837 VSS.n2153 VSS.n2152 5.2005
R7838 VSS.n2166 VSS.n2165 5.2005
R7839 VSS.n2163 VSS.n2153 5.2005
R7840 VSS.n2157 VSS.n2123 5.2005
R7841 VSS.n2170 VSS.n2169 5.2005
R7842 VSS.n2175 VSS.n2174 5.2005
R7843 VSS.n2178 VSS.n2177 5.2005
R7844 VSS.n2180 VSS.n1070 5.2005
R7845 VSS.n2579 VSS.n2578 5.2005
R7846 VSS.n2576 VSS.n2575 5.2005
R7847 VSS.n2582 VSS.n2574 5.2005
R7848 VSS.n2586 VSS.n2585 5.2005
R7849 VSS.n1422 VSS.n1357 5.2005
R7850 VSS.n1453 VSS.n1328 5.2005
R7851 VSS.n1449 VSS.n1329 5.2005
R7852 VSS.n1447 VSS.n1446 5.2005
R7853 VSS.n1944 VSS.n1122 5.2005
R7854 VSS.n1942 VSS.n1940 5.2005
R7855 VSS.n1425 VSS.n1424 5.2005
R7856 VSS.n1429 VSS.n1428 5.2005
R7857 VSS.n1920 VSS.n1919 5.2005
R7858 VSS.n1926 VSS.n1925 5.2005
R7859 VSS.n1918 VSS.n1917 5.2005
R7860 VSS.n1912 VSS.n1911 5.2005
R7861 VSS.n1889 VSS.n1233 5.2005
R7862 VSS.n1897 VSS.n1896 5.2005
R7863 VSS.n1231 VSS.n1230 5.2005
R7864 VSS.n1231 VSS.n1228 5.2005
R7865 VSS.n1231 VSS.n1226 5.2005
R7866 VSS.n1231 VSS.n1224 5.2005
R7867 VSS.n1905 VSS.n1232 5.2005
R7868 VSS.n1346 VSS.n1231 5.2005
R7869 VSS.n1344 VSS.n1231 5.2005
R7870 VSS.n1342 VSS.n1231 5.2005
R7871 VSS.n1340 VSS.n1231 5.2005
R7872 VSS.n1332 VSS.n1331 5.2005
R7873 VSS.n1335 VSS.n1334 5.2005
R7874 VSS.n1338 VSS.n1337 5.2005
R7875 VSS.n1445 VSS.n1351 5.2005
R7876 VSS.n1939 VSS.n1938 5.2005
R7877 VSS.n1936 VSS.n1123 5.2005
R7878 VSS.n1932 VSS.n1124 5.2005
R7879 VSS.n1929 VSS.n1907 5.2005
R7880 VSS.n1771 VSS.n1770 5.2005
R7881 VSS.n1776 VSS.n1775 5.2005
R7882 VSS.n1712 VSS.n1711 5.2005
R7883 VSS.n1714 VSS.n1710 5.2005
R7884 VSS.n1706 VSS.n1705 5.2005
R7885 VSS.n1703 VSS.n1554 5.2005
R7886 VSS.n1701 VSS.n1700 5.2005
R7887 VSS.n1698 VSS.n1697 5.2005
R7888 VSS.n1691 VSS.n1690 5.2005
R7889 VSS.n1686 VSS.n1553 5.2005
R7890 VSS.n827 VSS.n826 5.2005
R7891 VSS.n831 VSS.n830 5.2005
R7892 VSS.n833 VSS.n832 5.2005
R7893 VSS.n837 VSS.n836 5.2005
R7894 VSS.n843 VSS.n842 5.2005
R7895 VSS.n847 VSS.n846 5.2005
R7896 VSS.n849 VSS.n848 5.2005
R7897 VSS.n853 VSS.n852 5.2005
R7898 VSS.n2650 VSS.n2649 5.2005
R7899 VSS.n1642 VSS.n1641 5.2005
R7900 VSS.n804 VSS.n803 5.2005
R7901 VSS.n799 VSS.n798 5.2005
R7902 VSS.n794 VSS.n793 5.2005
R7903 VSS.n1670 VSS.n1576 5.2005
R7904 VSS.n1674 VSS.n1673 5.2005
R7905 VSS.n1561 VSS.n1560 5.2005
R7906 VSS.n1594 VSS.n1592 5.2005
R7907 VSS.n1676 VSS.n1675 5.2005
R7908 VSS.n1679 VSS.n1564 5.2005
R7909 VSS.n1682 VSS.n1559 5.2005
R7910 VSS.n1685 VSS.n1557 5.2005
R7911 VSS.n2674 VSS.n792 5.2005
R7912 VSS.n2671 VSS.n797 5.2005
R7913 VSS.n2668 VSS.n802 5.2005
R7914 VSS.n2665 VSS.n807 5.2005
R7915 VSS.n2698 VSS.n2697 5.2005
R7916 VSS.n2695 VSS.n774 5.2005
R7917 VSS.n2693 VSS.n775 5.2005
R7918 VSS.n2691 VSS.n776 5.2005
R7919 VSS.n822 VSS.n821 5.2005
R7920 VSS.n1587 VSS.n1586 5.2005
R7921 VSS.n1587 VSS.n1584 5.2005
R7922 VSS.n1587 VSS.n1582 5.2005
R7923 VSS.n1587 VSS.n1580 5.2005
R7924 VSS.n1666 VSS.n1665 5.2005
R7925 VSS.n2678 VSS.n789 5.2005
R7926 VSS.n2681 VSS.n782 5.2005
R7927 VSS.n2684 VSS.n780 5.2005
R7928 VSS.n2686 VSS.n779 5.2005
R7929 VSS.n1630 VSS.n1629 5.2005
R7930 VSS.n784 VSS.n783 5.2005
R7931 VSS.n1568 VSS.n1566 5.2005
R7932 VSS.n1571 VSS.n1570 5.2005
R7933 VSS.n839 VSS.n838 5.2005
R7934 VSS.n1718 VSS.n1716 5.2005
R7935 VSS.n1720 VSS.n1708 5.2005
R7936 VSS.n1523 VSS.n1506 5.2005
R7937 VSS.n1240 VSS.n1239 5.2005
R7938 VSS.n1872 VSS.n1871 5.2005
R7939 VSS.n1876 VSS.n1875 5.2005
R7940 VSS.n1878 VSS.n1877 5.2005
R7941 VSS.n1882 VSS.n1881 5.2005
R7942 VSS.n1850 VSS.n1849 5.2005
R7943 VSS.n1467 VSS.n1466 5.2005
R7944 VSS.n1864 VSS.n1863 5.2005
R7945 VSS.n1529 VSS.n1528 5.2005
R7946 VSS.n1535 VSS.n1534 5.2005
R7947 VSS.n1537 VSS.n1536 5.2005
R7948 VSS.n1543 VSS.n1542 5.2005
R7949 VSS.n1753 VSS.n1752 5.2005
R7950 VSS.n1756 VSS.n1755 5.2005
R7951 VSS.n1759 VSS.n1758 5.2005
R7952 VSS.n1764 VSS.n1763 5.2005
R7953 VSS.n1747 VSS.n1746 5.2005
R7954 VSS.n1844 VSS.n1486 5.2005
R7955 VSS.n1843 VSS.n1842 5.2005
R7956 VSS.n1840 VSS.n1490 5.2005
R7957 VSS.n1838 VSS.n1837 5.2005
R7958 VSS.n1834 VSS.n1495 5.2005
R7959 VSS.n1858 VSS.n1857 5.2005
R7960 VSS.n1855 VSS.n1854 5.2005
R7961 VSS.n1852 VSS.n1851 5.2005
R7962 VSS.n1868 VSS.n1867 5.2005
R7963 VSS.n1462 VSS.n1243 5.2005
R7964 VSS.n1461 VSS.n1460 5.2005
R7965 VSS.n1458 VSS.n1245 5.2005
R7966 VSS.n1456 VSS.n1246 5.2005
R7967 VSS.n1323 VSS.n1322 5.2005
R7968 VSS.n1955 VSS.n1954 5.2005
R7969 VSS.n1952 VSS.n1118 5.2005
R7970 VSS.n1950 VSS.n1119 5.2005
R7971 VSS.n1948 VSS.n1120 5.2005
R7972 VSS.n1353 VSS.n1352 5.2005
R7973 VSS.n1440 VSS.n1439 5.2005
R7974 VSS.n1437 VSS.n1354 5.2005
R7975 VSS.n1435 VSS.n1355 5.2005
R7976 VSS.n1433 VSS.n1356 5.2005
R7977 VSS.n1381 VSS.n1379 5.2005
R7978 VSS.n1382 VSS.n1376 5.2005
R7979 VSS.n1383 VSS.n1373 5.2005
R7980 VSS.n1384 VSS.n1370 5.2005
R7981 VSS.n1385 VSS.n1367 5.2005
R7982 VSS.n2328 VSS.n2327 5.2005
R7983 VSS.n2329 VSS.n2324 5.2005
R7984 VSS.n2330 VSS.n2321 5.2005
R7985 VSS.n2331 VSS.n2318 5.2005
R7986 VSS.n2333 VSS.n2332 5.2005
R7987 VSS.n1963 VSS.n1962 5.2005
R7988 VSS.n1965 VSS.n1115 5.2005
R7989 VSS.n1967 VSS.n1113 5.2005
R7990 VSS.n1969 VSS.n1111 5.2005
R7991 VSS.n2234 VSS.n2233 5.2005
R7992 VSS.n2239 VSS.n2238 5.2005
R7993 VSS.n2241 VSS.n2230 5.2005
R7994 VSS.n2243 VSS.n2228 5.2005
R7995 VSS.n2245 VSS.n2226 5.2005
R7996 VSS.n2258 VSS.n2257 5.2005
R7997 VSS.n2269 VSS.n2268 5.2005
R7998 VSS.n2272 VSS.n2271 5.2005
R7999 VSS.n2287 VSS.n1106 5.2005
R8000 VSS.n2285 VSS.n1107 5.2005
R8001 VSS.n2283 VSS.n2282 5.2005
R8002 VSS.n2311 VSS.n2310 5.2005
R8003 VSS.n2343 VSS.n2342 5.2005
R8004 VSS.n2346 VSS.n2345 5.2005
R8005 VSS.n2357 VSS.n2356 5.2005
R8006 VSS.n2360 VSS.n2359 5.2005
R8007 VSS.n2381 VSS.n1074 5.2005
R8008 VSS.n2379 VSS.n1075 5.2005
R8009 VSS.n2377 VSS.n2376 5.2005
R8010 VSS.n2405 VSS.n2404 5.2005
R8011 VSS.n2260 VSS.n2259 5.2005
R8012 VSS.n2267 VSS.n2266 5.2005
R8013 VSS.n2264 VSS.n2263 5.2005
R8014 VSS.n2274 VSS.n2273 5.2005
R8015 VSS.n2278 VSS.n2277 5.2005
R8016 VSS.n2281 VSS.n2280 5.2005
R8017 VSS.n2313 VSS.n2312 5.2005
R8018 VSS.n2339 VSS.n2338 5.2005
R8019 VSS.n2348 VSS.n2347 5.2005
R8020 VSS.n2355 VSS.n2354 5.2005
R8021 VSS.n2352 VSS.n2351 5.2005
R8022 VSS.n2362 VSS.n2361 5.2005
R8023 VSS.n2366 VSS.n2365 5.2005
R8024 VSS.n2375 VSS.n2374 5.2005
R8025 VSS.n2372 VSS.n2369 5.2005
R8026 VSS.n1095 VSS.n1094 5.2005
R8027 VSS.n1097 VSS.n1096 5.2005
R8028 VSS.n1101 VSS.n1100 5.2005
R8029 VSS.n1103 VSS.n1102 5.2005
R8030 VSS.n2291 VSS.n2290 5.2005
R8031 VSS.n2296 VSS.n2295 5.2005
R8032 VSS.n2298 VSS.n2297 5.2005
R8033 VSS.n2301 VSS.n2300 5.2005
R8034 VSS.n2304 VSS.n2303 5.2005
R8035 VSS.n2306 VSS.n2305 5.2005
R8036 VSS.n2058 VSS.n2048 5.2005
R8037 VSS.n2057 VSS.n2056 5.2005
R8038 VSS.n2054 VSS.n2050 5.2005
R8039 VSS.n2052 VSS.n2051 5.2005
R8040 VSS.n2385 VSS.n2384 5.2005
R8041 VSS.n2390 VSS.n2389 5.2005
R8042 VSS.n2392 VSS.n2391 5.2005
R8043 VSS.n2395 VSS.n2394 5.2005
R8044 VSS.n2399 VSS.n2398 5.2005
R8045 VSS.n2140 VSS.n2138 5.2005
R8046 VSS.n2141 VSS.n2135 5.2005
R8047 VSS.n2142 VSS.n2132 5.2005
R8048 VSS.n2143 VSS.n2129 5.2005
R8049 VSS.n2144 VSS.n2126 5.2005
R8050 VSS.n2095 VSS.n2094 5.2005
R8051 VSS.n2096 VSS.n2091 5.2005
R8052 VSS.n2097 VSS.n2088 5.2005
R8053 VSS.n2098 VSS.n2085 5.2005
R8054 VSS.n2099 VSS.n2082 5.2005
R8055 VSS.n2079 VSS.n2078 5.2005
R8056 VSS.n2076 VSS.n2075 5.2005
R8057 VSS.n2074 VSS.n2073 5.2005
R8058 VSS.n2071 VSS.n2070 5.2005
R8059 VSS.n2036 VSS.n2035 5.2005
R8060 VSS.n2016 VSS.n2015 5.2005
R8061 VSS.n2018 VSS.n2012 5.2005
R8062 VSS.n2020 VSS.n2010 5.2005
R8063 VSS.n2022 VSS.n2008 5.2005
R8064 VSS.n2216 VSS.n2025 5.2005
R8065 VSS.n2214 VSS.n2027 5.2005
R8066 VSS.n2212 VSS.n2029 5.2005
R8067 VSS.n2210 VSS.n2031 5.2005
R8068 VSS.n2207 VSS.n2039 5.2005
R8069 VSS.n2205 VSS.n2041 5.2005
R8070 VSS.n2203 VSS.n2043 5.2005
R8071 VSS.n2201 VSS.n2045 5.2005
R8072 VSS.n2198 VSS.n2102 5.2005
R8073 VSS.n2196 VSS.n2104 5.2005
R8074 VSS.n2194 VSS.n2106 5.2005
R8075 VSS.n2192 VSS.n2108 5.2005
R8076 VSS.n2189 VSS.n2111 5.2005
R8077 VSS.n2187 VSS.n2113 5.2005
R8078 VSS.n2185 VSS.n2115 5.2005
R8079 VSS.n2183 VSS.n2117 5.2005
R8080 VSS.n2220 VSS.n2219 5.2005
R8081 VSS.n2255 VSS.n2254 5.2005
R8082 VSS.n2251 VSS.n2250 5.2005
R8083 VSS.n1846 VSS.n1485 5.2005
R8084 VSS.n1738 VSS.n1737 5.2005
R8085 VSS.n1740 VSS.n1739 5.2005
R8086 VSS.n1743 VSS.n1742 5.2005
R8087 VSS.n1598 VSS.n1597 5.2005
R8088 VSS.n1604 VSS.n1603 5.2005
R8089 VSS.n1602 VSS.n1601 5.2005
R8090 VSS.n1606 VSS.n1589 5.2005
R8091 VSS.n1614 VSS.n1613 5.2005
R8092 VSS.n1615 VSS.n1614 5.2005
R8093 VSS.n1618 VSS.n1617 5.2005
R8094 VSS.n1650 VSS.n1649 5.2005
R8095 VSS.n1651 VSS.n1639 5.2005
R8096 VSS.n1652 VSS.n1637 5.2005
R8097 VSS.n1653 VSS.n1635 5.2005
R8098 VSS.n1646 VSS.n1645 5.2005
R8099 VSS.n1657 VSS.n1627 5.2005
R8100 VSS.n1658 VSS.n1625 5.2005
R8101 VSS.n1659 VSS.n1623 5.2005
R8102 VSS.n1660 VSS.n1621 5.2005
R8103 VSS.n1656 VSS.n1634 5.2005
R8104 VSS.n2640 VSS.n2639 5.2005
R8105 VSS.n2638 VSS.n2637 5.2005
R8106 VSS.n2634 VSS.n2633 5.2005
R8107 VSS.n2632 VSS.n2631 5.2005
R8108 VSS.n2656 VSS.n813 5.2005
R8109 VSS.n2659 VSS.n811 5.2005
R8110 VSS.n2661 VSS.n810 5.2005
R8111 VSS.n2646 VSS.n2645 5.2005
R8112 VSS.n2643 VSS.n2642 5.2005
R8113 VSS.n817 VSS.n815 5.2005
R8114 VSS.n820 VSS.n819 5.2005
R8115 VSS.n881 VSS.n880 5.2005
R8116 VSS.n883 VSS.n882 5.2005
R8117 VSS.n887 VSS.n886 5.2005
R8118 VSS.n889 VSS.n888 5.2005
R8119 VSS.n1779 VSS.n1778 5.2005
R8120 VSS.n1782 VSS.n1781 5.2005
R8121 VSS.n1796 VSS.n1785 5.2005
R8122 VSS.n1794 VSS.n1787 5.2005
R8123 VSS.n1792 VSS.n1789 5.2005
R8124 VSS.n2596 VSS.n911 5.2005
R8125 VSS.n1826 VSS.n1507 5.2005
R8126 VSS.n1825 VSS.n1824 5.2005
R8127 VSS.n1822 VSS.n1511 5.2005
R8128 VSS.n1820 VSS.n1819 5.2005
R8129 VSS.n1815 VSS.n1801 5.2005
R8130 VSS.n1814 VSS.n1804 5.2005
R8131 VSS.n1813 VSS.n1807 5.2005
R8132 VSS.n1812 VSS.n1810 5.2005
R8133 VSS.n1816 VSS.n1514 5.2005
R8134 VSS.n2927 VSS.n2926 5.2005
R8135 VSS.n2925 VSS.n2924 5.2005
R8136 VSS.n949 VSS.n948 5.2005
R8137 VSS.n951 VSS.n917 5.2005
R8138 VSS.n953 VSS.n916 5.2005
R8139 VSS.n955 VSS.n915 5.2005
R8140 VSS.n921 VSS.n920 5.2005
R8141 VSS.n923 VSS.n922 5.2005
R8142 VSS.n926 VSS.n925 5.2005
R8143 VSS.n930 VSS.n929 5.2005
R8144 VSS.n932 VSS.n931 5.2005
R8145 VSS.n944 VSS.n933 5.2005
R8146 VSS.n943 VSS.n935 5.2005
R8147 VSS.n942 VSS.n937 5.2005
R8148 VSS.n941 VSS.n940 5.2005
R8149 VSS.n1174 VSS.n1173 5.2005
R8150 VSS.n2934 VSS.n2933 5.2005
R8151 VSS.n2930 VSS.n2929 5.2005
R8152 VSS.n893 VSS.n892 5.2005
R8153 VSS.n895 VSS.n894 5.2005
R8154 VSS.n2804 VSS.n2803 5.2005
R8155 VSS.n876 VSS.n875 5.2005
R8156 VSS.n901 VSS.n900 5.2005
R8157 VSS.n488 VSS.n487 5.2005
R8158 VSS.n489 VSS.n484 5.2005
R8159 VSS.n490 VSS.n481 5.2005
R8160 VSS.n491 VSS.n478 5.2005
R8161 VSS.n492 VSS.n474 5.2005
R8162 VSS.n471 VSS.n470 5.2005
R8163 VSS.n468 VSS.n467 5.2005
R8164 VSS.n466 VSS.n465 5.2005
R8165 VSS.n463 VSS.n462 5.2005
R8166 VSS.n461 VSS.n460 5.2005
R8167 VSS.n456 VSS.n455 5.2005
R8168 VSS.n453 VSS.n452 5.2005
R8169 VSS.n450 VSS.n449 5.2005
R8170 VSS.n448 VSS.n447 5.2005
R8171 VSS.n444 VSS.n443 5.2005
R8172 VSS.n437 VSS.n436 5.2005
R8173 VSS.n434 VSS.n433 5.2005
R8174 VSS.n432 VSS.n431 5.2005
R8175 VSS.n429 VSS.n428 5.2005
R8176 VSS.n427 VSS.n426 5.2005
R8177 VSS.n727 VSS.n361 5.2005
R8178 VSS.n731 VSS.n358 5.2005
R8179 VSS.n735 VSS.n355 5.2005
R8180 VSS.n739 VSS.n352 5.2005
R8181 VSS.n721 VSS.n366 5.2005
R8182 VSS.n717 VSS.n369 5.2005
R8183 VSS.n713 VSS.n371 5.2005
R8184 VSS.n709 VSS.n374 5.2005
R8185 VSS.n706 VSS.n376 5.2005
R8186 VSS.n710 VSS.n373 5.2005
R8187 VSS.n718 VSS.n368 5.2005
R8188 VSS.n722 VSS.n365 5.2005
R8189 VSS.n726 VSS.n362 5.2005
R8190 VSS.n730 VSS.n359 5.2005
R8191 VSS.n736 VSS.n354 5.2005
R8192 VSS.n740 VSS.n351 5.2005
R8193 VSS.n331 VSS.n330 5.2005
R8194 VSS.n1 VSS.n0 5.2005
R8195 VSS.n771 VSS.n770 5.15718
R8196 VSS.n763 VSS.n762 5.15718
R8197 VSS.n2793 VSS.n2792 5.15281
R8198 VSS.n761 VSS.n760 5.15281
R8199 VSS.n688 VSS.t1816 5.03731
R8200 VSS.n3119 VSS.n3118 4.93566
R8201 VSS.n1907 VSS.n1906 4.90616
R8202 VSS.n1665 VSS.n1664 4.61862
R8203 VSS.n870 VSS.n869 4.5005
R8204 VSS.n627 VSS.n626 4.5005
R8205 VSS.n3490 VSS.n3489 4.5005
R8206 VSS.n3489 VSS.n3488 4.5005
R8207 VSS.n3441 VSS.n3440 4.47093
R8208 VSS.n3449 VSS.n3448 4.3559
R8209 VSS.n1357 VSS.t2537 4.31466
R8210 VSS.n525 VSS.n512 4.30229
R8211 VSS VSS.n870 4.12455
R8212 VSS.n627 VSS 4.12355
R8213 VSS.n1846 VSS.n1845 4.08444
R8214 VSS.n2571 VSS.n2570 3.83432
R8215 VSS.n3422 VSS.n32 3.82133
R8216 VSS.n1416 VSS.t1910 3.81142
R8217 VSS.n1978 VSS.t1949 3.81141
R8218 VSS.n1252 VSS.t1831 3.81141
R8219 VSS.n2176 VSS.t1821 3.81141
R8220 VSS.n1596 VSS.t2106 3.81141
R8221 VSS.t1207 VSS.t1211 3.68113
R8222 VSS.n1130 VSS.t537 3.68113
R8223 VSS.t2447 VSS.t2436 3.68113
R8224 VSS.t759 VSS.n1187 3.68113
R8225 VSS.t2441 VSS.t2439 3.68113
R8226 VSS.t1198 VSS.t1201 3.68113
R8227 VSS.t1209 VSS.t1213 3.68113
R8228 VSS.n1159 VSS.t1186 3.68113
R8229 VSS.t2445 VSS.t2442 3.68113
R8230 VSS.t1276 VSS.n1139 3.68113
R8231 VSS.t2443 VSS.t1163 3.68113
R8232 VSS.t1497 VSS.t918 3.67489
R8233 VSS.n1700 VSS.n1554 3.67489
R8234 VSS.t2297 VSS.t767 3.67489
R8235 VSS.n3488 VSS.n5 3.67489
R8236 VSS.n2763 VSS.n2762 3.56644
R8237 VSS.n1149 VSS.n1141 3.37613
R8238 VSS.n1157 VSS.n1140 3.37613
R8239 VSS.n1166 VSS.n1164 3.37613
R8240 VSS.n1180 VSS.n1170 3.37613
R8241 VSS.n1196 VSS.n1127 3.37613
R8242 VSS.n1189 VSS.n1132 3.37613
R8243 VSS.n1185 VSS.n1135 3.37613
R8244 VSS.n1828 VSS.n1827 3.36838
R8245 VSS.n3260 VSS.n222 3.36453
R8246 VSS.n2005 VSS.n1977 3.36323
R8247 VSS.n1279 VSS.n1251 3.36323
R8248 VSS.n2416 VSS.n1066 3.36323
R8249 VSS.n1419 VSS.n1359 3.36323
R8250 VSS.n2179 VSS.n2119 3.36323
R8251 VSS.n1595 VSS.n1591 3.36323
R8252 VSS.n1689 VSS.n1556 3.28959
R8253 VSS.n335 VSS.n334 3.28959
R8254 VSS.n2252 VSS.n2251 3.27176
R8255 VSS VSS.n957 3.25698
R8256 VSS.n1762 VSS.n1761 3.20563
R8257 VSS.n2408 VSS.n957 3.2003
R8258 VSS.n2921 VSS.n2920 3.1685
R8259 VSS.n2411 VSS.n2408 3.07634
R8260 VSS.n1699 VSS.n1698 3.03722
R8261 VSS.n241 VSS.t1626 3.0114
R8262 VSS.n3073 VSS 2.96937
R8263 VSS.n2510 VSS.t2524 2.94368
R8264 VSS.n129 VSS 2.84263
R8265 VSS.t1690 VSS.n3140 2.73236
R8266 VSS.n3141 VSS.t1004 2.73236
R8267 VSS.n3255 VSS.n3254 2.6035
R8268 VSS.n3239 VSS.n3238 2.6035
R8269 VSS.n3247 VSS.n3246 2.6035
R8270 VSS VSS.n1144 2.6035
R8271 VSS.n1197 VSS 2.6035
R8272 VSS.n1186 VSS 2.6035
R8273 VSS VSS.n1131 2.6035
R8274 VSS VSS.n1152 2.6035
R8275 VSS.n1169 VSS 2.6035
R8276 VSS VSS.n1160 2.6035
R8277 VSS VSS.n3232 2.60126
R8278 VSS.n2603 VSS.n2602 2.6005
R8279 VSS.n2602 VSS.n2601 2.6005
R8280 VSS.n3236 VSS.n3235 2.6005
R8281 VSS.t610 VSS.n3236 2.6005
R8282 VSS.n3232 VSS.n3231 2.6005
R8283 VSS.n632 VSS.n631 2.6005
R8284 VSS.n633 VSS.n632 2.6005
R8285 VSS.n1185 VSS.n1184 2.6005
R8286 VSS.t2439 VSS.n1185 2.6005
R8287 VSS.n1191 VSS.n1132 2.6005
R8288 VSS.n1132 VSS.t2447 2.6005
R8289 VSS.n1196 VSS.n1195 2.6005
R8290 VSS.t1211 VSS.n1196 2.6005
R8291 VSS VSS.n1135 2.6005
R8292 VSS.n1135 VSS.n1134 2.6005
R8293 VSS VSS.n1189 2.6005
R8294 VSS.n1189 VSS.n1188 2.6005
R8295 VSS VSS.n1127 2.6005
R8296 VSS.n1129 VSS.n1127 2.6005
R8297 VSS VSS.n1180 2.6005
R8298 VSS.n1180 VSS.n1179 2.6005
R8299 VSS VSS.n1166 2.6005
R8300 VSS.n1166 VSS.n1165 2.6005
R8301 VSS.n1157 VSS 2.6005
R8302 VSS.n1158 VSS.n1157 2.6005
R8303 VSS.n1149 VSS 2.6005
R8304 VSS.n1150 VSS.n1149 2.6005
R8305 VSS.n1170 VSS.n1138 2.6005
R8306 VSS.n1170 VSS.t2443 2.6005
R8307 VSS.n1164 VSS.n1163 2.6005
R8308 VSS.n1164 VSS.t2445 2.6005
R8309 VSS.n1154 VSS.n1140 2.6005
R8310 VSS.t1213 VSS.n1140 2.6005
R8311 VSS.n1146 VSS.n1141 2.6005
R8312 VSS.t1201 VSS.n1141 2.6005
R8313 VSS.n769 VSS.n768 2.59576
R8314 VSS.n2789 VSS.n2788 2.59576
R8315 VSS.t1816 VSS.t1255 2.5189
R8316 VSS.n3488 VSS.n4 2.4849
R8317 VSS VSS.n2005 2.40845
R8318 VSS VSS.n1279 2.40845
R8319 VSS.n1595 VSS 2.40845
R8320 VSS.n875 VSS.t899 2.40257
R8321 VSS.n2807 VSS.t1301 2.40257
R8322 VSS.n3389 VSS.n3388 2.38977
R8323 VSS.n1906 VSS.n1905 2.38977
R8324 VSS VSS.n2572 2.38278
R8325 VSS.n2570 VSS.n2569 2.2505
R8326 VSS.n2920 VSS.n755 2.2505
R8327 VSS.n2918 VSS.n2915 2.24865
R8328 VSS.n2918 VSS.n2835 2.24839
R8329 VSS VSS.n108 2.24014
R8330 VSS.n716 VSS 2.24014
R8331 VSS.n1765 VSS 2.24014
R8332 VSS.n1928 VSS.n1927 2.2128
R8333 VSS.t2334 VSS.t1641 2.19348
R8334 VSS.t1397 VSS.t852 2.19348
R8335 VSS.n1888 VSS 2.14127
R8336 VSS.n3491 VSS.n3490 2.13837
R8337 VSS.n1693 VSS.n1692 2.13725
R8338 VSS.n1420 VSS 2.1304
R8339 VSS VSS.n2182 2.1304
R8340 VSS.n3446 VSS 2.0829
R8341 VSS.n1688 VSS 2.03762
R8342 VSS.n1421 VSS 1.99132
R8343 VSS VSS.n2181 1.99132
R8344 VSS.n3172 VSS 1.98504
R8345 VSS.n3032 VSS.t451 1.97859
R8346 VSS.n3408 VSS 1.92724
R8347 VSS.n1927 VSS.n956 1.85846
R8348 VSS.n2569 VSS.n958 1.71863
R8349 VSS.n1178 VSS.n1177 1.69233
R8350 VSS.n3209 VSS.n237 1.56287
R8351 VSS.n2920 VSS.n2919 1.53562
R8352 VSS.n754 VSS.n336 1.46066
R8353 VSS.n2415 VSS.n2411 1.4385
R8354 VSS.n2415 VSS.n2414 1.37944
R8355 VSS.n1733 VSS.n1732 1.36907
R8356 VSS.n2798 VSS.n2797 1.30375
R8357 VSS.n2800 VSS.n2799 1.30375
R8358 VSS.n2802 VSS.n2801 1.30375
R8359 VSS.n757 VSS.n756 1.30375
R8360 VSS.n2809 VSS.n2808 1.30375
R8361 VSS.n2812 VSS.n2811 1.30375
R8362 VSS.n2816 VSS.n2815 1.30375
R8363 VSS.n2913 VSS.n2838 1.3005
R8364 VSS.n2912 VSS.n2839 1.3005
R8365 VSS.n2911 VSS.n2840 1.3005
R8366 VSS.n2910 VSS.n2841 1.3005
R8367 VSS.n2909 VSS.n2842 1.3005
R8368 VSS.n2908 VSS.n2843 1.3005
R8369 VSS.n2907 VSS.n2844 1.3005
R8370 VSS.n2906 VSS.n2849 1.3005
R8371 VSS.n2905 VSS.n2850 1.3005
R8372 VSS.n2904 VSS.n2851 1.3005
R8373 VSS.n2903 VSS.n2852 1.3005
R8374 VSS.n2902 VSS.n2853 1.3005
R8375 VSS.n2901 VSS.n2854 1.3005
R8376 VSS.n2900 VSS.n2855 1.3005
R8377 VSS.n2899 VSS.n2856 1.3005
R8378 VSS.n2898 VSS.n2857 1.3005
R8379 VSS.n2897 VSS.n2858 1.3005
R8380 VSS.n2896 VSS.n2859 1.3005
R8381 VSS.n2895 VSS.n2860 1.3005
R8382 VSS.n2894 VSS.n2861 1.3005
R8383 VSS.n2893 VSS.n2862 1.3005
R8384 VSS.n2892 VSS.n2863 1.3005
R8385 VSS.n2891 VSS.n2864 1.3005
R8386 VSS.n2890 VSS.n2865 1.3005
R8387 VSS.n2889 VSS.n2866 1.3005
R8388 VSS.n2888 VSS.n2867 1.3005
R8389 VSS.n2887 VSS.n2868 1.3005
R8390 VSS.n2886 VSS.n2869 1.3005
R8391 VSS.n2885 VSS.n2870 1.3005
R8392 VSS.n2884 VSS.n2871 1.3005
R8393 VSS.n2883 VSS.n2872 1.3005
R8394 VSS.n2882 VSS.n2873 1.3005
R8395 VSS.n2881 VSS.n2874 1.3005
R8396 VSS.n2880 VSS.n2875 1.3005
R8397 VSS.n2879 VSS.n2876 1.3005
R8398 VSS.n2704 VSS.n2703 1.3005
R8399 VSS.n2706 VSS.n2705 1.3005
R8400 VSS.n2709 VSS.n2708 1.3005
R8401 VSS.n2711 VSS.n2710 1.3005
R8402 VSS.n2713 VSS.n2712 1.3005
R8403 VSS.n2715 VSS.n2714 1.3005
R8404 VSS.n2717 VSS.n2716 1.3005
R8405 VSS.n2719 VSS.n2718 1.3005
R8406 VSS.n2721 VSS.n2720 1.3005
R8407 VSS.n2723 VSS.n2722 1.3005
R8408 VSS.n2725 VSS.n2724 1.3005
R8409 VSS.n2727 VSS.n2726 1.3005
R8410 VSS.n2729 VSS.n2728 1.3005
R8411 VSS.n2732 VSS.n2731 1.3005
R8412 VSS.n2734 VSS.n2733 1.3005
R8413 VSS.n2736 VSS.n2735 1.3005
R8414 VSS.n2738 VSS.n2737 1.3005
R8415 VSS.n2741 VSS.n2740 1.3005
R8416 VSS.n2743 VSS.n2742 1.3005
R8417 VSS.n2745 VSS.n2744 1.3005
R8418 VSS.n2747 VSS.n2746 1.3005
R8419 VSS.n2749 VSS.n2748 1.3005
R8420 VSS.n2751 VSS.n2750 1.3005
R8421 VSS.n2753 VSS.n2752 1.3005
R8422 VSS.n2755 VSS.n2754 1.3005
R8423 VSS.n2757 VSS.n2756 1.3005
R8424 VSS.n2759 VSS.n2758 1.3005
R8425 VSS.n2761 VSS.n2760 1.3005
R8426 VSS.n2764 VSS.n2763 1.3005
R8427 VSS.n2766 VSS.n2765 1.3005
R8428 VSS.n2768 VSS.n2767 1.3005
R8429 VSS.n2770 VSS.n2769 1.3005
R8430 VSS.n2772 VSS.n2771 1.3005
R8431 VSS.n2774 VSS.n2773 1.3005
R8432 VSS.n2776 VSS.n2775 1.3005
R8433 VSS.n2778 VSS.n2777 1.3005
R8434 VSS.n2780 VSS.n2779 1.3005
R8435 VSS.n2784 VSS.n2783 1.3005
R8436 VSS.n2818 VSS.n2817 1.3005
R8437 VSS.n2820 VSS.n2819 1.3005
R8438 VSS.n2822 VSS.n2821 1.3005
R8439 VSS.n2824 VSS.n2823 1.3005
R8440 VSS.n2826 VSS.n2825 1.3005
R8441 VSS.n2828 VSS.n2827 1.3005
R8442 VSS.n2832 VSS.n2831 1.12018
R8443 VSS.n2837 VSS.n2836 1.12018
R8444 VSS.n1761 VSS.t529 1.09297
R8445 VSS.n2609 VSS 1.09141
R8446 VSS VSS.n616 1.09141
R8447 VSS.n2648 VSS.n2647 1.03389
R8448 VSS.n1931 VSS.n1930 1.03389
R8449 VSS.n1431 VSS.n1430 1.03335
R8450 VSS.n2249 VSS.n2248 1.03307
R8451 VSS.n2218 VSS.n2217 1.03307
R8452 VSS.n1700 VSS.n1699 1.00481
R8453 VSS.n1177 VSS.n1171 0.944719
R8454 VSS.n3425 VSS.n3424 0.943665
R8455 VSS.n3265 VSS.n3260 0.919774
R8456 VSS.n2507 VSS.n2506 0.918836
R8457 VSS.n3412 VSS.n3411 0.917851
R8458 VSS.n130 VSS.n129 0.899322
R8459 VSS.n3455 VSS.n3454 0.850616
R8460 VSS.n3394 VSS.n79 0.846463
R8461 VSS.n3381 VSS.n3380 0.846463
R8462 VSS.n3354 VSS.n113 0.846463
R8463 VSS.n714 VSS.n370 0.846463
R8464 VSS.n476 VSS.n384 0.846463
R8465 VSS.n733 VSS.n356 0.846463
R8466 VSS.n425 VSS.n424 0.846463
R8467 VSS.n2363 VSS.n1078 0.846463
R8468 VSS.n2337 VSS.n2334 0.846463
R8469 VSS.n2275 VSS.n1971 0.846463
R8470 VSS.n2191 VSS.n2109 0.846463
R8471 VSS.n2200 VSS.n2046 0.846463
R8472 VSS.n2209 VSS.n2032 0.846463
R8473 VSS.n1349 VSS.n1348 0.846463
R8474 VSS.n1647 VSS.n1644 0.846463
R8475 VSS.n1633 VSS.n1632 0.846463
R8476 VSS.n1668 VSS.n1667 0.846463
R8477 VSS.n1733 VSS.n1730 0.845914
R8478 VSS.n1748 VSS.n1550 0.845914
R8479 VSS.n2289 VSS.n2288 0.845914
R8480 VSS.n2308 VSS.n2307 0.845914
R8481 VSS.n2383 VSS.n2382 0.845914
R8482 VSS.n1305 VSS.n1291 0.845914
R8483 VSS.n1454 VSS.n1324 0.845914
R8484 VSS.n1946 VSS.n1945 0.845914
R8485 VSS.n3048 VSS.n3047 0.845914
R8486 VSS.n3201 VSS.n243 0.845914
R8487 VSS.n2460 VSS.n2459 0.845914
R8488 VSS.n3185 VSS.n254 0.845914
R8489 VSS.n2530 VSS.n969 0.845914
R8490 VSS.n2922 VSS.n327 0.845914
R8491 VSS.n3061 VSS.n3060 0.845914
R8492 VSS.n2407 VSS.n1067 0.845914
R8493 VSS.n1766 VSS.n1524 0.845914
R8494 VSS.n1799 VSS.n1798 0.845914
R8495 VSS.n3438 VSS.n3437 0.844811
R8496 VSS.n742 VSS.n349 0.843955
R8497 VSS.n2689 VSS.n2688 0.843955
R8498 VSS.n2570 VSS.n957 0.828588
R8499 VSS.n3172 VSS.n3171 0.825821
R8500 VSS.n1866 VSS.n1865 0.819492
R8501 VSS.n1887 VSS.n1236 0.817015
R8502 VSS.n2560 VSS.n965 0.807932
R8503 VSS.n3151 VSS.n3150 0.807932
R8504 VSS.n903 VSS.n902 0.796031
R8505 VSS.n2675 VSS.n791 0.73944
R8506 VSS.n676 VSS.n497 0.734346
R8507 VSS.n901 VSS.n899 0.734346
R8508 VSS.n3120 VSS.n3119 0.729114
R8509 VSS.n724 VSS.n363 0.70444
R8510 VSS.n3160 VSS.n279 0.692427
R8511 VSS.n3484 VSS 0.676801
R8512 VSS VSS.n1704 0.676801
R8513 VSS.n898 VSS.n896 0.645242
R8514 VSS.n2936 VSS.n325 0.637841
R8515 VSS.n691 VSS.n690 0.623774
R8516 VSS.n1688 VSS.n1687 0.616742
R8517 VSS.n336 VSS.n332 0.616742
R8518 VSS.n2662 VSS.n809 0.605183
R8519 VSS.n705 VSS.n377 0.574895
R8520 VSS.n2408 VSS.n2407 0.567839
R8521 VSS.n2416 VSS.n2415 0.534803
R8522 VSS VSS.n2337 0.520683
R8523 VSS.n2363 VSS 0.520683
R8524 VSS VSS.n2200 0.520683
R8525 VSS VSS.n2191 0.520683
R8526 VSS.n2288 VSS 0.519858
R8527 VSS.n2308 VSS 0.519858
R8528 VSS.n1291 VSS 0.519858
R8529 VSS.n1454 VSS 0.519858
R8530 VSS.n1698 VSS.n1694 0.486611
R8531 VSS.n2269 VSS.n1974 0.480225
R8532 VSS.n2271 VSS.n2270 0.480225
R8533 VSS.n2284 VSS.n2283 0.480225
R8534 VSS.n2310 VSS.n1088 0.480225
R8535 VSS.n2357 VSS.n1081 0.480225
R8536 VSS.n2359 VSS.n2358 0.480225
R8537 VSS.n1286 VSS.n1285 0.480225
R8538 VSS.n1289 VSS.n1249 0.480225
R8539 VSS.n1459 VSS.n1458 0.480225
R8540 VSS.n1457 VSS.n1456 0.480225
R8541 VSS.n1450 VSS.n1449 0.480225
R8542 VSS.n1448 VSS.n1447 0.480225
R8543 VSS.n2525 VSS.n2524 0.480225
R8544 VSS.n2528 VSS.n970 0.480225
R8545 VSS.n2538 VSS.n2537 0.480225
R8546 VSS.n2536 VSS.n2535 0.480225
R8547 VSS.n1429 VSS.n1423 0.480225
R8548 VSS.n2261 VSS.n2260 0.480225
R8549 VSS.n2266 VSS.n2265 0.480225
R8550 VSS.n2279 VSS.n2278 0.480225
R8551 VSS.n2280 VSS.n1087 0.480225
R8552 VSS.n2349 VSS.n2348 0.480225
R8553 VSS.n2354 VSS.n2353 0.480225
R8554 VSS.n2367 VSS.n2366 0.480225
R8555 VSS.n2374 VSS.n2373 0.480225
R8556 VSS.n2216 VSS.n2215 0.480225
R8557 VSS.n2214 VSS.n2213 0.480225
R8558 VSS.n2207 VSS.n2206 0.480225
R8559 VSS.n2205 VSS.n2204 0.480225
R8560 VSS.n2198 VSS.n2197 0.480225
R8561 VSS.n2196 VSS.n2195 0.480225
R8562 VSS.n2189 VSS.n2188 0.480225
R8563 VSS.n2187 VSS.n2186 0.480225
R8564 VSS.n1338 VSS.n1336 0.480225
R8565 VSS.n1351 VSS.n1339 0.480225
R8566 VSS.n1935 VSS.n1934 0.480225
R8567 VSS.n1933 VSS.n1932 0.480225
R8568 VSS.n2646 VSS.n2644 0.480225
R8569 VSS.n1865 VSS 0.473
R8570 VSS.n3480 VSS.n3479 0.439554
R8571 VSS.n1716 VSS.n1709 0.439554
R8572 VSS VSS.n790 0.43894
R8573 VSS VSS.n1888 0.438387
R8574 VSS.n754 VSS 0.432899
R8575 VSS.n1927 VSS 0.413056
R8576 VSS.n1392 VSS.n1389 0.396541
R8577 VSS.n1403 VSS.n1402 0.396541
R8578 VSS.n1398 VSS.n1397 0.396541
R8579 VSS.n2152 VSS.n2149 0.396541
R8580 VSS.n2163 VSS.n2162 0.396541
R8581 VSS.n2159 VSS.n2158 0.396541
R8582 VSS.n1989 VSS.n1988 0.396455
R8583 VSS.n1993 VSS.n1992 0.396455
R8584 VSS.n1997 VSS.n1996 0.396455
R8585 VSS.n1264 VSS.n1263 0.396455
R8586 VSS.n1268 VSS.n1267 0.396455
R8587 VSS.n1272 VSS.n1271 0.396455
R8588 VSS.n2437 VSS.n2436 0.396455
R8589 VSS.n2441 VSS.n2440 0.396455
R8590 VSS.n2431 VSS.n2429 0.396455
R8591 VSS.n1616 VSS.n1615 0.395692
R8592 VSS.n1613 VSS.n1611 0.395692
R8593 VSS.n1608 VSS.n1607 0.395692
R8594 VSS.n3408 VSS 0.392281
R8595 VSS.n2003 VSS 0.379596
R8596 VSS VSS.n1253 0.379596
R8597 VSS VSS.n2420 0.379596
R8598 VSS VSS.n1413 0.378121
R8599 VSS VSS.n2173 0.378121
R8600 VSS VSS.n1599 0.378121
R8601 VSS.n866 VSS.n865 0.365463
R8602 VSS.n607 VSS.n606 0.365463
R8603 VSS.n1855 VSS.n1853 0.363625
R8604 VSS.n1857 VSS.n1856 0.363625
R8605 VSS.n1468 VSS.n1467 0.363625
R8606 VSS.n1885 VSS.n1237 0.363625
R8607 VSS VSS.n1420 0.357797
R8608 VSS.n2182 VSS 0.357797
R8609 VSS.n1668 VSS.n778 0.35472
R8610 VSS.n2378 VSS.n2377 0.353977
R8611 VSS.n903 VSS.n755 0.348751
R8612 VSS.n1671 VSS.n1670 0.348115
R8613 VSS VSS.n1841 0.343161
R8614 VSS VSS.n1839 0.343161
R8615 VSS.n1479 VSS 0.343161
R8616 VSS.n1477 VSS 0.343161
R8617 VSS.n1501 VSS 0.343161
R8618 VSS.n1504 VSS 0.343161
R8619 VSS.n1229 VSS 0.343161
R8620 VSS.n1227 VSS 0.343161
R8621 VSS.n1093 VSS 0.343161
R8622 VSS VSS.n1098 0.343161
R8623 VSS.n2294 VSS 0.343161
R8624 VSS VSS.n2299 0.343161
R8625 VSS VSS.n2049 0.343161
R8626 VSS.n2055 VSS 0.343161
R8627 VSS VSS.n2256 0.343161
R8628 VSS.n2286 VSS 0.343161
R8629 VSS VSS.n2344 0.343161
R8630 VSS.n2380 VSS 0.343161
R8631 VSS.n1438 VSS 0.343161
R8632 VSS.n1436 VSS 0.343161
R8633 VSS.n1293 VSS 0.343161
R8634 VSS VSS.n1298 0.343161
R8635 VSS.n1310 VSS 0.343161
R8636 VSS VSS.n1315 0.343161
R8637 VSS.n1953 VSS 0.343161
R8638 VSS.n1951 VSS 0.343161
R8639 VSS.n1280 VSS 0.343161
R8640 VSS VSS.n1244 0.343161
R8641 VSS.n1452 VSS 0.343161
R8642 VSS.n1943 VSS 0.343161
R8643 VSS VSS.n3016 0.343161
R8644 VSS.n3053 VSS 0.343161
R8645 VSS VSS.n1007 0.343161
R8646 VSS.n1008 VSS 0.343161
R8647 VSS.n2446 VSS 0.343161
R8648 VSS VSS.n2451 0.343161
R8649 VSS.n2465 VSS 0.343161
R8650 VSS VSS.n2470 0.343161
R8651 VSS.n99 VSS 0.343161
R8652 VSS.n102 VSS 0.343161
R8653 VSS.n87 VSS 0.343161
R8654 VSS.n90 VSS 0.343161
R8655 VSS VSS.n3344 0.343161
R8656 VSS VSS.n3342 0.343161
R8657 VSS VSS.n120 0.343161
R8658 VSS.n3286 VSS 0.343161
R8659 VSS.n56 VSS 0.343161
R8660 VSS VSS.n61 0.343161
R8661 VSS VSS.n273 0.343161
R8662 VSS VSS.n271 0.343161
R8663 VSS VSS.n1032 0.343161
R8664 VSS VSS.n1034 0.343161
R8665 VSS.n2519 VSS 0.343161
R8666 VSS VSS.n2532 0.343161
R8667 VSS VSS.n1037 0.343161
R8668 VSS.n1043 VSS 0.343161
R8669 VSS VSS.n992 0.343161
R8670 VSS VSS.n990 0.343161
R8671 VSS VSS.n2479 0.343161
R8672 VSS VSS.n2481 0.343161
R8673 VSS.n919 VSS 0.343161
R8674 VSS VSS.n924 0.343161
R8675 VSS VSS.n934 0.343161
R8676 VSS VSS.n936 0.343161
R8677 VSS VSS.n1019 0.343161
R8678 VSS VSS.n1021 0.343161
R8679 VSS VSS.n3004 0.343161
R8680 VSS VSS.n3002 0.343161
R8681 VSS VSS.n43 0.343161
R8682 VSS VSS.n41 0.343161
R8683 VSS.n3462 VSS 0.343161
R8684 VSS.n3460 VSS 0.343161
R8685 VSS VSS.n389 0.343161
R8686 VSS.n469 VSS 0.343161
R8687 VSS.n483 VSS 0.343161
R8688 VSS.n486 VSS 0.343161
R8689 VSS.n451 VSS 0.343161
R8690 VSS.n454 VSS 0.343161
R8691 VSS VSS.n419 0.343161
R8692 VSS.n435 VSS 0.343161
R8693 VSS VSS.n2983 0.343161
R8694 VSS.n2984 VSS 0.343161
R8695 VSS.n2549 VSS 0.343161
R8696 VSS.n2547 VSS 0.343161
R8697 VSS.n1375 VSS 0.343161
R8698 VSS.n1378 VSS 0.343161
R8699 VSS.n2323 VSS 0.343161
R8700 VSS.n2326 VSS 0.343161
R8701 VSS VSS.n1966 0.343161
R8702 VSS VSS.n1964 0.343161
R8703 VSS VSS.n2242 0.343161
R8704 VSS VSS.n2240 0.343161
R8705 VSS VSS.n1973 0.343161
R8706 VSS.n2314 VSS 0.343161
R8707 VSS VSS.n1080 0.343161
R8708 VSS VSS.n2371 0.343161
R8709 VSS.n2134 VSS 0.343161
R8710 VSS.n2137 VSS 0.343161
R8711 VSS.n2090 VSS 0.343161
R8712 VSS.n2093 VSS 0.343161
R8713 VSS VSS.n2066 0.343161
R8714 VSS.n2077 VSS 0.343161
R8715 VSS VSS.n2019 0.343161
R8716 VSS VSS.n2017 0.343161
R8717 VSS VSS.n2211 0.343161
R8718 VSS VSS.n2202 0.343161
R8719 VSS VSS.n2193 0.343161
R8720 VSS VSS.n2184 0.343161
R8721 VSS.n2388 VSS 0.343161
R8722 VSS VSS.n2393 0.343161
R8723 VSS VSS.n1341 0.343161
R8724 VSS VSS.n1343 0.343161
R8725 VSS.n1330 VSS 0.343161
R8726 VSS.n1937 VSS 0.343161
R8727 VSS VSS.n1823 0.343161
R8728 VSS VSS.n1821 0.343161
R8729 VSS.n1806 VSS 0.343161
R8730 VSS.n1809 VSS 0.343161
R8731 VSS.n2630 VSS 0.343161
R8732 VSS VSS.n2635 0.343161
R8733 VSS VSS.n1636 0.343161
R8734 VSS VSS.n1638 0.343161
R8735 VSS VSS.n1622 0.343161
R8736 VSS VSS.n1624 0.343161
R8737 VSS VSS.n1581 0.343161
R8738 VSS VSS.n1583 0.343161
R8739 VSS.n1569 VSS 0.343161
R8740 VSS.n818 VSS 0.343161
R8741 VSS VSS.n1873 0.343161
R8742 VSS.n1874 VSS 0.343161
R8743 VSS.n891 VSS.n873 0.338437
R8744 VSS.n682 VSS.n681 0.338437
R8745 VSS.n2560 VSS 0.336214
R8746 VSS.n1673 VSS.n1563 0.325821
R8747 VSS.n755 VSS.n754 0.320599
R8748 VSS.n3482 VSS.n3481 0.316175
R8749 VSS.n1708 VSS.n1707 0.316175
R8750 VSS.n784 VSS.n781 0.313436
R8751 VSS.n3478 VSS 0.311851
R8752 VSS.n1715 VSS 0.311851
R8753 VSS.n1411 VSS 0.311509
R8754 VSS.n2171 VSS 0.311509
R8755 VSS.n2001 VSS 0.310668
R8756 VSS VSS.n1255 0.310668
R8757 VSS VSS.n2423 0.310668
R8758 VSS.n1600 VSS 0.310668
R8759 VSS.n3329 VSS.n3328 0.310174
R8760 VSS.n3311 VSS.n3310 0.310174
R8761 VSS.n647 VSS.n646 0.310174
R8762 VSS.n401 VSS.n400 0.310174
R8763 VSS.n1915 VSS.n1914 0.310174
R8764 VSS.n1532 VSS.n1531 0.310174
R8765 VSS.n2514 VSS.n2513 0.309418
R8766 VSS.n2581 VSS.n2580 0.309418
R8767 VSS.n1894 VSS.n1893 0.309418
R8768 VSS.n3176 VSS.n3175 0.308088
R8769 VSS.n3177 VSS.n71 0.308088
R8770 VSS.n1888 VSS.n1887 0.3055
R8771 VSS.n2643 VSS.n812 0.294445
R8772 VSS.n3437 VSS 0.290741
R8773 VSS VSS.n1486 0.289491
R8774 VSS VSS.n1474 0.289491
R8775 VSS VSS.n1496 0.289491
R8776 VSS VSS.n1224 0.289491
R8777 VSS.n1103 VSS 0.289491
R8778 VSS.n2303 VSS 0.289491
R8779 VSS VSS.n2052 0.289491
R8780 VSS VSS.n1433 0.289491
R8781 VSS.n1303 VSS 0.289491
R8782 VSS.n1319 VSS 0.289491
R8783 VSS VSS.n1948 0.289491
R8784 VSS VSS.n3050 0.289491
R8785 VSS.n1015 VSS 0.289491
R8786 VSS.n2456 VSS 0.289491
R8787 VSS.n2475 VSS 0.289491
R8788 VSS VSS.n94 0.289491
R8789 VSS VSS.n82 0.289491
R8790 VSS.n3347 VSS 0.289491
R8791 VSS VSS.n3280 0.289491
R8792 VSS.n66 VSS 0.289491
R8793 VSS VSS.n263 0.289491
R8794 VSS VSS.n1051 0.289491
R8795 VSS VSS.n1040 0.289491
R8796 VSS.n995 VSS 0.289491
R8797 VSS.n2484 VSS 0.289491
R8798 VSS.n929 VSS 0.289491
R8799 VSS.n940 VSS 0.289491
R8800 VSS VSS.n1024 0.289491
R8801 VSS VSS.n2994 0.289491
R8802 VSS.n46 VSS 0.289491
R8803 VSS VSS.n3457 0.289491
R8804 VSS VSS.n463 0.289491
R8805 VSS VSS.n478 0.289491
R8806 VSS.n447 VSS 0.289491
R8807 VSS VSS.n429 0.289491
R8808 VSS.n2990 VSS 0.289491
R8809 VSS.n3153 VSS 0.289491
R8810 VSS VSS.n1370 0.289491
R8811 VSS VSS.n2318 0.289491
R8812 VSS.n1969 VSS 0.289491
R8813 VSS.n2245 VSS 0.289491
R8814 VSS VSS.n2129 0.289491
R8815 VSS VSS.n2085 0.289491
R8816 VSS VSS.n2071 0.289491
R8817 VSS.n2022 VSS 0.289491
R8818 VSS.n2398 VSS 0.289491
R8819 VSS.n1346 VSS 0.289491
R8820 VSS VSS.n1507 0.289491
R8821 VSS VSS.n1801 0.289491
R8822 VSS.n2640 VSS 0.289491
R8823 VSS.n1649 VSS 0.289491
R8824 VSS.n1627 VSS 0.289491
R8825 VSS.n1586 VSS 0.289491
R8826 VSS.n1881 VSS 0.289491
R8827 VSS.n2657 VSS.n2656 0.286539
R8828 VSS.n661 VSS.n660 0.284276
R8829 VSS.n2806 VSS.n2805 0.284276
R8830 VSS.n1420 VSS.n1419 0.280231
R8831 VSS.n2182 VSS.n2179 0.280231
R8832 VSS.n1991 VSS 0.27984
R8833 VSS.n1995 VSS 0.27984
R8834 VSS.n1266 VSS 0.27984
R8835 VSS.n1270 VSS 0.27984
R8836 VSS.n2439 VSS 0.27984
R8837 VSS VSS.n2432 0.27984
R8838 VSS VSS.n1404 0.27984
R8839 VSS VSS.n1400 0.27984
R8840 VSS VSS.n2164 0.27984
R8841 VSS VSS.n2160 0.27984
R8842 VSS.n1612 VSS 0.27984
R8843 VSS VSS.n1609 0.27984
R8844 VSS.n906 VSS.n905 0.277931
R8845 VSS.n680 VSS.n679 0.277931
R8846 VSS.n2565 VSS.n2564 0.277167
R8847 VSS.n2563 VSS.n2562 0.277167
R8848 VSS.n3126 VSS.n285 0.277167
R8849 VSS.n3128 VSS.n3127 0.277167
R8850 VSS.n3243 VSS.n3241 0.273398
R8851 VSS.n873 VSS.n872 0.272151
R8852 VSS.n681 VSS.n602 0.272151
R8853 VSS.n1630 VSS.n786 0.268849
R8854 VSS VSS.n543 0.265394
R8855 VSS VSS.n561 0.265394
R8856 VSS.n898 VSS.n897 0.262771
R8857 VSS.n3251 VSS.n3249 0.262705
R8858 VSS VSS.n828 0.261689
R8859 VSS.n829 VSS 0.261689
R8860 VSS VSS.n579 0.259875
R8861 VSS.n580 VSS 0.259875
R8862 VSS.n879 VSS 0.259875
R8863 VSS VSS.n884 0.259875
R8864 VSS.n1848 VSS 0.259875
R8865 VSS.n1470 VSS 0.259875
R8866 VSS VSS.n844 0.258086
R8867 VSS.n845 VSS 0.258086
R8868 VSS.n1532 VSS.n1529 0.255008
R8869 VSS.n2513 VSS.n2512 0.255008
R8870 VSS.n2580 VSS.n2579 0.255008
R8871 VSS.n1915 VSS.n1912 0.255008
R8872 VSS VSS.n528 0.254582
R8873 VSS.n529 VSS 0.254582
R8874 VSS.n2696 VSS 0.254582
R8875 VSS.n2694 VSS 0.254582
R8876 VSS.n3329 VSS.n3321 0.254245
R8877 VSS.n3311 VSS.n3303 0.254245
R8878 VSS.n401 VSS.n398 0.254245
R8879 VSS.n647 VSS.n644 0.254245
R8880 VSS.n1894 VSS.n1234 0.254245
R8881 VSS.n1424 VSS.n958 0.253161
R8882 VSS.n3435 VSS.n3434 0.253109
R8883 VSS.n3433 VSS.n3432 0.253109
R8884 VSS.n1642 VSS.n806 0.252335
R8885 VSS.n3123 VSS.n3122 0.251894
R8886 VSS.n3132 VSS.n3131 0.251894
R8887 VSS.n3161 VSS.n3160 0.251419
R8888 VSS.n3146 VSS.n3145 0.250691
R8889 VSS.n3426 VSS.n51 0.250691
R8890 VSS.n801 VSS.n800 0.250683
R8891 VSS.n1999 VSS 0.250123
R8892 VSS VSS.n1257 0.250123
R8893 VSS.n2424 VSS 0.250123
R8894 VSS VSS.n1362 0.250123
R8895 VSS VSS.n2122 0.250123
R8896 VSS VSS.n1605 0.250123
R8897 VSS.n3258 VSS.n3257 0.249789
R8898 VSS.n2000 VSS.n1999 0.247195
R8899 VSS.n1257 VSS.n1256 0.247195
R8900 VSS.n2425 VSS.n2424 0.247195
R8901 VSS.n1410 VSS.n1362 0.247195
R8902 VSS.n2170 VSS.n2122 0.247195
R8903 VSS.n1605 VSS.n1604 0.247195
R8904 VSS.n3159 VSS.n262 0.246335
R8905 VSS.n2505 VSS.n2504 0.245993
R8906 VSS.n2503 VSS.n2502 0.245993
R8907 VSS VSS.n1991 0.243604
R8908 VSS VSS.n1995 0.243604
R8909 VSS VSS.n1266 0.243604
R8910 VSS VSS.n1270 0.243604
R8911 VSS VSS.n2439 0.243604
R8912 VSS.n2432 VSS 0.243604
R8913 VSS.n1404 VSS 0.243604
R8914 VSS.n1400 VSS 0.243604
R8915 VSS.n2164 VSS 0.243604
R8916 VSS.n2160 VSS 0.243604
R8917 VSS VSS.n1612 0.243604
R8918 VSS.n1609 VSS 0.243604
R8919 VSS VSS.n1558 0.240775
R8920 VSS.n3235 VSS.n3233 0.240248
R8921 VSS VSS.n796 0.23417
R8922 VSS.n4 VSS.n3 0.233202
R8923 VSS.n804 VSS.n801 0.230041
R8924 VSS.n806 VSS.n805 0.22839
R8925 VSS.n552 VSS 0.223904
R8926 VSS.n570 VSS 0.223904
R8927 VSS.n3476 VSS 0.223676
R8928 VSS.n1713 VSS 0.223676
R8929 VSS.n956 VSS 0.222572
R8930 VSS.n836 VSS 0.22078
R8931 VSS.n3417 VSS 0.220206
R8932 VSS.n586 VSS 0.21925
R8933 VSS.n889 VSS 0.21925
R8934 VSS.n852 VSS 0.217741
R8935 VSS.n2275 VSS 0.217656
R8936 VSS VSS.n2209 0.217656
R8937 VSS.n2382 VSS 0.21683
R8938 VSS.n1945 VSS 0.21683
R8939 VSS.n2571 VSS.n956 0.215457
R8940 VSS.n536 VSS 0.214786
R8941 VSS VSS.n2691 0.214786
R8942 VSS.n786 VSS.n785 0.211876
R8943 VSS.n696 VSS.n695 0.203
R8944 VSS.n133 VSS.n131 0.202392
R8945 VSS.n138 VSS.n137 0.202392
R8946 VSS.n3358 VSS.n3357 0.202392
R8947 VSS.n3362 VSS.n3361 0.202392
R8948 VSS.n3378 VSS.n3377 0.202392
R8949 VSS.n3376 VSS.n3375 0.202392
R8950 VSS.n3398 VSS.n3397 0.202392
R8951 VSS.n3402 VSS.n3401 0.202392
R8952 VSS.n596 VSS.n595 0.202392
R8953 VSS.n599 VSS.n598 0.202392
R8954 VSS.n1644 VSS.n808 0.201142
R8955 VSS.n2459 VSS 0.199831
R8956 VSS.n2567 VSS 0.198119
R8957 VSS.n2558 VSS 0.198119
R8958 VSS.n2411 VSS 0.194611
R8959 VSS.n3160 VSS.n3159 0.194066
R8960 VSS.n3380 VSS.n108 0.193357
R8961 VSS.n2675 VSS 0.192251
R8962 VSS.n665 VSS.n664 0.19152
R8963 VSS.n878 VSS.n877 0.19152
R8964 VSS.n1488 VSS 0.191234
R8965 VSS.n1475 VSS 0.191234
R8966 VSS.n1498 VSS 0.191234
R8967 VSS.n1225 VSS 0.191234
R8968 VSS.n1099 VSS 0.191234
R8969 VSS VSS.n2302 0.191234
R8970 VSS.n2053 VSS 0.191234
R8971 VSS.n1434 VSS 0.191234
R8972 VSS.n1299 VSS 0.191234
R8973 VSS VSS.n1318 0.191234
R8974 VSS.n1949 VSS 0.191234
R8975 VSS.n3051 VSS 0.191234
R8976 VSS VSS.n1013 0.191234
R8977 VSS.n2452 VSS 0.191234
R8978 VSS VSS.n2473 0.191234
R8979 VSS.n96 VSS 0.191234
R8980 VSS.n84 VSS 0.191234
R8981 VSS VSS.n3346 0.191234
R8982 VSS.n3281 VSS 0.191234
R8983 VSS.n62 VSS 0.191234
R8984 VSS.n265 VSS 0.191234
R8985 VSS.n1052 VSS 0.191234
R8986 VSS.n1041 VSS 0.191234
R8987 VSS VSS.n994 0.191234
R8988 VSS VSS.n2483 0.191234
R8989 VSS VSS.n927 0.191234
R8990 VSS VSS.n938 0.191234
R8991 VSS.n1025 VSS 0.191234
R8992 VSS.n2996 VSS 0.191234
R8993 VSS VSS.n45 0.191234
R8994 VSS.n3458 VSS 0.191234
R8995 VSS.n464 VSS 0.191234
R8996 VSS.n480 VSS 0.191234
R8997 VSS VSS.n415 0.191234
R8998 VSS.n430 VSS 0.191234
R8999 VSS VSS.n2989 0.191234
R9000 VSS.n2545 VSS 0.191234
R9001 VSS.n1372 VSS 0.191234
R9002 VSS.n2320 VSS 0.191234
R9003 VSS VSS.n1968 0.191234
R9004 VSS VSS.n2244 0.191234
R9005 VSS.n2131 VSS 0.191234
R9006 VSS.n2087 VSS 0.191234
R9007 VSS.n2072 VSS 0.191234
R9008 VSS VSS.n2021 0.191234
R9009 VSS VSS.n2396 0.191234
R9010 VSS VSS.n1345 0.191234
R9011 VSS.n1509 VSS 0.191234
R9012 VSS.n1803 VSS 0.191234
R9013 VSS.n2636 VSS 0.191234
R9014 VSS VSS.n1640 0.191234
R9015 VSS VSS.n1626 0.191234
R9016 VSS VSS.n1585 0.191234
R9017 VSS VSS.n1879 0.191234
R9018 VSS.n2288 VSS.n1105 0.187931
R9019 VSS.n2309 VSS.n2308 0.187931
R9020 VSS.n2382 VSS.n1073 0.187931
R9021 VSS.n1291 VSS.n1290 0.187931
R9022 VSS.n1455 VSS.n1454 0.187931
R9023 VSS.n1945 VSS.n1121 0.187931
R9024 VSS.n2530 VSS.n2529 0.187931
R9025 VSS.n1350 VSS.n1349 0.187931
R9026 VSS.n1669 VSS.n1668 0.187931
R9027 VSS.n1632 VSS.n1631 0.187931
R9028 VSS.n1644 VSS.n1643 0.187931
R9029 VSS.n2606 VSS.n860 0.187704
R9030 VSS.n623 VSS.n622 0.187704
R9031 VSS.n2276 VSS.n2275 0.187105
R9032 VSS.n2337 VSS.n2336 0.187105
R9033 VSS.n2364 VSS.n2363 0.187105
R9034 VSS.n2209 VSS.n2208 0.187105
R9035 VSS.n2200 VSS.n2199 0.187105
R9036 VSS.n2191 VSS.n2190 0.187105
R9037 VSS.n816 VSS.n812 0.18628
R9038 VSS.n3206 VSS.n3205 0.18462
R9039 VSS.n3204 VSS.n3203 0.18462
R9040 VSS.n3197 VSS.n3196 0.18462
R9041 VSS.n250 VSS.n249 0.18462
R9042 VSS.n3190 VSS.n3189 0.18462
R9043 VSS.n3188 VSS.n3187 0.18462
R9044 VSS.n3181 VSS.n3180 0.18462
R9045 VSS.n3413 VSS.n72 0.18462
R9046 VSS.n2612 VSS.n2611 0.184546
R9047 VSS.n613 VSS.n612 0.184546
R9048 VSS VSS.n2530 0.183803
R9049 VSS.n1349 VSS 0.183803
R9050 VSS VSS.n7 0.182492
R9051 VSS.n1695 VSS 0.182492
R9052 VSS VSS.n31 0.180935
R9053 VSS.n1689 VSS.n1688 0.180913
R9054 VSS.n336 VSS.n335 0.180913
R9055 VSS.n3138 VSS 0.180067
R9056 VSS.n3148 VSS 0.179208
R9057 VSS.n2414 VSS.n2413 0.177259
R9058 VSS VSS.n2500 0.175852
R9059 VSS.n3267 VSS.n3266 0.175279
R9060 VSS.n3244 VSS.n3228 0.175279
R9061 VSS.n3237 VSS.n3229 0.175279
R9062 VSS.n3234 VSS.n3229 0.175279
R9063 VSS.n3242 VSS.n3228 0.175279
R9064 VSS.n3250 VSS.n3227 0.175279
R9065 VSS.n3266 VSS.n3259 0.175279
R9066 VSS.n3252 VSS.n3227 0.173855
R9067 VSS.n2517 VSS.n2516 0.168119
R9068 VSS.n2584 VSS.n2583 0.168119
R9069 VSS.n1891 VSS.n1890 0.168119
R9070 VSS.n2405 VSS.n1068 0.168096
R9071 VSS.n3326 VSS.n3325 0.168072
R9072 VSS.n3308 VSS.n3307 0.168072
R9073 VSS.n654 VSS.n653 0.168072
R9074 VSS.n408 VSS.n407 0.168072
R9075 VSS.n1922 VSS.n1921 0.168072
R9076 VSS.n1539 VSS.n1538 0.168072
R9077 VSS.n1567 VSS.n781 0.167289
R9078 VSS.n663 VSS.n662 0.165806
R9079 VSS.n2804 VSS.n759 0.165806
R9080 VSS VSS.n778 0.165638
R9081 VSS VSS.n904 0.158206
R9082 VSS VSS.n678 0.158206
R9083 VSS.n2655 VSS.n2654 0.156125
R9084 VSS.n1563 VSS.n1562 0.154904
R9085 VSS.n3263 VSS.n3262 0.15424
R9086 VSS.n227 VSS 0.152427
R9087 VSS VSS.n3219 0.152427
R9088 VSS.n2002 VSS.n2001 0.152211
R9089 VSS.n1255 VSS.n1254 0.152211
R9090 VSS.n2423 VSS.n2422 0.152211
R9091 VSS.n1601 VSS.n1600 0.152211
R9092 VSS.n1414 VSS.n1411 0.15137
R9093 VSS.n2174 VSS.n2171 0.15137
R9094 VSS.n952 VSS.n951 0.151192
R9095 VSS.n950 VSS.n949 0.151192
R9096 VSS.n2929 VSS.n2928 0.151192
R9097 VSS.n2934 VSS.n326 0.151192
R9098 VSS.n318 VSS 0.151087
R9099 VSS.n315 VSS 0.150362
R9100 VSS VSS.n550 0.147947
R9101 VSS VSS.n568 0.147947
R9102 VSS VSS.n834 0.145885
R9103 VSS VSS.n585 0.144875
R9104 VSS.n885 VSS 0.144875
R9105 VSS VSS.n115 0.144708
R9106 VSS.n3365 VSS 0.144708
R9107 VSS VSS.n81 0.144708
R9108 VSS VSS.n76 0.144708
R9109 VSS.n656 VSS 0.144708
R9110 VSS.n2666 VSS.n2665 0.144447
R9111 VSS VSS.n850 0.143879
R9112 VSS VSS.n108 0.142971
R9113 VSS.n3330 VSS.n3329 0.142796
R9114 VSS.n3312 VSS.n3311 0.142796
R9115 VSS.n648 VSS.n647 0.142796
R9116 VSS.n402 VSS.n401 0.142796
R9117 VSS.n1916 VSS.n1915 0.142796
R9118 VSS.n1533 VSS.n1532 0.142796
R9119 VSS.n1865 VSS.n1465 0.142375
R9120 VSS.n1887 VSS.n1886 0.142375
R9121 VSS.n320 VSS 0.141998
R9122 VSS VSS.n534 0.141929
R9123 VSS.n2692 VSS 0.141929
R9124 VSS.n2513 VSS.n976 0.141461
R9125 VSS.n2580 VSS.n2577 0.141461
R9126 VSS.n1895 VSS.n1894 0.141455
R9127 VSS VSS.n661 0.140092
R9128 VSS.n2805 VSS 0.140092
R9129 VSS.n2572 VSS.n2571 0.140035
R9130 VSS.n2005 VSS.n2004 0.138903
R9131 VSS.n1279 VSS.n1278 0.138903
R9132 VSS.n2419 VSS.n2416 0.138903
R9133 VSS.n1419 VSS.n1418 0.138903
R9134 VSS.n2179 VSS.n2178 0.138903
R9135 VSS.n1598 VSS.n1595 0.138903
R9136 VSS.n2682 VSS.n2681 0.138304
R9137 VSS.n1730 VSS 0.137685
R9138 VSS VSS.n1866 0.137685
R9139 VSS VSS.n1236 0.137685
R9140 VSS.n1550 VSS 0.137685
R9141 VSS VSS.n2289 0.137685
R9142 VSS.n2307 VSS 0.137685
R9143 VSS VSS.n2383 0.137685
R9144 VSS.n1324 VSS 0.137685
R9145 VSS VSS.n1305 0.137685
R9146 VSS.n1946 VSS 0.137685
R9147 VSS.n3060 VSS 0.137685
R9148 VSS.n3048 VSS 0.137685
R9149 VSS VSS.n243 0.137685
R9150 VSS VSS.n2460 0.137685
R9151 VSS VSS.n254 0.137685
R9152 VSS.n3411 VSS 0.137685
R9153 VSS.n3424 VSS 0.137685
R9154 VSS.n3151 VSS 0.137685
R9155 VSS VSS.n969 0.137685
R9156 VSS VSS.n3161 0.137685
R9157 VSS VSS.n327 0.137685
R9158 VSS VSS.n325 0.137685
R9159 VSS VSS.n965 0.137685
R9160 VSS.n1431 VSS 0.137685
R9161 VSS VSS.n1067 0.137685
R9162 VSS.n1524 VSS 0.137685
R9163 VSS.n1799 VSS 0.137685
R9164 VSS.n3327 VSS.n3326 0.137391
R9165 VSS.n3309 VSS.n3308 0.137391
R9166 VSS.n653 VSS.n652 0.137391
R9167 VSS.n407 VSS.n406 0.137391
R9168 VSS.n1921 VSS.n1920 0.137391
R9169 VSS.n1538 VSS.n1537 0.137391
R9170 VSS.n2669 VSS.n2668 0.137236
R9171 VSS.n1348 VSS 0.137136
R9172 VSS VSS.n79 0.137136
R9173 VSS VSS.n3381 0.137136
R9174 VSS VSS.n113 0.137136
R9175 VSS.n3171 VSS 0.137136
R9176 VSS VSS.n2507 0.137136
R9177 VSS VSS.n287 0.137136
R9178 VSS VSS.n3438 0.137136
R9179 VSS VSS.n370 0.137136
R9180 VSS.n476 VSS 0.137136
R9181 VSS VSS.n356 0.137136
R9182 VSS VSS.n425 0.137136
R9183 VSS VSS.n1078 0.137136
R9184 VSS.n2334 VSS 0.137136
R9185 VSS VSS.n1971 0.137136
R9186 VSS VSS.n2249 0.137136
R9187 VSS VSS.n2109 0.137136
R9188 VSS VSS.n2046 0.137136
R9189 VSS VSS.n2032 0.137136
R9190 VSS VSS.n2218 0.137136
R9191 VSS.n1930 VSS 0.137136
R9192 VSS VSS.n2648 0.137136
R9193 VSS.n1647 VSS 0.137136
R9194 VSS VSS.n1633 0.137136
R9195 VSS.n1667 VSS 0.137136
R9196 VSS.n2611 VSS.n2610 0.136634
R9197 VSS.n2516 VSS.n2515 0.136634
R9198 VSS.n2583 VSS.n2582 0.136634
R9199 VSS.n615 VSS.n613 0.136634
R9200 VSS.n3214 VSS.n3213 0.136634
R9201 VSS.n1892 VSS.n1891 0.136634
R9202 VSS.n129 VSS.n128 0.136196
R9203 VSS.n3456 VSS.n3455 0.135964
R9204 VSS.n545 VSS.n544 0.133266
R9205 VSS.n563 VSS.n562 0.133266
R9206 VSS.n544 VSS 0.132628
R9207 VSS.n562 VSS 0.132628
R9208 VSS.n1672 VSS.n1671 0.13261
R9209 VSS.n2409 VSS 0.132014
R9210 VSS.n3199 VSS 0.132014
R9211 VSS.n3192 VSS 0.132014
R9212 VSS.n3183 VSS 0.132014
R9213 VSS.n1146 VSS.n1145 0.131017
R9214 VSS.n1154 VSS.n1153 0.131017
R9215 VSS.n1163 VSS.n1161 0.131017
R9216 VSS.n1168 VSS.n1138 0.131017
R9217 VSS.n1184 VSS.n1136 0.131017
R9218 VSS.n1192 VSS.n1191 0.131017
R9219 VSS.n1195 VSS.n1128 0.131017
R9220 VSS.n1737 VSS.n1736 0.130899
R9221 VSS.n1741 VSS.n1740 0.130899
R9222 VSS.n1752 VSS.n1751 0.130899
R9223 VSS.n1757 VSS.n1756 0.130899
R9224 VSS.n694 VSS.n693 0.130643
R9225 VSS.n1770 VSS.n1769 0.130575
R9226 VSS.n1777 VSS.n1776 0.130575
R9227 VSS.n1796 VSS.n1795 0.130575
R9228 VSS.n1794 VSS.n1793 0.130575
R9229 VSS.n690 VSS 0.127807
R9230 VSS.n896 VSS 0.127807
R9231 VSS.n2689 VSS 0.127258
R9232 VSS VSS.n349 0.127258
R9233 VSS.n907 VSS.n906 0.12579
R9234 VSS.n680 VSS.n638 0.12579
R9235 VSS.n2679 VSS.n2678 0.123883
R9236 VSS.n3150 VSS 0.123833
R9237 VSS.n3173 VSS.n3172 0.120147
R9238 VSS.n3239 VSS.n3229 0.119812
R9239 VSS.n3247 VSS.n3228 0.119812
R9240 VSS.n3255 VSS.n3227 0.119812
R9241 VSS.n3266 VSS.n3265 0.119812
R9242 VSS.n1842 VSS.n1488 0.118573
R9243 VSS.n1841 VSS.n1840 0.118573
R9244 VSS.n1839 VSS.n1838 0.118573
R9245 VSS.n1480 VSS.n1479 0.118573
R9246 VSS.n1478 VSS.n1477 0.118573
R9247 VSS.n1476 VSS.n1475 0.118573
R9248 VSS.n1499 VSS.n1498 0.118573
R9249 VSS.n1502 VSS.n1501 0.118573
R9250 VSS.n1505 VSS.n1504 0.118573
R9251 VSS.n1230 VSS.n1229 0.118573
R9252 VSS.n1228 VSS.n1227 0.118573
R9253 VSS.n1226 VSS.n1225 0.118573
R9254 VSS.n1094 VSS.n1093 0.118573
R9255 VSS.n1098 VSS.n1097 0.118573
R9256 VSS.n1100 VSS.n1099 0.118573
R9257 VSS.n2295 VSS.n2294 0.118573
R9258 VSS.n2299 VSS.n2298 0.118573
R9259 VSS.n2302 VSS.n2301 0.118573
R9260 VSS.n2049 VSS.n2048 0.118573
R9261 VSS.n2056 VSS.n2055 0.118573
R9262 VSS.n2054 VSS.n2053 0.118573
R9263 VSS.n2256 VSS.n2255 0.118573
R9264 VSS.n2257 VSS.n1974 0.118573
R9265 VSS.n2287 VSS.n2286 0.118573
R9266 VSS.n2285 VSS.n2284 0.118573
R9267 VSS.n2344 VSS.n2343 0.118573
R9268 VSS.n2345 VSS.n1081 0.118573
R9269 VSS.n2381 VSS.n2380 0.118573
R9270 VSS.n2379 VSS.n2378 0.118573
R9271 VSS.n1439 VSS.n1438 0.118573
R9272 VSS.n1437 VSS.n1436 0.118573
R9273 VSS.n1435 VSS.n1434 0.118573
R9274 VSS.n1294 VSS.n1293 0.118573
R9275 VSS.n1298 VSS.n1297 0.118573
R9276 VSS.n1300 VSS.n1299 0.118573
R9277 VSS.n1311 VSS.n1310 0.118573
R9278 VSS.n1315 VSS.n1314 0.118573
R9279 VSS.n1318 VSS.n1317 0.118573
R9280 VSS.n1954 VSS.n1953 0.118573
R9281 VSS.n1952 VSS.n1951 0.118573
R9282 VSS.n1950 VSS.n1949 0.118573
R9283 VSS.n1281 VSS.n1280 0.118573
R9284 VSS.n1285 VSS.n1284 0.118573
R9285 VSS.n1244 VSS.n1243 0.118573
R9286 VSS.n1460 VSS.n1459 0.118573
R9287 VSS.n1453 VSS.n1452 0.118573
R9288 VSS.n1451 VSS.n1450 0.118573
R9289 VSS.n1944 VSS.n1943 0.118573
R9290 VSS.n1942 VSS.n1941 0.118573
R9291 VSS.n3016 VSS.n3015 0.118573
R9292 VSS.n3054 VSS.n3053 0.118573
R9293 VSS.n3052 VSS.n3051 0.118573
R9294 VSS.n1007 VSS.n1006 0.118573
R9295 VSS.n1009 VSS.n1008 0.118573
R9296 VSS.n1013 VSS.n1012 0.118573
R9297 VSS.n2447 VSS.n2446 0.118573
R9298 VSS.n2451 VSS.n2450 0.118573
R9299 VSS.n2453 VSS.n2452 0.118573
R9300 VSS.n2466 VSS.n2465 0.118573
R9301 VSS.n2470 VSS.n2469 0.118573
R9302 VSS.n2473 VSS.n2472 0.118573
R9303 VSS.n97 VSS.n96 0.118573
R9304 VSS.n100 VSS.n99 0.118573
R9305 VSS.n103 VSS.n102 0.118573
R9306 VSS.n85 VSS.n84 0.118573
R9307 VSS.n88 VSS.n87 0.118573
R9308 VSS.n91 VSS.n90 0.118573
R9309 VSS.n3346 VSS.n3345 0.118573
R9310 VSS.n3344 VSS.n3343 0.118573
R9311 VSS.n3342 VSS.n3341 0.118573
R9312 VSS.n3282 VSS.n3281 0.118573
R9313 VSS.n3285 VSS.n120 0.118573
R9314 VSS.n3287 VSS.n3286 0.118573
R9315 VSS.n57 VSS.n56 0.118573
R9316 VSS.n61 VSS.n60 0.118573
R9317 VSS.n63 VSS.n62 0.118573
R9318 VSS.n274 VSS.n265 0.118573
R9319 VSS.n273 VSS.n272 0.118573
R9320 VSS.n271 VSS.n270 0.118573
R9321 VSS.n1032 VSS.n1031 0.118573
R9322 VSS.n1034 VSS.n1033 0.118573
R9323 VSS.n1053 VSS.n1052 0.118573
R9324 VSS.n2520 VSS.n2519 0.118573
R9325 VSS.n2524 VSS.n2523 0.118573
R9326 VSS.n2532 VSS.n2531 0.118573
R9327 VSS.n2539 VSS.n2538 0.118573
R9328 VSS.n1037 VSS.n1036 0.118573
R9329 VSS.n1044 VSS.n1043 0.118573
R9330 VSS.n1042 VSS.n1041 0.118573
R9331 VSS.n994 VSS.n993 0.118573
R9332 VSS.n992 VSS.n991 0.118573
R9333 VSS.n990 VSS.n989 0.118573
R9334 VSS.n2479 VSS.n2478 0.118573
R9335 VSS.n2481 VSS.n2480 0.118573
R9336 VSS.n2483 VSS.n2482 0.118573
R9337 VSS.n920 VSS.n919 0.118573
R9338 VSS.n924 VSS.n923 0.118573
R9339 VSS.n927 VSS.n926 0.118573
R9340 VSS.n934 VSS.n933 0.118573
R9341 VSS.n936 VSS.n935 0.118573
R9342 VSS.n938 VSS.n937 0.118573
R9343 VSS.n1019 VSS.n1018 0.118573
R9344 VSS.n1021 VSS.n1020 0.118573
R9345 VSS.n1026 VSS.n1025 0.118573
R9346 VSS.n3005 VSS.n2996 0.118573
R9347 VSS.n3004 VSS.n3003 0.118573
R9348 VSS.n3002 VSS.n3001 0.118573
R9349 VSS.n45 VSS.n44 0.118573
R9350 VSS.n43 VSS.n42 0.118573
R9351 VSS.n41 VSS.n40 0.118573
R9352 VSS.n3463 VSS.n3462 0.118573
R9353 VSS.n3461 VSS.n3460 0.118573
R9354 VSS.n3459 VSS.n3458 0.118573
R9355 VSS.n465 VSS.n464 0.118573
R9356 VSS.n468 VSS.n389 0.118573
R9357 VSS.n470 VSS.n469 0.118573
R9358 VSS.n481 VSS.n480 0.118573
R9359 VSS.n484 VSS.n483 0.118573
R9360 VSS.n487 VSS.n486 0.118573
R9361 VSS.n450 VSS.n415 0.118573
R9362 VSS.n453 VSS.n451 0.118573
R9363 VSS.n455 VSS.n454 0.118573
R9364 VSS.n431 VSS.n430 0.118573
R9365 VSS.n434 VSS.n419 0.118573
R9366 VSS.n436 VSS.n435 0.118573
R9367 VSS.n2983 VSS.n2982 0.118573
R9368 VSS.n2985 VSS.n2984 0.118573
R9369 VSS.n2989 VSS.n2988 0.118573
R9370 VSS.n2550 VSS.n2549 0.118573
R9371 VSS.n2548 VSS.n2547 0.118573
R9372 VSS.n2546 VSS.n2545 0.118573
R9373 VSS.n1373 VSS.n1372 0.118573
R9374 VSS.n1376 VSS.n1375 0.118573
R9375 VSS.n1379 VSS.n1378 0.118573
R9376 VSS.n2321 VSS.n2320 0.118573
R9377 VSS.n2324 VSS.n2323 0.118573
R9378 VSS.n2327 VSS.n2326 0.118573
R9379 VSS.n1968 VSS.n1967 0.118573
R9380 VSS.n1966 VSS.n1965 0.118573
R9381 VSS.n1964 VSS.n1963 0.118573
R9382 VSS.n2244 VSS.n2243 0.118573
R9383 VSS.n2242 VSS.n2241 0.118573
R9384 VSS.n2240 VSS.n2239 0.118573
R9385 VSS.n2265 VSS.n2264 0.118573
R9386 VSS.n2274 VSS.n1973 0.118573
R9387 VSS.n2313 VSS.n1087 0.118573
R9388 VSS.n2338 VSS.n2314 0.118573
R9389 VSS.n2353 VSS.n2352 0.118573
R9390 VSS.n2362 VSS.n1080 0.118573
R9391 VSS.n2373 VSS.n2372 0.118573
R9392 VSS.n2371 VSS.n1069 0.118573
R9393 VSS.n2132 VSS.n2131 0.118573
R9394 VSS.n2135 VSS.n2134 0.118573
R9395 VSS.n2138 VSS.n2137 0.118573
R9396 VSS.n2088 VSS.n2087 0.118573
R9397 VSS.n2091 VSS.n2090 0.118573
R9398 VSS.n2094 VSS.n2093 0.118573
R9399 VSS.n2073 VSS.n2072 0.118573
R9400 VSS.n2076 VSS.n2066 0.118573
R9401 VSS.n2078 VSS.n2077 0.118573
R9402 VSS.n2021 VSS.n2020 0.118573
R9403 VSS.n2019 VSS.n2018 0.118573
R9404 VSS.n2017 VSS.n2016 0.118573
R9405 VSS.n2213 VSS.n2212 0.118573
R9406 VSS.n2211 VSS.n2210 0.118573
R9407 VSS.n2204 VSS.n2203 0.118573
R9408 VSS.n2202 VSS.n2201 0.118573
R9409 VSS.n2195 VSS.n2194 0.118573
R9410 VSS.n2193 VSS.n2192 0.118573
R9411 VSS.n2186 VSS.n2185 0.118573
R9412 VSS.n2184 VSS.n2183 0.118573
R9413 VSS.n2389 VSS.n2388 0.118573
R9414 VSS.n2393 VSS.n2392 0.118573
R9415 VSS.n2396 VSS.n2395 0.118573
R9416 VSS.n1341 VSS.n1340 0.118573
R9417 VSS.n1343 VSS.n1342 0.118573
R9418 VSS.n1345 VSS.n1344 0.118573
R9419 VSS.n1331 VSS.n1330 0.118573
R9420 VSS.n1336 VSS.n1335 0.118573
R9421 VSS.n1938 VSS.n1937 0.118573
R9422 VSS.n1936 VSS.n1935 0.118573
R9423 VSS.n1824 VSS.n1509 0.118573
R9424 VSS.n1823 VSS.n1822 0.118573
R9425 VSS.n1821 VSS.n1820 0.118573
R9426 VSS.n1804 VSS.n1803 0.118573
R9427 VSS.n1807 VSS.n1806 0.118573
R9428 VSS.n1810 VSS.n1809 0.118573
R9429 VSS.n2631 VSS.n2630 0.118573
R9430 VSS.n2635 VSS.n2634 0.118573
R9431 VSS.n2637 VSS.n2636 0.118573
R9432 VSS.n1636 VSS.n1635 0.118573
R9433 VSS.n1638 VSS.n1637 0.118573
R9434 VSS.n1640 VSS.n1639 0.118573
R9435 VSS.n1622 VSS.n1621 0.118573
R9436 VSS.n1624 VSS.n1623 0.118573
R9437 VSS.n1626 VSS.n1625 0.118573
R9438 VSS.n1581 VSS.n1580 0.118573
R9439 VSS.n1583 VSS.n1582 0.118573
R9440 VSS.n1585 VSS.n1584 0.118573
R9441 VSS.n1594 VSS.n1593 0.118573
R9442 VSS.n1562 VSS.n1561 0.118573
R9443 VSS.n1570 VSS.n1569 0.118573
R9444 VSS.n1568 VSS.n1567 0.118573
R9445 VSS.n795 VSS.n794 0.118573
R9446 VSS.n800 VSS.n799 0.118573
R9447 VSS.n819 VSS.n818 0.118573
R9448 VSS.n817 VSS.n816 0.118573
R9449 VSS.n1873 VSS.n1872 0.118573
R9450 VSS.n1875 VSS.n1874 0.118573
R9451 VSS.n1879 VSS.n1878 0.118573
R9452 VSS VSS.n1765 0.116501
R9453 VSS.n2688 VSS.n2687 0.116405
R9454 VSS VSS.n2609 0.115458
R9455 VSS VSS.n2514 0.115458
R9456 VSS VSS.n2581 0.115458
R9457 VSS.n616 VSS 0.115458
R9458 VSS.n1893 VSS 0.115458
R9459 VSS.n1729 VSS 0.115271
R9460 VSS VSS.n1464 0.115271
R9461 VSS.n1549 VSS 0.115271
R9462 VSS VSS.n1125 0.115271
R9463 VSS.n1104 VSS 0.115271
R9464 VSS VSS.n1089 0.115271
R9465 VSS VSS.n1072 0.115271
R9466 VSS.n2270 VSS 0.115271
R9467 VSS VSS.n1105 0.115271
R9468 VSS VSS.n1088 0.115271
R9469 VSS VSS.n2309 0.115271
R9470 VSS.n2358 VSS 0.115271
R9471 VSS VSS.n1073 0.115271
R9472 VSS VSS.n1432 0.115271
R9473 VSS.n1304 VSS 0.115271
R9474 VSS VSS.n1247 0.115271
R9475 VSS VSS.n1947 0.115271
R9476 VSS VSS.n1249 0.115271
R9477 VSS.n1290 VSS 0.115271
R9478 VSS VSS.n1457 0.115271
R9479 VSS VSS.n1455 0.115271
R9480 VSS VSS.n1448 0.115271
R9481 VSS VSS.n1121 0.115271
R9482 VSS VSS.n3049 0.115271
R9483 VSS VSS.n1014 0.115271
R9484 VSS.n2457 VSS 0.115271
R9485 VSS VSS.n2474 0.115271
R9486 VSS VSS.n93 0.115271
R9487 VSS.n107 VSS 0.115271
R9488 VSS VSS.n3293 0.115271
R9489 VSS.n128 VSS 0.115271
R9490 VSS.n67 VSS 0.115271
R9491 VSS VSS.n260 0.115271
R9492 VSS VSS.n1050 0.115271
R9493 VSS VSS.n970 0.115271
R9494 VSS.n2529 VSS 0.115271
R9495 VSS VSS.n2536 0.115271
R9496 VSS VSS.n279 0.115271
R9497 VSS VSS.n278 0.115271
R9498 VSS.n996 VSS 0.115271
R9499 VSS VSS.n73 0.115271
R9500 VSS VSS.n928 0.115271
R9501 VSS VSS.n939 0.115271
R9502 VSS VSS.n1023 0.115271
R9503 VSS VSS.n2993 0.115271
R9504 VSS.n47 VSS 0.115271
R9505 VSS VSS.n3456 0.115271
R9506 VSS VSS.n392 0.115271
R9507 VSS VSS.n477 0.115271
R9508 VSS VSS.n446 0.115271
R9509 VSS.n423 VSS 0.115271
R9510 VSS VSS.n2975 0.115271
R9511 VSS VSS.n3152 0.115271
R9512 VSS VSS.n1423 0.115271
R9513 VSS.n1430 VSS 0.115271
R9514 VSS VSS.n1369 0.115271
R9515 VSS VSS.n2316 0.115271
R9516 VSS.n1970 VSS 0.115271
R9517 VSS.n2246 VSS 0.115271
R9518 VSS.n2248 VSS 0.115271
R9519 VSS VSS.n2261 0.115271
R9520 VSS VSS.n2276 0.115271
R9521 VSS VSS.n2279 0.115271
R9522 VSS.n2336 VSS 0.115271
R9523 VSS VSS.n2349 0.115271
R9524 VSS VSS.n2364 0.115271
R9525 VSS VSS.n2367 0.115271
R9526 VSS VSS.n2128 0.115271
R9527 VSS VSS.n2084 0.115271
R9528 VSS VSS.n2069 0.115271
R9529 VSS.n2023 VSS 0.115271
R9530 VSS.n2217 VSS 0.115271
R9531 VSS.n2215 VSS 0.115271
R9532 VSS.n2208 VSS 0.115271
R9533 VSS.n2206 VSS 0.115271
R9534 VSS.n2199 VSS 0.115271
R9535 VSS.n2197 VSS 0.115271
R9536 VSS.n2190 VSS 0.115271
R9537 VSS.n2188 VSS 0.115271
R9538 VSS VSS.n2397 0.115271
R9539 VSS.n1347 VSS 0.115271
R9540 VSS.n1339 VSS 0.115271
R9541 VSS VSS.n1350 0.115271
R9542 VSS VSS.n1933 0.115271
R9543 VSS VSS.n1931 0.115271
R9544 VSS.n1521 VSS 0.115271
R9545 VSS VSS.n1800 0.115271
R9546 VSS.n2641 VSS 0.115271
R9547 VSS VSS.n1648 0.115271
R9548 VSS.n1628 VSS 0.115271
R9549 VSS VSS.n1577 0.115271
R9550 VSS VSS.n1672 0.115271
R9551 VSS VSS.n1669 0.115271
R9552 VSS.n785 VSS 0.115271
R9553 VSS.n1631 VSS 0.115271
R9554 VSS.n805 VSS 0.115271
R9555 VSS.n1643 VSS 0.115271
R9556 VSS.n2644 VSS 0.115271
R9557 VSS.n2647 VSS 0.115271
R9558 VSS VSS.n1880 0.115271
R9559 VSS.n3328 VSS 0.114702
R9560 VSS.n3310 VSS 0.114702
R9561 VSS.n646 VSS 0.114702
R9562 VSS.n400 VSS 0.114702
R9563 VSS.n1914 VSS 0.114702
R9564 VSS.n1531 VSS 0.114702
R9565 VSS.n3201 VSS 0.114268
R9566 VSS VSS.n2003 0.113945
R9567 VSS.n1253 VSS 0.113945
R9568 VSS.n2420 VSS 0.113945
R9569 VSS.n1413 VSS 0.113945
R9570 VSS.n2173 VSS 0.113945
R9571 VSS.n1599 VSS 0.113945
R9572 VSS VSS.n3077 0.111993
R9573 VSS.n1677 VSS.n1676 0.111598
R9574 VSS.n2685 VSS 0.111331
R9575 VSS.n2672 VSS 0.111331
R9576 VSS.n3486 VSS 0.109909
R9577 VSS VSS.n1702 0.109909
R9578 VSS.n796 VSS.n795 0.109491
R9579 VSS.n3477 VSS.n3476 0.109351
R9580 VSS.n1714 VSS.n1713 0.109351
R9581 VSS.n2561 VSS.n2560 0.108595
R9582 VSS.n3150 VSS.n282 0.108595
R9583 VSS.n954 VSS 0.108137
R9584 VSS.n2923 VSS 0.108137
R9585 VSS VSS.n791 0.106575
R9586 VSS VSS.n554 0.106075
R9587 VSS.n3064 VSS.n3063 0.10529
R9588 VSS.n3024 VSS.n3022 0.10508
R9589 VSS.n1680 VSS.n1679 0.104387
R9590 VSS.n3096 VSS.n290 0.103269
R9591 VSS.n3104 VSS.n289 0.103269
R9592 VSS.n3112 VSS.n288 0.103269
R9593 VSS.n1593 VSS.n1558 0.102885
R9594 VSS.n3047 VSS.n3046 0.102565
R9595 VSS.n1730 VSS.n1729 0.10206
R9596 VSS.n1866 VSS.n1464 0.10206
R9597 VSS.n1550 VSS.n1549 0.10206
R9598 VSS.n1930 VSS.n1125 0.10206
R9599 VSS.n2289 VSS.n1104 0.10206
R9600 VSS.n2307 VSS.n1089 0.10206
R9601 VSS.n2383 VSS.n1072 0.10206
R9602 VSS.n1432 VSS.n1431 0.10206
R9603 VSS.n1305 VSS.n1304 0.10206
R9604 VSS.n1324 VSS.n1247 0.10206
R9605 VSS.n1947 VSS.n1946 0.10206
R9606 VSS.n3049 VSS.n3048 0.10206
R9607 VSS.n1014 VSS.n243 0.10206
R9608 VSS.n2460 VSS.n2457 0.10206
R9609 VSS.n2474 VSS.n254 0.10206
R9610 VSS.n93 VSS.n79 0.10206
R9611 VSS.n3381 VSS.n107 0.10206
R9612 VSS.n3293 VSS.n113 0.10206
R9613 VSS.n3424 VSS.n67 0.10206
R9614 VSS.n3171 VSS.n260 0.10206
R9615 VSS.n1050 VSS.n969 0.10206
R9616 VSS.n3161 VSS.n278 0.10206
R9617 VSS.n2507 VSS.n996 0.10206
R9618 VSS.n3411 VSS.n73 0.10206
R9619 VSS.n928 VSS.n327 0.10206
R9620 VSS.n939 VSS.n325 0.10206
R9621 VSS.n1023 VSS.n965 0.10206
R9622 VSS.n2993 VSS.n287 0.10206
R9623 VSS.n3438 VSS.n47 0.10206
R9624 VSS.n392 VSS.n370 0.10206
R9625 VSS.n477 VSS.n476 0.10206
R9626 VSS.n446 VSS.n356 0.10206
R9627 VSS.n425 VSS.n423 0.10206
R9628 VSS.n3060 VSS.n2975 0.10206
R9629 VSS.n3152 VSS.n3151 0.10206
R9630 VSS.n1369 VSS.n1078 0.10206
R9631 VSS.n2334 VSS.n2316 0.10206
R9632 VSS.n1971 VSS.n1970 0.10206
R9633 VSS.n2249 VSS.n2246 0.10206
R9634 VSS.n2128 VSS.n2109 0.10206
R9635 VSS.n2084 VSS.n2046 0.10206
R9636 VSS.n2069 VSS.n2032 0.10206
R9637 VSS.n2218 VSS.n2023 0.10206
R9638 VSS.n2397 VSS.n1067 0.10206
R9639 VSS.n1348 VSS.n1347 0.10206
R9640 VSS.n1524 VSS.n1521 0.10206
R9641 VSS.n1800 VSS.n1799 0.10206
R9642 VSS.n2648 VSS.n2641 0.10206
R9643 VSS.n1648 VSS.n1647 0.10206
R9644 VSS.n1633 VSS.n1628 0.10206
R9645 VSS.n1667 VSS.n1577 0.10206
R9646 VSS.n1880 VSS.n1236 0.10206
R9647 VSS.n3037 VSS.n29 0.101682
R9648 VSS.n3437 VSS.n3436 0.0985362
R9649 VSS.n2572 VSS 0.0983618
R9650 VSS.n3067 VSS.n3066 0.0971733
R9651 VSS VSS.n1552 0.0936421
R9652 VSS VSS.n1545 0.0936421
R9653 VSS.n1780 VSS 0.0934104
R9654 VSS VSS.n1791 0.0934104
R9655 VSS.n1765 VSS 0.09252
R9656 VSS.n543 VSS.n542 0.0917766
R9657 VSS.n546 VSS.n545 0.0917766
R9658 VSS.n550 VSS.n549 0.0917766
R9659 VSS.n561 VSS.n560 0.0917766
R9660 VSS.n564 VSS.n563 0.0917766
R9661 VSS.n568 VSS.n567 0.0917766
R9662 VSS.n828 VSS.n827 0.0905
R9663 VSS.n830 VSS.n829 0.0905
R9664 VSS.n834 VSS.n833 0.0905
R9665 VSS.n2687 VSS 0.0905
R9666 VSS.n579 VSS.n578 0.089875
R9667 VSS.n581 VSS.n580 0.089875
R9668 VSS.n585 VSS.n584 0.089875
R9669 VSS.n880 VSS.n879 0.089875
R9670 VSS.n884 VSS.n883 0.089875
R9671 VSS.n886 VSS.n885 0.089875
R9672 VSS.n1849 VSS.n1848 0.089875
R9673 VSS.n1853 VSS.n1852 0.089875
R9674 VSS.n1864 VSS.n1470 0.089875
R9675 VSS.n1469 VSS.n1468 0.089875
R9676 VSS.n3487 VSS.n3486 0.0895055
R9677 VSS.n1702 VSS.n1701 0.0895055
R9678 VSS.n844 VSS.n843 0.0892586
R9679 VSS.n846 VSS.n845 0.0892586
R9680 VSS.n850 VSS.n849 0.0892586
R9681 VSS.n553 VSS 0.0892234
R9682 VSS.n571 VSS 0.0892234
R9683 VSS.n528 VSS.n527 0.088051
R9684 VSS.n530 VSS.n529 0.088051
R9685 VSS.n534 VSS.n533 0.088051
R9686 VSS.n2697 VSS.n2696 0.088051
R9687 VSS.n2695 VSS.n2694 0.088051
R9688 VSS.n2693 VSS.n2692 0.088051
R9689 VSS.n677 VSS 0.0879825
R9690 VSS VSS.n835 0.0879825
R9691 VSS.n902 VSS 0.0879825
R9692 VSS VSS.n498 0.087375
R9693 VSS.n890 VSS 0.087375
R9694 VSS.n1856 VSS 0.087375
R9695 VSS VSS.n1465 0.087375
R9696 VSS VSS.n1237 0.087375
R9697 VSS.n1886 VSS 0.087375
R9698 VSS.n7 VSS.n6 0.0869264
R9699 VSS.n1696 VSS.n1695 0.0869264
R9700 VSS VSS.n851 0.0867759
R9701 VSS VSS.n535 0.085602
R9702 VSS VSS.n2690 0.085602
R9703 VSS VSS.n3480 0.085027
R9704 VSS VSS.n3478 0.085027
R9705 VSS.n1709 VSS 0.085027
R9706 VSS VSS.n1715 0.085027
R9707 VSS.n1680 VSS.n1563 0.0847202
R9708 VSS.n1677 VSS.n1671 0.0847202
R9709 VSS.n2687 VSS.n778 0.0847202
R9710 VSS.n2682 VSS.n781 0.0847202
R9711 VSS.n2679 VSS.n786 0.0847202
R9712 VSS.n2676 VSS.n790 0.0847202
R9713 VSS.n2673 VSS.n796 0.0847202
R9714 VSS.n2669 VSS.n801 0.0847202
R9715 VSS.n2666 VSS.n806 0.0847202
R9716 VSS.n2663 VSS.n808 0.0847202
R9717 VSS.n2658 VSS.n812 0.0847202
R9718 VSS.n1683 VSS.n1558 0.0847202
R9719 VSS.n3215 VSS.n3214 0.0844496
R9720 VSS.n3185 VSS 0.0835282
R9721 VSS.n3030 VSS.n3027 0.08348
R9722 VSS.n1632 VSS.n790 0.0814174
R9723 VSS.n3355 VSS.n3354 0.0790328
R9724 VSS.n3380 VSS.n3379 0.0790328
R9725 VSS.n3395 VSS.n3394 0.0790328
R9726 VSS.n592 VSS.n384 0.0790328
R9727 VSS.n554 VSS.n553 0.0790106
R9728 VSS.n572 VSS.n571 0.0790106
R9729 VSS.n3354 VSS 0.0779904
R9730 VSS.n3394 VSS 0.0779904
R9731 VSS.n835 VSS.n791 0.0779126
R9732 VSS.n906 VSS.n873 0.0777727
R9733 VSS.n681 VSS.n680 0.0777727
R9734 VSS.n690 VSS.n498 0.077375
R9735 VSS.n896 VSS.n890 0.077375
R9736 VSS.n1683 VSS 0.0768798
R9737 VSS.n851 VSS.n809 0.0768448
R9738 VSS.n3416 VSS.n71 0.0762059
R9739 VSS.n3418 VSS.n3417 0.0762059
R9740 VSS.n2662 VSS 0.0760786
R9741 VSS.n1691 VSS.n1689 0.0760505
R9742 VSS.n335 VSS.n1 0.0760505
R9743 VSS.n535 VSS.n349 0.0758061
R9744 VSS.n2690 VSS.n2689 0.0758061
R9745 VSS.n3044 VSS 0.0753497
R9746 VSS.n3069 VSS 0.0753497
R9747 VSS VSS.n16 0.0752
R9748 VSS VSS.n3173 0.0740882
R9749 VSS VSS.n3176 0.0740882
R9750 VSS.n317 VSS.n315 0.0739862
R9751 VSS.n3220 VSS.n227 0.0739862
R9752 VSS.n3219 VSS.n3218 0.0739862
R9753 VSS.n3071 VSS 0.0733657
R9754 VSS.n715 VSS.n714 0.0730937
R9755 VSS.n666 VSS.n665 0.073051
R9756 VSS.n877 VSS.n876 0.073051
R9757 VSS.n854 VSS.n809 0.0727596
R9758 VSS.n3202 VSS.n3201 0.0724366
R9759 VSS.n2459 VSS.n2458 0.0724366
R9760 VSS.n3186 VSS.n3185 0.0724366
R9761 VSS.n573 VSS.n572 0.0718942
R9762 VSS VSS.n2936 0.0717187
R9763 VSS.n2602 VSS.n866 0.071566
R9764 VSS.n632 VSS.n607 0.071566
R9765 VSS.n1941 VSS.n958 0.0715092
R9766 VSS.n729 VSS.n728 0.0714745
R9767 VSS.n2605 VSS.n2604 0.0706762
R9768 VSS.n625 VSS.n624 0.0706762
R9769 VSS.n705 VSS.n704 0.0699903
R9770 VSS.n752 VSS 0.0695388
R9771 VSS.n3490 VSS 0.0691188
R9772 VSS VSS.n1693 0.0691188
R9773 VSS.n3248 VSS 0.0690321
R9774 VSS.n2568 VSS.n2567 0.0685952
R9775 VSS.n2566 VSS.n2565 0.0685952
R9776 VSS.n2559 VSS.n2558 0.0685952
R9777 VSS.n2557 VSS.n285 0.0685952
R9778 VSS.n3264 VSS.n3263 0.0682064
R9779 VSS.n892 VSS.n891 0.0675755
R9780 VSS.n908 VSS.n907 0.0675755
R9781 VSS.n2613 VSS.n2612 0.0675755
R9782 VSS.n860 VSS.n859 0.0675755
R9783 VSS.n1990 VSS.n1989 0.0675755
R9784 VSS.n1994 VSS.n1993 0.0675755
R9785 VSS.n1998 VSS.n1997 0.0675755
R9786 VSS.n1265 VSS.n1264 0.0675755
R9787 VSS.n1269 VSS.n1268 0.0675755
R9788 VSS.n1273 VSS.n1272 0.0675755
R9789 VSS.n3410 VSS.n3409 0.0675755
R9790 VSS.n3158 VSS.n3157 0.0675755
R9791 VSS.n2438 VSS.n2437 0.0675755
R9792 VSS.n2442 VSS.n2441 0.0675755
R9793 VSS.n2429 VSS.n2428 0.0675755
R9794 VSS.n683 VSS.n682 0.0675755
R9795 VSS.n638 VSS.n637 0.0675755
R9796 VSS.n622 VSS.n621 0.0675755
R9797 VSS.n612 VSS.n611 0.0675755
R9798 VSS.n3483 VSS.n3482 0.0675755
R9799 VSS.n1422 VSS.n1421 0.0675755
R9800 VSS.n2181 VSS.n2180 0.0675755
R9801 VSS.n1929 VSS.n1928 0.0675755
R9802 VSS.n1707 VSS.n1706 0.0675755
R9803 VSS.n1687 VSS.n1686 0.0675755
R9804 VSS.n1617 VSS.n1616 0.0675755
R9805 VSS.n1611 VSS.n1610 0.0675755
R9806 VSS.n1607 VSS.n1606 0.0675755
R9807 VSS.n332 VSS.n331 0.0675755
R9808 VSS VSS.n694 0.0671607
R9809 VSS.n747 VSS.n746 0.0671567
R9810 VSS.n319 VSS.n318 0.066973
R9811 VSS.n1732 VSS.n1485 0.0667264
R9812 VSS.n3331 VSS.n3330 0.0667264
R9813 VSS.n3313 VSS.n3312 0.0667264
R9814 VSS.n1405 VSS.n1389 0.0667264
R9815 VSS.n1397 VSS.n1396 0.0667264
R9816 VSS.n1402 VSS.n1401 0.0667264
R9817 VSS.n649 VSS.n648 0.0667264
R9818 VSS.n403 VSS.n402 0.0667264
R9819 VSS.n2165 VSS.n2149 0.0667264
R9820 VSS.n2162 VSS.n2161 0.0667264
R9821 VSS.n2158 VSS.n2157 0.0667264
R9822 VSS.n1917 VSS.n1916 0.0667264
R9823 VSS.n1534 VSS.n1533 0.0667264
R9824 VSS.n3072 VSS.n322 0.0666983
R9825 VSS VSS.n2563 0.0666905
R9826 VSS VSS.n2561 0.0666905
R9827 VSS.n3127 VSS 0.0666905
R9828 VSS VSS.n282 0.0666905
R9829 VSS VSS.n2655 0.0666607
R9830 VSS.n3095 VSS.n3094 0.0664039
R9831 VSS.n3170 VSS.n262 0.066226
R9832 VSS.n2407 VSS.n2406 0.0659808
R9833 VSS VSS.n3267 0.0647857
R9834 VSS VSS.n3252 0.0647857
R9835 VSS VSS.n3244 0.0647857
R9836 VSS VSS.n3237 0.0647857
R9837 VSS.n3233 VSS 0.0647857
R9838 VSS VSS.n3234 0.0647857
R9839 VSS VSS.n3242 0.0647857
R9840 VSS VSS.n3250 0.0647857
R9841 VSS.n3259 VSS 0.0647857
R9842 VSS.n3103 VSS.n3102 0.0637265
R9843 VSS.n2664 VSS.n2663 0.0635267
R9844 VSS.n3432 VSS.n3431 0.0626739
R9845 VSS.n3445 VSS.n31 0.0626739
R9846 VSS.n1692 VSS 0.0624266
R9847 VSS VSS.n3491 0.0624266
R9848 VSS.n3137 VSS.n3132 0.062375
R9849 VSS.n3139 VSS.n3138 0.062375
R9850 VSS.n3149 VSS.n3148 0.0620789
R9851 VSS.n3147 VSS.n3146 0.0620789
R9852 VSS.n3078 VSS.n320 0.0618793
R9853 VSS.n3087 VSS.n305 0.061873
R9854 VSS.n2688 VSS.n777 0.0611231
R9855 VSS.n3436 VSS 0.0609348
R9856 VSS.n3434 VSS 0.0609348
R9857 VSS.n2502 VSS.n2501 0.0609225
R9858 VSS.n2500 VSS.n2499 0.0609225
R9859 VSS VSS.n3120 0.0606442
R9860 VSS.n3122 VSS 0.0606442
R9861 VSS VSS.n51 0.0603565
R9862 VSS VSS.n3425 0.0603565
R9863 VSS.n742 VSS.n741 0.0600053
R9864 VSS.n3119 VSS.n287 0.059582
R9865 VSS.n1145 VSS 0.0595367
R9866 VSS.n1153 VSS 0.0595367
R9867 VSS.n1161 VSS 0.0595367
R9868 VSS VSS.n1168 0.0595367
R9869 VSS.n1136 VSS 0.0595367
R9870 VSS VSS.n1192 0.0595367
R9871 VSS.n1128 VSS 0.0595367
R9872 VSS.n2506 VSS 0.0592324
R9873 VSS.n2504 VSS 0.0592324
R9874 VSS.n1896 VSS.n1895 0.0589403
R9875 VSS.n976 VSS.n975 0.0589274
R9876 VSS.n2577 VSS.n2576 0.0589274
R9877 VSS VSS.n2922 0.0580792
R9878 VSS.n3039 VSS.n3038 0.0573136
R9879 VSS VSS.n1148 0.0569474
R9880 VSS VSS.n1156 0.0569474
R9881 VSS.n1167 VSS 0.0569474
R9882 VSS.n1181 VSS 0.0569474
R9883 VSS VSS.n1182 0.0569474
R9884 VSS VSS.n1133 0.0569474
R9885 VSS VSS.n1193 0.0569474
R9886 VSS.n2518 VSS.n2517 0.0564843
R9887 VSS.n2585 VSS.n2584 0.0564843
R9888 VSS.n1890 VSS.n1889 0.0564843
R9889 VSS.n3240 VSS 0.0562339
R9890 VSS VSS.n3264 0.0562339
R9891 VSS.n3325 VSS.n3324 0.0557756
R9892 VSS.n3307 VSS.n3306 0.0557756
R9893 VSS.n670 VSS.n654 0.0557756
R9894 VSS.n409 VSS.n408 0.0557756
R9895 VSS.n1926 VSS.n1922 0.0557756
R9896 VSS.n1543 VSS.n1539 0.0557756
R9897 VSS.n2922 VSS.n2921 0.055745
R9898 VSS VSS.n2946 0.0553671
R9899 VSS VSS.n2962 0.0553671
R9900 VSS.n2947 VSS 0.0552176
R9901 VSS.n3256 VSS 0.0549954
R9902 VSS.n867 VSS 0.0548172
R9903 VSS VSS.n629 0.0548172
R9904 VSS.n710 VSS.n709 0.0542031
R9905 VSS.n3217 VSS.n3215 0.0540556
R9906 VSS.n3061 VSS 0.0537064
R9907 VSS VSS.n3110 0.053635
R9908 VSS.n424 VSS 0.0535035
R9909 VSS.n2936 VSS.n2935 0.0533747
R9910 VSS VSS.n14 0.0532782
R9911 VSS.n1766 VSS 0.0526154
R9912 VSS.n1681 VSS.n1680 0.051776
R9913 VSS.n3074 VSS.n3073 0.0514681
R9914 VSS.n1734 VSS.n1733 0.0512232
R9915 VSS.n1749 VSS.n1748 0.0512232
R9916 VSS.n1767 VSS.n1766 0.051097
R9917 VSS.n1798 VSS.n1797 0.051097
R9918 VSS.n2677 VSS.n2676 0.0507077
R9919 VSS.n1748 VSS 0.0505499
R9920 VSS.n1798 VSS 0.0504254
R9921 VSS.n3087 VSS 0.0502725
R9922 VSS.n137 VSS.n136 0.0501911
R9923 VSS.n3353 VSS.n115 0.0501911
R9924 VSS.n3364 VSS.n3362 0.0501911
R9925 VSS.n3366 VSS.n3365 0.0501911
R9926 VSS.n3375 VSS.n3374 0.0501911
R9927 VSS.n3393 VSS.n81 0.0501911
R9928 VSS.n3403 VSS.n3402 0.0501911
R9929 VSS.n3407 VSS.n76 0.0501911
R9930 VSS.n600 VSS.n599 0.0501911
R9931 VSS.n669 VSS.n656 0.0501911
R9932 VSS.n2955 VSS 0.0495365
R9933 VSS VSS.n130 0.0488012
R9934 VSS VSS.n133 0.0488012
R9935 VSS VSS.n3355 0.0488012
R9936 VSS.n3357 VSS 0.0488012
R9937 VSS.n3379 VSS 0.0488012
R9938 VSS.n3377 VSS 0.0488012
R9939 VSS VSS.n3395 0.0488012
R9940 VSS.n3397 VSS 0.0488012
R9941 VSS VSS.n592 0.0488012
R9942 VSS VSS.n596 0.0488012
R9943 VSS.n3040 VSS.n3039 0.048476
R9944 VSS.n2410 VSS.n2409 0.0458169
R9945 VSS.n3207 VSS.n3206 0.0458169
R9946 VSS.n3200 VSS.n3199 0.0458169
R9947 VSS.n3198 VSS.n3197 0.0458169
R9948 VSS.n3193 VSS.n3192 0.0458169
R9949 VSS.n3191 VSS.n3190 0.0458169
R9950 VSS.n3184 VSS.n3183 0.0458169
R9951 VSS.n3182 VSS.n3181 0.0458169
R9952 VSS.n2942 VSS.n2941 0.0455
R9953 VSS.n2606 VSS.n2605 0.0449053
R9954 VSS.n624 VSS.n623 0.0449053
R9955 VSS.n1678 VSS.n1677 0.0445653
R9956 VSS VSS.n3204 0.0445493
R9957 VSS VSS.n3202 0.0445493
R9958 VSS.n249 VSS 0.0445493
R9959 VSS.n2458 VSS 0.0445493
R9960 VSS VSS.n3188 0.0445493
R9961 VSS VSS.n3186 0.0445493
R9962 VSS VSS.n72 0.0445493
R9963 VSS VSS.n3412 0.0445493
R9964 VSS.n3088 VSS.n3087 0.0423182
R9965 VSS.n3062 VSS.n3061 0.0414419
R9966 VSS.n3047 VSS.n3031 0.04136
R9967 VSS VSS.n1068 0.0405962
R9968 VSS.n2406 VSS 0.0405962
R9969 VSS.n3485 VSS.n3484 0.04
R9970 VSS.n1704 VSS.n1703 0.04
R9971 VSS.n724 VSS.n723 0.0397654
R9972 VSS.n1685 VSS.n1684 0.0386899
R9973 VSS.n1682 VSS.n1681 0.0386899
R9974 VSS.n2686 VSS.n2685 0.0386899
R9975 VSS.n2684 VSS.n2683 0.0386899
R9976 VSS.n2671 VSS.n2670 0.0386899
R9977 VSS.n2661 VSS.n2660 0.0386899
R9978 VSS.n696 VSS.n384 0.0383764
R9979 VSS.n897 VSS 0.0377321
R9980 VSS VSS.n1678 0.0376217
R9981 VSS VSS.n777 0.0376217
R9982 VSS VSS.n2680 0.0376217
R9983 VSS VSS.n2677 0.0376217
R9984 VSS VSS.n2667 0.0376217
R9985 VSS VSS.n2664 0.0376217
R9986 VSS.n955 VSS.n954 0.0375893
R9987 VSS.n953 VSS.n952 0.0375893
R9988 VSS.n2924 VSS.n2923 0.0375893
R9989 VSS.n2928 VSS.n2927 0.0375893
R9990 VSS.n3241 VSS.n3240 0.0372431
R9991 VSS.n3257 VSS.n3256 0.0372431
R9992 VSS.n3076 VSS 0.0366794
R9993 VSS VSS.n950 0.0365519
R9994 VSS VSS.n328 0.0365519
R9995 VSS VSS.n326 0.0365519
R9996 VSS.n2935 VSS 0.0365519
R9997 VSS.n2602 VSS.n864 0.036033
R9998 VSS.n632 VSS.n605 0.036033
R9999 VSS.n554 VSS.n363 0.036
R10000 VSS.n1684 VSS.n1683 0.034951
R10001 VSS.n2658 VSS.n2657 0.0344169
R10002 VSS.n1147 VSS 0.0340526
R10003 VSS.n1155 VSS 0.0340526
R10004 VSS VSS.n1162 0.0340526
R10005 VSS VSS.n1137 0.0340526
R10006 VSS VSS.n1183 0.0340526
R10007 VSS VSS.n1194 0.0340526
R10008 VSS.n1742 VSS.n1741 0.0325948
R10009 VSS.n1747 VSS.n1552 0.0325948
R10010 VSS.n1758 VSS.n1757 0.0325948
R10011 VSS.n1764 VSS.n1545 0.0325948
R10012 VSS.n1779 VSS.n1777 0.0325149
R10013 VSS.n1781 VSS.n1780 0.0325149
R10014 VSS.n1793 VSS.n1792 0.0325149
R10015 VSS.n1791 VSS.n911 0.0325149
R10016 VSS.n3217 VSS.n231 0.032289
R10017 VSS.n2680 VSS.n2679 0.0322804
R10018 VSS.n725 VSS.n724 0.0322091
R10019 VSS VSS.n1190 0.0320789
R10020 VSS VSS.n1734 0.031697
R10021 VSS.n1736 VSS 0.031697
R10022 VSS VSS.n1749 0.031697
R10023 VSS.n1751 VSS 0.031697
R10024 VSS.n572 VSS.n377 0.0316538
R10025 VSS VSS.n1767 0.0316194
R10026 VSS.n1769 VSS 0.0316194
R10027 VSS.n1797 VSS 0.0316194
R10028 VSS.n1795 VSS 0.0316194
R10029 VSS VSS.n3088 0.0311818
R10030 VSS.n733 VSS.n732 0.0309948
R10031 VSS VSS.n733 0.03059
R10032 VSS.n3455 VSS 0.030089
R10033 VSS.n3088 VSS.n307 0.0295323
R10034 VSS.n3093 VSS 0.0289211
R10035 VSS.n3101 VSS 0.0289211
R10036 VSS.n3109 VSS 0.0289211
R10037 VSS.n3117 VSS 0.0289211
R10038 VSS VSS.n2953 0.0278588
R10039 VSS.n2673 VSS.n2672 0.0277404
R10040 VSS.n2941 VSS.n2940 0.0272608
R10041 VSS.n2946 VSS.n2945 0.0272608
R10042 VSS.n2948 VSS.n2947 0.0272608
R10043 VSS.n2953 VSS.n2952 0.0272608
R10044 VSS.n2957 VSS.n2956 0.0272608
R10045 VSS.n2962 VSS.n2961 0.0272608
R10046 VSS.n2963 VSS.n323 0.0272608
R10047 VSS.n3075 VSS.n3074 0.0272608
R10048 VSS.n697 VSS 0.0270817
R10049 VSS VSS.n3217 0.026922
R10050 VSS.n693 VSS.n496 0.0265597
R10051 VSS.n2608 VSS.n2607 0.0263107
R10052 VSS.n619 VSS.n618 0.0263107
R10053 VSS.n3045 VSS.n3044 0.0262916
R10054 VSS.n3043 VSS.n3040 0.0262916
R10055 VSS.n3070 VSS.n3069 0.0262916
R10056 VSS.n3068 VSS.n3067 0.0262916
R10057 VSS.n16 VSS.n15 0.02624
R10058 VSS.n3022 VSS.n17 0.02624
R10059 VSS VSS.n3037 0.0255701
R10060 VSS.n3454 VSS 0.0255701
R10061 VSS VSS.n3064 0.0255701
R10062 VSS VSS.n3062 0.0255701
R10063 VSS.n3077 VSS.n322 0.0255299
R10064 VSS.n3025 VSS 0.02552
R10065 VSS.n3031 VSS 0.02552
R10066 VSS.n2794 VSS.n2793 0.0250946
R10067 VSS.n2787 VSS.n2786 0.0250946
R10068 VSS.n2790 VSS.n761 0.0250946
R10069 VSS.n3447 VSS.n3446 0.0248493
R10070 VSS.n753 VSS.n752 0.0242893
R10071 VSS.n751 VSS.n338 0.0242893
R10072 VSS.n3249 VSS.n3248 0.0242273
R10073 VSS.n765 VSS.n764 0.0229091
R10074 VSS.n767 VSS.n763 0.0229091
R10075 VSS.n772 VSS.n771 0.0229091
R10076 VSS.n3027 VSS.n3025 0.0221
R10077 VSS.n2879 VSS.n2878 0.0220932
R10078 VSS.n2704 VSS.n772 0.0214902
R10079 VSS.n2706 VSS.n2704 0.0214902
R10080 VSS.n2709 VSS.n2706 0.0214902
R10081 VSS.n2711 VSS.n2709 0.0214902
R10082 VSS.n2713 VSS.n2711 0.0214902
R10083 VSS.n2715 VSS.n2713 0.0214902
R10084 VSS.n2717 VSS.n2715 0.0214902
R10085 VSS.n2719 VSS.n2717 0.0214902
R10086 VSS.n2721 VSS.n2719 0.0214902
R10087 VSS.n2723 VSS.n2721 0.0214902
R10088 VSS.n2725 VSS.n2723 0.0214902
R10089 VSS.n2727 VSS.n2725 0.0214902
R10090 VSS.n2729 VSS.n2727 0.0214902
R10091 VSS.n2732 VSS.n2729 0.0214902
R10092 VSS.n2734 VSS.n2732 0.0214902
R10093 VSS.n2736 VSS.n2734 0.0214902
R10094 VSS.n2738 VSS.n2736 0.0214902
R10095 VSS.n2741 VSS.n2738 0.0214902
R10096 VSS.n2743 VSS.n2741 0.0214902
R10097 VSS.n2745 VSS.n2743 0.0214902
R10098 VSS.n2747 VSS.n2745 0.0214902
R10099 VSS.n2749 VSS.n2747 0.0214902
R10100 VSS.n2751 VSS.n2749 0.0214902
R10101 VSS.n2753 VSS.n2751 0.0214902
R10102 VSS.n2755 VSS.n2753 0.0214902
R10103 VSS.n2757 VSS.n2755 0.0214902
R10104 VSS.n2759 VSS.n2757 0.0214902
R10105 VSS.n2761 VSS.n2759 0.0214902
R10106 VSS.n2764 VSS.n2761 0.0214902
R10107 VSS.n2766 VSS.n2764 0.0214902
R10108 VSS.n2768 VSS.n2766 0.0214902
R10109 VSS.n2770 VSS.n2768 0.0214902
R10110 VSS.n2772 VSS.n2770 0.0214902
R10111 VSS.n2774 VSS.n2772 0.0214902
R10112 VSS.n2776 VSS.n2774 0.0214902
R10113 VSS.n2778 VSS.n2776 0.0214902
R10114 VSS.n2780 VSS.n2778 0.0214902
R10115 VSS.n2784 VSS.n2780 0.0214902
R10116 VSS.n2785 VSS.n2784 0.0214902
R10117 VSS.n2787 VSS.n2785 0.0214902
R10118 VSS.n2798 VSS.n2794 0.0214902
R10119 VSS.n2800 VSS.n2798 0.0214902
R10120 VSS.n2801 VSS.n2800 0.0214902
R10121 VSS.n2801 VSS.n757 0.0214902
R10122 VSS.n2809 VSS.n757 0.0214902
R10123 VSS.n2812 VSS.n2809 0.0214902
R10124 VSS.n2816 VSS.n2812 0.0214902
R10125 VSS.n2818 VSS.n2816 0.0214902
R10126 VSS.n2820 VSS.n2818 0.0214902
R10127 VSS.n2822 VSS.n2820 0.0214902
R10128 VSS.n2824 VSS.n2822 0.0214902
R10129 VSS.n2825 VSS.n2824 0.0214902
R10130 VSS.n2913 VSS.n2912 0.0214902
R10131 VSS.n2912 VSS.n2911 0.0214902
R10132 VSS.n2911 VSS.n2910 0.0214902
R10133 VSS.n2910 VSS.n2909 0.0214902
R10134 VSS.n2909 VSS.n2908 0.0214902
R10135 VSS.n2908 VSS.n2907 0.0214902
R10136 VSS.n2907 VSS.n2906 0.0214902
R10137 VSS.n2906 VSS.n2905 0.0214902
R10138 VSS.n2905 VSS.n2904 0.0214902
R10139 VSS.n2904 VSS.n2903 0.0214902
R10140 VSS.n2903 VSS.n2902 0.0214902
R10141 VSS.n2902 VSS.n2901 0.0214902
R10142 VSS.n2901 VSS.n2900 0.0214902
R10143 VSS.n2900 VSS.n2899 0.0214902
R10144 VSS.n2899 VSS.n2898 0.0214902
R10145 VSS.n2898 VSS.n2897 0.0214902
R10146 VSS.n2897 VSS.n2896 0.0214902
R10147 VSS.n2896 VSS.n2895 0.0214902
R10148 VSS.n2895 VSS.n2894 0.0214902
R10149 VSS.n2894 VSS.n2893 0.0214902
R10150 VSS.n2893 VSS.n2892 0.0214902
R10151 VSS.n2892 VSS.n2891 0.0214902
R10152 VSS.n2891 VSS.n2890 0.0214902
R10153 VSS.n2890 VSS.n2889 0.0214902
R10154 VSS.n2889 VSS.n2888 0.0214902
R10155 VSS.n2888 VSS.n2887 0.0214902
R10156 VSS.n2887 VSS.n2886 0.0214902
R10157 VSS.n2886 VSS.n2885 0.0214902
R10158 VSS.n2885 VSS.n2884 0.0214902
R10159 VSS.n2884 VSS.n2883 0.0214902
R10160 VSS.n2883 VSS.n2882 0.0214902
R10161 VSS.n2882 VSS.n2881 0.0214902
R10162 VSS.n2881 VSS.n2880 0.0214902
R10163 VSS.n2880 VSS.n2879 0.0214902
R10164 VSS.n870 VSS.n868 0.0211167
R10165 VSS.n628 VSS.n627 0.0211167
R10166 VSS VSS.n700 0.0206049
R10167 VSS.n3095 VSS 0.0205495
R10168 VSS VSS.n3096 0.0205495
R10169 VSS.n741 VSS.n740 0.0197954
R10170 VSS.n739 VSS.n738 0.0197954
R10171 VSS.n737 VSS.n736 0.0197954
R10172 VSS.n735 VSS.n734 0.0197954
R10173 VSS.n723 VSS.n722 0.0197954
R10174 VSS.n704 VSS.n703 0.0197954
R10175 VSS.n702 VSS.n701 0.0197954
R10176 VSS.n700 VSS.n699 0.0197954
R10177 VSS.n698 VSS.n697 0.0197954
R10178 VSS.n664 VSS.n663 0.0197857
R10179 VSS.n878 VSS.n759 0.0197857
R10180 VSS.n743 VSS.n742 0.0193906
R10181 VSS VSS.n338 0.0192985
R10182 VSS.n424 VSS.n339 0.0192556
R10183 VSS VSS.n712 0.0192556
R10184 VSS.n711 VSS 0.0192556
R10185 VSS VSS.n708 0.0192556
R10186 VSS.n707 VSS 0.0192556
R10187 VSS.n3076 VSS.n323 0.0191877
R10188 VSS.n2670 VSS.n2669 0.0189273
R10189 VSS.n721 VSS.n720 0.0181762
R10190 VSS.n719 VSS.n718 0.0181762
R10191 VSS.n2917 VSS.n2916 0.0179878
R10192 VSS.n2683 VSS.n2682 0.017859
R10193 VSS VSS.n14 0.01778
R10194 VSS.n717 VSS.n716 0.0175015
R10195 VSS.n3046 VSS 0.0163717
R10196 VSS VSS.n808 0.0161881
R10197 VSS.n1148 VSS 0.0158947
R10198 VSS.n1156 VSS 0.0158947
R10199 VSS VSS.n1167 0.0158947
R10200 VSS VSS.n1181 0.0158947
R10201 VSS.n1182 VSS 0.0158947
R10202 VSS VSS.n1133 0.0158947
R10203 VSS.n1193 VSS 0.0158947
R10204 VSS VSS.n696 0.0158823
R10205 VSS.n2660 VSS 0.0154555
R10206 VSS.n2829 VSS.n2828 0.0147144
R10207 VSS.n2919 VSS.n2918 0.0143015
R10208 VSS VSS.n307 0.0135645
R10209 VSS.n2825 VSS 0.013536
R10210 VSS.n2918 VSS.n2917 0.0131167
R10211 VSS.n2676 VSS.n2675 0.0130519
R10212 VSS.n2914 VSS.n2913 0.012063
R10213 VSS.n738 VSS.n737 0.0119693
R10214 VSS.n2667 VSS.n2666 0.0117166
R10215 VSS.n341 VSS 0.0116994
R10216 VSS VSS.n342 0.0116994
R10217 VSS VSS.n745 0.0116994
R10218 VSS.n744 VSS 0.0116994
R10219 VSS.n766 VSS.n765 0.011474
R10220 VSS.n772 VSS.n769 0.011474
R10221 VSS.n2789 VSS.n2787 0.011474
R10222 VSS.n2791 VSS.n2790 0.011474
R10223 VSS.n769 VSS.n767 0.011474
R10224 VSS.n2790 VSS.n2789 0.011474
R10225 VSS.n2794 VSS.n2791 0.011474
R10226 VSS.n767 VSS.n766 0.011474
R10227 VSS.n2674 VSS.n2673 0.0114496
R10228 VSS.n734 VSS 0.0108898
R10229 VSS.n2942 VSS 0.0103671
R10230 VSS.n2607 VSS.n2606 0.00961702
R10231 VSS.n623 VSS.n619 0.00961702
R10232 VSS.n706 VSS.n705 0.00940555
R10233 VSS.n3111 VSS 0.00935583
R10234 VSS.n3066 VSS.n3065 0.00861623
R10235 VSS.n2828 VSS 0.00845417
R10236 VSS.n342 VSS.n341 0.00805622
R10237 VSS.n745 VSS.n744 0.00805622
R10238 VSS.n701 VSS 0.00805622
R10239 VSS.n732 VSS.n731 0.00792129
R10240 VSS.n730 VSS.n729 0.00792129
R10241 VSS.n728 VSS.n727 0.00792129
R10242 VSS.n726 VSS.n725 0.00792129
R10243 VSS.n308 VSS 0.00654839
R10244 VSS.n868 VSS.n867 0.00644714
R10245 VSS.n629 VSS.n628 0.00644714
R10246 VSS.n2956 VSS.n2955 0.00633057
R10247 VSS.n714 VSS.n713 0.0063021
R10248 VSS.n3073 VSS.n3071 0.00627154
R10249 VSS.n2835 VSS.n2832 0.00622306
R10250 VSS.n2835 VSS.n2834 0.00622306
R10251 VSS.n712 VSS.n711 0.0058973
R10252 VSS.n708 VSS.n707 0.0058973
R10253 VSS.n2915 VSS.n2837 0.00570865
R10254 VSS.n2915 VSS.n2914 0.00570865
R10255 VSS.n1842 VSS 0.00545413
R10256 VSS.n1840 VSS 0.00545413
R10257 VSS.n1838 VSS 0.00545413
R10258 VSS.n1480 VSS 0.00545413
R10259 VSS VSS.n1478 0.00545413
R10260 VSS VSS.n1476 0.00545413
R10261 VSS VSS.n1499 0.00545413
R10262 VSS VSS.n1502 0.00545413
R10263 VSS.n1505 VSS 0.00545413
R10264 VSS.n1230 VSS 0.00545413
R10265 VSS VSS.n1228 0.00545413
R10266 VSS VSS.n1226 0.00545413
R10267 VSS.n1094 VSS 0.00545413
R10268 VSS.n1097 VSS 0.00545413
R10269 VSS.n1100 VSS 0.00545413
R10270 VSS.n2295 VSS 0.00545413
R10271 VSS.n2298 VSS 0.00545413
R10272 VSS.n2301 VSS 0.00545413
R10273 VSS.n2048 VSS 0.00545413
R10274 VSS.n2056 VSS 0.00545413
R10275 VSS VSS.n2054 0.00545413
R10276 VSS.n2255 VSS 0.00545413
R10277 VSS.n2257 VSS 0.00545413
R10278 VSS VSS.n2287 0.00545413
R10279 VSS VSS.n2285 0.00545413
R10280 VSS.n2343 VSS 0.00545413
R10281 VSS.n2345 VSS 0.00545413
R10282 VSS VSS.n2381 0.00545413
R10283 VSS VSS.n2379 0.00545413
R10284 VSS.n1439 VSS 0.00545413
R10285 VSS VSS.n1437 0.00545413
R10286 VSS VSS.n1435 0.00545413
R10287 VSS.n1294 VSS 0.00545413
R10288 VSS.n1297 VSS 0.00545413
R10289 VSS.n1300 VSS 0.00545413
R10290 VSS.n1311 VSS 0.00545413
R10291 VSS.n1314 VSS 0.00545413
R10292 VSS.n1317 VSS 0.00545413
R10293 VSS.n1954 VSS 0.00545413
R10294 VSS VSS.n1952 0.00545413
R10295 VSS VSS.n1950 0.00545413
R10296 VSS.n1281 VSS 0.00545413
R10297 VSS.n1284 VSS 0.00545413
R10298 VSS VSS.n1243 0.00545413
R10299 VSS.n1460 VSS 0.00545413
R10300 VSS VSS.n1453 0.00545413
R10301 VSS VSS.n1451 0.00545413
R10302 VSS VSS.n1944 0.00545413
R10303 VSS VSS.n1942 0.00545413
R10304 VSS.n3015 VSS 0.00545413
R10305 VSS.n3054 VSS 0.00545413
R10306 VSS VSS.n3052 0.00545413
R10307 VSS.n1006 VSS 0.00545413
R10308 VSS.n1009 VSS 0.00545413
R10309 VSS.n1012 VSS 0.00545413
R10310 VSS.n2447 VSS 0.00545413
R10311 VSS.n2450 VSS 0.00545413
R10312 VSS.n2453 VSS 0.00545413
R10313 VSS.n2466 VSS 0.00545413
R10314 VSS.n2469 VSS 0.00545413
R10315 VSS.n2472 VSS 0.00545413
R10316 VSS VSS.n97 0.00545413
R10317 VSS VSS.n100 0.00545413
R10318 VSS.n103 VSS 0.00545413
R10319 VSS VSS.n85 0.00545413
R10320 VSS VSS.n88 0.00545413
R10321 VSS.n91 VSS 0.00545413
R10322 VSS.n3345 VSS 0.00545413
R10323 VSS.n3343 VSS 0.00545413
R10324 VSS.n3341 VSS 0.00545413
R10325 VSS.n3282 VSS 0.00545413
R10326 VSS VSS.n3285 0.00545413
R10327 VSS.n3287 VSS 0.00545413
R10328 VSS.n57 VSS 0.00545413
R10329 VSS.n60 VSS 0.00545413
R10330 VSS.n63 VSS 0.00545413
R10331 VSS.n274 VSS 0.00545413
R10332 VSS.n272 VSS 0.00545413
R10333 VSS.n270 VSS 0.00545413
R10334 VSS.n1031 VSS 0.00545413
R10335 VSS.n1033 VSS 0.00545413
R10336 VSS.n1053 VSS 0.00545413
R10337 VSS.n2520 VSS 0.00545413
R10338 VSS.n2523 VSS 0.00545413
R10339 VSS.n2531 VSS 0.00545413
R10340 VSS.n2539 VSS 0.00545413
R10341 VSS.n1036 VSS 0.00545413
R10342 VSS.n1044 VSS 0.00545413
R10343 VSS VSS.n1042 0.00545413
R10344 VSS.n993 VSS 0.00545413
R10345 VSS.n991 VSS 0.00545413
R10346 VSS.n989 VSS 0.00545413
R10347 VSS.n2478 VSS 0.00545413
R10348 VSS.n2480 VSS 0.00545413
R10349 VSS.n2482 VSS 0.00545413
R10350 VSS.n920 VSS 0.00545413
R10351 VSS.n923 VSS 0.00545413
R10352 VSS.n926 VSS 0.00545413
R10353 VSS.n933 VSS 0.00545413
R10354 VSS.n935 VSS 0.00545413
R10355 VSS.n937 VSS 0.00545413
R10356 VSS.n1018 VSS 0.00545413
R10357 VSS.n1020 VSS 0.00545413
R10358 VSS.n1026 VSS 0.00545413
R10359 VSS.n3005 VSS 0.00545413
R10360 VSS.n3003 VSS 0.00545413
R10361 VSS.n3001 VSS 0.00545413
R10362 VSS.n44 VSS 0.00545413
R10363 VSS.n42 VSS 0.00545413
R10364 VSS.n40 VSS 0.00545413
R10365 VSS.n3463 VSS 0.00545413
R10366 VSS VSS.n3461 0.00545413
R10367 VSS VSS.n3459 0.00545413
R10368 VSS.n465 VSS 0.00545413
R10369 VSS VSS.n468 0.00545413
R10370 VSS.n470 VSS 0.00545413
R10371 VSS VSS.n481 0.00545413
R10372 VSS VSS.n484 0.00545413
R10373 VSS.n487 VSS 0.00545413
R10374 VSS VSS.n450 0.00545413
R10375 VSS VSS.n453 0.00545413
R10376 VSS.n455 VSS 0.00545413
R10377 VSS.n431 VSS 0.00545413
R10378 VSS VSS.n434 0.00545413
R10379 VSS.n436 VSS 0.00545413
R10380 VSS.n2982 VSS 0.00545413
R10381 VSS.n2985 VSS 0.00545413
R10382 VSS.n2988 VSS 0.00545413
R10383 VSS.n2550 VSS 0.00545413
R10384 VSS VSS.n2548 0.00545413
R10385 VSS VSS.n2546 0.00545413
R10386 VSS VSS.n1373 0.00545413
R10387 VSS VSS.n1376 0.00545413
R10388 VSS.n1379 VSS 0.00545413
R10389 VSS VSS.n2321 0.00545413
R10390 VSS VSS.n2324 0.00545413
R10391 VSS.n2327 VSS 0.00545413
R10392 VSS.n1967 VSS 0.00545413
R10393 VSS.n1965 VSS 0.00545413
R10394 VSS.n1963 VSS 0.00545413
R10395 VSS.n2243 VSS 0.00545413
R10396 VSS.n2241 VSS 0.00545413
R10397 VSS.n2239 VSS 0.00545413
R10398 VSS.n2264 VSS 0.00545413
R10399 VSS VSS.n2274 0.00545413
R10400 VSS VSS.n2313 0.00545413
R10401 VSS.n2338 VSS 0.00545413
R10402 VSS.n2352 VSS 0.00545413
R10403 VSS VSS.n2362 0.00545413
R10404 VSS.n2372 VSS 0.00545413
R10405 VSS VSS.n1069 0.00545413
R10406 VSS VSS.n2132 0.00545413
R10407 VSS VSS.n2135 0.00545413
R10408 VSS.n2138 VSS 0.00545413
R10409 VSS VSS.n2088 0.00545413
R10410 VSS VSS.n2091 0.00545413
R10411 VSS.n2094 VSS 0.00545413
R10412 VSS.n2073 VSS 0.00545413
R10413 VSS VSS.n2076 0.00545413
R10414 VSS.n2078 VSS 0.00545413
R10415 VSS.n2020 VSS 0.00545413
R10416 VSS.n2018 VSS 0.00545413
R10417 VSS.n2016 VSS 0.00545413
R10418 VSS.n2212 VSS 0.00545413
R10419 VSS.n2210 VSS 0.00545413
R10420 VSS.n2203 VSS 0.00545413
R10421 VSS.n2201 VSS 0.00545413
R10422 VSS.n2194 VSS 0.00545413
R10423 VSS.n2192 VSS 0.00545413
R10424 VSS.n2185 VSS 0.00545413
R10425 VSS.n2183 VSS 0.00545413
R10426 VSS.n2389 VSS 0.00545413
R10427 VSS.n2392 VSS 0.00545413
R10428 VSS.n2395 VSS 0.00545413
R10429 VSS.n1340 VSS 0.00545413
R10430 VSS.n1342 VSS 0.00545413
R10431 VSS.n1344 VSS 0.00545413
R10432 VSS.n1331 VSS 0.00545413
R10433 VSS.n1335 VSS 0.00545413
R10434 VSS.n1938 VSS 0.00545413
R10435 VSS VSS.n1936 0.00545413
R10436 VSS.n1824 VSS 0.00545413
R10437 VSS.n1822 VSS 0.00545413
R10438 VSS.n1820 VSS 0.00545413
R10439 VSS VSS.n1804 0.00545413
R10440 VSS VSS.n1807 0.00545413
R10441 VSS.n1810 VSS 0.00545413
R10442 VSS.n2631 VSS 0.00545413
R10443 VSS.n2634 VSS 0.00545413
R10444 VSS.n2637 VSS 0.00545413
R10445 VSS.n1635 VSS 0.00545413
R10446 VSS.n1637 VSS 0.00545413
R10447 VSS.n1639 VSS 0.00545413
R10448 VSS.n1621 VSS 0.00545413
R10449 VSS.n1623 VSS 0.00545413
R10450 VSS.n1625 VSS 0.00545413
R10451 VSS.n1580 VSS 0.00545413
R10452 VSS.n1582 VSS 0.00545413
R10453 VSS.n1584 VSS 0.00545413
R10454 VSS VSS.n1594 0.00545413
R10455 VSS.n1561 VSS 0.00545413
R10456 VSS.n1570 VSS 0.00545413
R10457 VSS VSS.n1568 0.00545413
R10458 VSS.n794 VSS 0.00545413
R10459 VSS.n799 VSS 0.00545413
R10460 VSS.n819 VSS 0.00545413
R10461 VSS VSS.n817 0.00545413
R10462 VSS.n1872 VSS 0.00545413
R10463 VSS.n1875 VSS 0.00545413
R10464 VSS.n1878 VSS 0.00545413
R10465 VSS.n2659 VSS.n2658 0.004773
R10466 VSS.n2830 VSS.n2829 0.00438534
R10467 VSS.n2832 VSS.n2830 0.00438534
R10468 VSS.n542 VSS 0.00432979
R10469 VSS.n546 VSS 0.00432979
R10470 VSS.n549 VSS 0.00432979
R10471 VSS.n560 VSS 0.00432979
R10472 VSS.n564 VSS 0.00432979
R10473 VSS.n567 VSS 0.00432979
R10474 VSS.n3215 VSS 0.00427778
R10475 VSS.n827 VSS 0.00427622
R10476 VSS.n830 VSS 0.00427622
R10477 VSS.n833 VSS 0.00427622
R10478 VSS.n578 VSS 0.00425
R10479 VSS.n581 VSS 0.00425
R10480 VSS.n584 VSS 0.00425
R10481 VSS.n880 VSS 0.00425
R10482 VSS.n883 VSS 0.00425
R10483 VSS.n886 VSS 0.00425
R10484 VSS.n1849 VSS 0.00425
R10485 VSS.n1852 VSS 0.00425
R10486 VSS VSS.n1864 0.00425
R10487 VSS VSS.n1469 0.00425
R10488 VSS.n843 VSS 0.00422414
R10489 VSS.n846 VSS 0.00422414
R10490 VSS.n849 VSS 0.00422414
R10491 VSS.n527 VSS 0.00417347
R10492 VSS.n530 VSS 0.00417347
R10493 VSS.n533 VSS 0.00417347
R10494 VSS.n662 VSS 0.00417347
R10495 VSS.n660 VSS 0.00417347
R10496 VSS VSS.n2804 0.00417347
R10497 VSS VSS.n2806 0.00417347
R10498 VSS.n2697 VSS 0.00417347
R10499 VSS VSS.n2695 0.00417347
R10500 VSS VSS.n2693 0.00417347
R10501 VSS.n2921 VSS.n328 0.00413112
R10502 VSS.n3453 VSS.n29 0.00410721
R10503 VSS VSS.n1147 0.00405263
R10504 VSS VSS.n1155 0.00405263
R10505 VSS VSS.n1137 0.00405263
R10506 VSS.n1183 VSS 0.00405263
R10507 VSS.n1194 VSS 0.00405263
R10508 VSS.n2663 VSS.n2662 0.00397181
R10509 VSS.n872 VSS 0.00380275
R10510 VSS.n905 VSS 0.00380275
R10511 VSS VSS.n1486 0.00380275
R10512 VSS.n1529 VSS 0.00380275
R10513 VSS.n1474 VSS 0.00380275
R10514 VSS VSS.n1496 0.00380275
R10515 VSS.n1224 VSS 0.00380275
R10516 VSS.n1988 VSS 0.00380275
R10517 VSS.n1992 VSS 0.00380275
R10518 VSS.n1996 VSS 0.00380275
R10519 VSS VSS.n1103 0.00380275
R10520 VSS.n2303 VSS 0.00380275
R10521 VSS.n2052 VSS 0.00380275
R10522 VSS VSS.n2269 0.00380275
R10523 VSS.n2271 VSS 0.00380275
R10524 VSS.n2283 VSS 0.00380275
R10525 VSS.n2310 VSS 0.00380275
R10526 VSS VSS.n2357 0.00380275
R10527 VSS.n2359 VSS 0.00380275
R10528 VSS.n1433 VSS 0.00380275
R10529 VSS VSS.n1303 0.00380275
R10530 VSS.n1263 VSS 0.00380275
R10531 VSS.n1267 VSS 0.00380275
R10532 VSS.n1271 VSS 0.00380275
R10533 VSS.n1319 VSS 0.00380275
R10534 VSS.n1948 VSS 0.00380275
R10535 VSS.n1286 VSS 0.00380275
R10536 VSS VSS.n1289 0.00380275
R10537 VSS.n1458 VSS 0.00380275
R10538 VSS.n1456 VSS 0.00380275
R10539 VSS.n1449 VSS 0.00380275
R10540 VSS.n1447 VSS 0.00380275
R10541 VSS.n3050 VSS 0.00380275
R10542 VSS.n1015 VSS 0.00380275
R10543 VSS VSS.n2456 0.00380275
R10544 VSS.n2475 VSS 0.00380275
R10545 VSS.n3321 VSS 0.00380275
R10546 VSS.n94 VSS 0.00380275
R10547 VSS VSS.n82 0.00380275
R10548 VSS.n3347 VSS 0.00380275
R10549 VSS.n3280 VSS 0.00380275
R10550 VSS.n3303 VSS 0.00380275
R10551 VSS VSS.n66 0.00380275
R10552 VSS.n263 VSS 0.00380275
R10553 VSS.n2512 VSS 0.00380275
R10554 VSS.n1051 VSS 0.00380275
R10555 VSS.n2525 VSS 0.00380275
R10556 VSS VSS.n2528 0.00380275
R10557 VSS.n2537 VSS 0.00380275
R10558 VSS.n2535 VSS 0.00380275
R10559 VSS.n1040 VSS 0.00380275
R10560 VSS VSS.n995 0.00380275
R10561 VSS.n2484 VSS 0.00380275
R10562 VSS.n2436 VSS 0.00380275
R10563 VSS.n2440 VSS 0.00380275
R10564 VSS VSS.n2431 0.00380275
R10565 VSS.n1392 VSS 0.00380275
R10566 VSS VSS.n1403 0.00380275
R10567 VSS VSS.n1398 0.00380275
R10568 VSS.n2579 VSS 0.00380275
R10569 VSS.n929 VSS 0.00380275
R10570 VSS.n940 VSS 0.00380275
R10571 VSS.n1024 VSS 0.00380275
R10572 VSS.n2994 VSS 0.00380275
R10573 VSS VSS.n46 0.00380275
R10574 VSS.n3457 VSS 0.00380275
R10575 VSS.n463 VSS 0.00380275
R10576 VSS.n398 VSS 0.00380275
R10577 VSS.n478 VSS 0.00380275
R10578 VSS.n644 VSS 0.00380275
R10579 VSS.n447 VSS 0.00380275
R10580 VSS.n429 VSS 0.00380275
R10581 VSS.n602 VSS 0.00380275
R10582 VSS.n679 VSS 0.00380275
R10583 VSS.n2990 VSS 0.00380275
R10584 VSS.n3153 VSS 0.00380275
R10585 VSS.n1424 VSS 0.00380275
R10586 VSS VSS.n1429 0.00380275
R10587 VSS.n1370 VSS 0.00380275
R10588 VSS.n2318 VSS 0.00380275
R10589 VSS VSS.n1969 0.00380275
R10590 VSS VSS.n2245 0.00380275
R10591 VSS.n2260 VSS 0.00380275
R10592 VSS.n2266 VSS 0.00380275
R10593 VSS.n2278 VSS 0.00380275
R10594 VSS.n2280 VSS 0.00380275
R10595 VSS.n2348 VSS 0.00380275
R10596 VSS.n2354 VSS 0.00380275
R10597 VSS.n2366 VSS 0.00380275
R10598 VSS.n2374 VSS 0.00380275
R10599 VSS.n2152 VSS 0.00380275
R10600 VSS VSS.n2163 0.00380275
R10601 VSS VSS.n2159 0.00380275
R10602 VSS.n2129 VSS 0.00380275
R10603 VSS.n2085 VSS 0.00380275
R10604 VSS.n2071 VSS 0.00380275
R10605 VSS VSS.n2022 0.00380275
R10606 VSS VSS.n2216 0.00380275
R10607 VSS VSS.n2214 0.00380275
R10608 VSS VSS.n2207 0.00380275
R10609 VSS VSS.n2205 0.00380275
R10610 VSS VSS.n2198 0.00380275
R10611 VSS VSS.n2196 0.00380275
R10612 VSS VSS.n2189 0.00380275
R10613 VSS VSS.n2187 0.00380275
R10614 VSS.n2398 VSS 0.00380275
R10615 VSS.n1912 VSS 0.00380275
R10616 VSS.n1234 VSS 0.00380275
R10617 VSS VSS.n1346 0.00380275
R10618 VSS VSS.n1338 0.00380275
R10619 VSS.n1351 VSS 0.00380275
R10620 VSS.n1934 VSS 0.00380275
R10621 VSS.n1932 VSS 0.00380275
R10622 VSS VSS.n1507 0.00380275
R10623 VSS.n1801 VSS 0.00380275
R10624 VSS VSS.n2640 0.00380275
R10625 VSS.n1649 VSS 0.00380275
R10626 VSS VSS.n1627 0.00380275
R10627 VSS.n1586 VSS 0.00380275
R10628 VSS.n1615 VSS 0.00380275
R10629 VSS.n1613 VSS 0.00380275
R10630 VSS VSS.n1608 0.00380275
R10631 VSS.n1673 VSS 0.00380275
R10632 VSS.n1670 VSS 0.00380275
R10633 VSS VSS.n784 0.00380275
R10634 VSS VSS.n1630 0.00380275
R10635 VSS VSS.n804 0.00380275
R10636 VSS VSS.n1642 0.00380275
R10637 VSS VSS.n2643 0.00380275
R10638 VSS VSS.n2646 0.00380275
R10639 VSS.n1881 VSS 0.00380275
R10640 VSS VSS.n3416 0.00367647
R10641 VSS.n3418 VSS 0.00367647
R10642 VSS.n2610 VSS 0.00352521
R10643 VSS.n2004 VSS 0.00352521
R10644 VSS.n1278 VSS 0.00352521
R10645 VSS VSS.n3327 0.00352521
R10646 VSS VSS.n3309 0.00352521
R10647 VSS.n2515 VSS 0.00352521
R10648 VSS VSS.n2419 0.00352521
R10649 VSS.n1418 VSS 0.00352521
R10650 VSS.n2582 VSS 0.00352521
R10651 VSS.n652 VSS 0.00352521
R10652 VSS.n406 VSS 0.00352521
R10653 VSS VSS.n615 0.00352521
R10654 VSS.n3213 VSS 0.00352521
R10655 VSS.n2178 VSS 0.00352521
R10656 VSS.n1920 VSS 0.00352521
R10657 VSS VSS.n1892 0.00352521
R10658 VSS VSS.n1598 0.00352521
R10659 VSS.n1537 VSS 0.00352521
R10660 VSS.n695 VSS 0.0035
R10661 VSS.n2656 VSS 0.0035
R10662 VSS VSS.n2568 0.00335714
R10663 VSS VSS.n2566 0.00335714
R10664 VSS VSS.n2559 0.00335714
R10665 VSS VSS.n2557 0.00335714
R10666 VSS.n664 VSS.n497 0.00324928
R10667 VSS.n899 VSS.n878 0.00324928
R10668 VSS.n2834 VSS.n2833 0.00322504
R10669 VSS.n3431 VSS 0.0031087
R10670 VSS VSS.n3445 0.0031087
R10671 VSS VSS.n3137 0.00309615
R10672 VSS.n3139 VSS 0.00309615
R10673 VSS VSS.n3149 0.00308373
R10674 VSS VSS.n3147 0.00308373
R10675 VSS VSS.n552 0.00305319
R10676 VSS VSS.n570 0.00305319
R10677 VSS.n2501 VSS 0.00303521
R10678 VSS.n2499 VSS 0.00303521
R10679 VSS VSS.n676 0.00301748
R10680 VSS.n836 VSS 0.00301748
R10681 VSS VSS.n901 0.00301748
R10682 VSS.n586 VSS 0.003
R10683 VSS VSS.n889 0.003
R10684 VSS VSS.n1855 0.003
R10685 VSS.n1857 VSS 0.003
R10686 VSS.n1467 VSS 0.003
R10687 VSS VSS.n1885 0.003
R10688 VSS.n1697 VSS.n1696 0.00298619
R10689 VSS.n852 VSS 0.00298276
R10690 VSS.n536 VSS 0.00294898
R10691 VSS.n2691 VSS 0.00294898
R10692 VSS.n3481 VSS 0.00293243
R10693 VSS.n3479 VSS 0.00293243
R10694 VSS VSS.n1708 0.00293243
R10695 VSS.n1716 VSS 0.00293243
R10696 VSS.n3103 VSS 0.00286842
R10697 VSS VSS.n3104 0.00286842
R10698 VSS.n716 VSS.n715 0.00279385
R10699 VSS.n3111 VSS 0.00279299
R10700 VSS VSS.n3112 0.00279299
R10701 VSS.n3175 VSS 0.00261765
R10702 VSS.n3177 VSS 0.00261765
R10703 VSS.n136 VSS 0.00258494
R10704 VSS VSS.n3353 0.00258494
R10705 VSS VSS.n3364 0.00258494
R10706 VSS.n3366 VSS 0.00258494
R10707 VSS.n3374 VSS 0.00258494
R10708 VSS VSS.n3393 0.00258494
R10709 VSS.n3403 VSS 0.00258494
R10710 VSS VSS.n3407 0.00258494
R10711 VSS VSS.n600 0.00258494
R10712 VSS VSS.n669 0.00258494
R10713 VSS.n1162 VSS 0.00247368
R10714 VSS.n1190 VSS 0.00247368
R10715 VSS.n2564 VSS 0.00240476
R10716 VSS.n2562 VSS 0.00240476
R10717 VSS VSS.n3126 0.00240476
R10718 VSS.n3128 VSS 0.00240476
R10719 VSS VSS.n2410 0.00240141
R10720 VSS.n3207 VSS 0.00240141
R10721 VSS VSS.n3200 0.00240141
R10722 VSS VSS.n3198 0.00240141
R10723 VSS.n3193 VSS 0.00240141
R10724 VSS VSS.n3191 0.00240141
R10725 VSS VSS.n3184 0.00240141
R10726 VSS VSS.n3182 0.00240141
R10727 VSS.n666 VSS 0.00233673
R10728 VSS.n876 VSS 0.00233673
R10729 VSS VSS.n3435 0.00223913
R10730 VSS VSS.n3433 0.00223913
R10731 VSS.n3123 VSS 0.00223077
R10732 VSS.n3131 VSS 0.00223077
R10733 VSS.n3145 VSS 0.00222249
R10734 VSS.n3426 VSS 0.00222249
R10735 VSS.n892 VSS 0.00219811
R10736 VSS.n908 VSS 0.00219811
R10737 VSS.n2613 VSS 0.00219811
R10738 VSS.n859 VSS 0.00219811
R10739 VSS VSS.n1485 0.00219811
R10740 VSS.n1867 VSS 0.00219811
R10741 VSS.n1239 VSS 0.00219811
R10742 VSS.n821 VSS 0.00219811
R10743 VSS.n838 VSS 0.00219811
R10744 VSS VSS.n1495 0.00219811
R10745 VSS VSS.n1232 0.00219811
R10746 VSS VSS.n1990 0.00219811
R10747 VSS VSS.n1994 0.00219811
R10748 VSS VSS.n1998 0.00219811
R10749 VSS VSS.n2000 0.00219811
R10750 VSS VSS.n2002 0.00219811
R10751 VSS.n2290 VSS 0.00219811
R10752 VSS VSS.n2306 0.00219811
R10753 VSS.n2384 VSS 0.00219811
R10754 VSS VSS.n1323 0.00219811
R10755 VSS.n1306 VSS 0.00219811
R10756 VSS VSS.n1265 0.00219811
R10757 VSS VSS.n1269 0.00219811
R10758 VSS.n1273 VSS 0.00219811
R10759 VSS.n1256 VSS 0.00219811
R10760 VSS.n1254 VSS 0.00219811
R10761 VSS.n1352 VSS 0.00219811
R10762 VSS VSS.n3059 0.00219811
R10763 VSS VSS.n3021 0.00219811
R10764 VSS.n1062 VSS 0.00219811
R10765 VSS.n2461 VSS 0.00219811
R10766 VSS.n2477 VSS 0.00219811
R10767 VSS VSS.n3410 0.00219811
R10768 VSS.n3331 VSS 0.00219811
R10769 VSS.n3386 VSS 0.00219811
R10770 VSS.n3382 VSS 0.00219811
R10771 VSS.n3291 VSS 0.00219811
R10772 VSS VSS.n123 0.00219811
R10773 VSS.n3313 VSS 0.00219811
R10774 VSS VSS.n3423 0.00219811
R10775 VSS.n3157 VSS 0.00219811
R10776 VSS.n975 VSS 0.00219811
R10777 VSS.n1035 VSS 0.00219811
R10778 VSS.n3162 VSS 0.00219811
R10779 VSS VSS.n3170 0.00219811
R10780 VSS.n2508 VSS 0.00219811
R10781 VSS VSS.n2438 0.00219811
R10782 VSS.n2442 VSS 0.00219811
R10783 VSS.n2428 VSS 0.00219811
R10784 VSS.n2425 VSS 0.00219811
R10785 VSS.n2422 VSS 0.00219811
R10786 VSS.n1405 VSS 0.00219811
R10787 VSS.n1414 VSS 0.00219811
R10788 VSS VSS.n1410 0.00219811
R10789 VSS.n1396 VSS 0.00219811
R10790 VSS.n1401 VSS 0.00219811
R10791 VSS.n2576 VSS 0.00219811
R10792 VSS.n931 VSS 0.00219811
R10793 VSS.n1173 VSS 0.00219811
R10794 VSS.n966 VSS 0.00219811
R10795 VSS.n3011 VSS 0.00219811
R10796 VSS.n3439 VSS 0.00219811
R10797 VSS.n508 VSS 0.00219811
R10798 VSS.n555 VSS 0.00219811
R10799 VSS.n460 VSS 0.00219811
R10800 VSS VSS.n474 0.00219811
R10801 VSS.n649 VSS 0.00219811
R10802 VSS.n403 VSS 0.00219811
R10803 VSS.n443 VSS 0.00219811
R10804 VSS.n426 VSS 0.00219811
R10805 VSS VSS.n689 0.00219811
R10806 VSS.n683 VSS 0.00219811
R10807 VSS.n637 VSS 0.00219811
R10808 VSS.n621 VSS 0.00219811
R10809 VSS.n611 VSS 0.00219811
R10810 VSS VSS.n3483 0.00219811
R10811 VSS VSS.n1422 0.00219811
R10812 VSS.n1367 VSS 0.00219811
R10813 VSS VSS.n2333 0.00219811
R10814 VSS.n2233 VSS 0.00219811
R10815 VSS.n2250 VSS 0.00219811
R10816 VSS.n2165 VSS 0.00219811
R10817 VSS.n2161 VSS 0.00219811
R10818 VSS.n2157 VSS 0.00219811
R10819 VSS VSS.n2170 0.00219811
R10820 VSS.n2174 VSS 0.00219811
R10821 VSS.n2126 VSS 0.00219811
R10822 VSS.n2082 VSS 0.00219811
R10823 VSS.n2035 VSS 0.00219811
R10824 VSS.n2219 VSS 0.00219811
R10825 VSS.n2180 VSS 0.00219811
R10826 VSS.n1917 VSS 0.00219811
R10827 VSS.n1896 VSS 0.00219811
R10828 VSS VSS.n1929 0.00219811
R10829 VSS VSS.n1523 0.00219811
R10830 VSS VSS.n1514 0.00219811
R10831 VSS.n1706 VSS 0.00219811
R10832 VSS.n1686 VSS 0.00219811
R10833 VSS VSS.n895 0.00219811
R10834 VSS.n2649 VSS 0.00219811
R10835 VSS VSS.n1646 0.00219811
R10836 VSS.n1634 VSS 0.00219811
R10837 VSS VSS.n1666 0.00219811
R10838 VSS.n1617 VSS 0.00219811
R10839 VSS.n1610 VSS 0.00219811
R10840 VSS.n1606 VSS 0.00219811
R10841 VSS.n1604 VSS 0.00219811
R10842 VSS.n1601 VSS 0.00219811
R10843 VSS.n1534 VSS 0.00219811
R10844 VSS.n331 VSS 0.00219811
R10845 VSS VSS.n2505 0.00219014
R10846 VSS VSS.n2503 0.00219014
R10847 VSS VSS.n3239 0.00215138
R10848 VSS VSS.n3247 0.00215138
R10849 VSS VSS.n3255 0.00215138
R10850 VSS.n3265 VSS 0.00215138
R10851 VSS VSS.n1691 0.00215138
R10852 VSS VSS.n1 0.00215138
R10853 VSS.n720 VSS.n719 0.00211919
R10854 VSS VSS.n1685 0.00210237
R10855 VSS VSS.n1682 0.00210237
R10856 VSS VSS.n2686 0.00210237
R10857 VSS VSS.n2684 0.00210237
R10858 VSS VSS.n2674 0.00210237
R10859 VSS VSS.n2671 0.00210237
R10860 VSS VSS.n2661 0.00210237
R10861 VSS VSS.n2659 0.00210237
R10862 VSS VSS.n955 0.0020562
R10863 VSS VSS.n953 0.0020562
R10864 VSS.n2924 VSS 0.0020562
R10865 VSS.n2927 VSS 0.0020562
R10866 VSS.n3324 VSS 0.00191732
R10867 VSS.n3306 VSS 0.00191732
R10868 VSS VSS.n2518 0.00191732
R10869 VSS.n2585 VSS 0.00191732
R10870 VSS.n670 VSS 0.00191732
R10871 VSS.n409 VSS 0.00191732
R10872 VSS VSS.n1926 0.00191732
R10873 VSS.n1889 VSS 0.00191732
R10874 VSS VSS.n1543 0.00191732
R10875 VSS.n131 VSS 0.00188996
R10876 VSS.n138 VSS 0.00188996
R10877 VSS.n3358 VSS 0.00188996
R10878 VSS.n3361 VSS 0.00188996
R10879 VSS VSS.n3378 0.00188996
R10880 VSS VSS.n3376 0.00188996
R10881 VSS.n3398 VSS 0.00188996
R10882 VSS.n3401 VSS 0.00188996
R10883 VSS.n595 VSS 0.00188996
R10884 VSS.n598 VSS 0.00188996
R10885 VSS.n1742 VSS 0.00184663
R10886 VSS VSS.n1747 0.00184663
R10887 VSS.n1758 VSS 0.00184663
R10888 VSS VSS.n1764 0.00184663
R10889 VSS VSS.n1779 0.00184328
R10890 VSS.n1781 VSS 0.00184328
R10891 VSS.n1792 VSS 0.00184328
R10892 VSS VSS.n911 0.00184328
R10893 VSS.n3205 VSS 0.00176761
R10894 VSS.n3203 VSS 0.00176761
R10895 VSS.n3196 VSS 0.00176761
R10896 VSS VSS.n250 0.00176761
R10897 VSS.n3189 VSS 0.00176761
R10898 VSS.n3187 VSS 0.00176761
R10899 VSS.n3180 VSS 0.00176761
R10900 VSS.n3413 VSS 0.00176761
R10901 VSS VSS.n3477 0.00171622
R10902 VSS VSS.n3475 0.00171622
R10903 VSS VSS.n1714 0.00171622
R10904 VSS VSS.n1712 0.00171622
R10905 VSS VSS.n3086 0.00168421
R10906 VSS.n291 VSS 0.00168421
R10907 VSS.n3105 VSS 0.00168421
R10908 VSS.n2377 VSS 0.00165385
R10909 VSS VSS.n2405 0.00165385
R10910 VSS.n294 VSS 0.0016465
R10911 VSS.n3113 VSS 0.0016465
R10912 VSS VSS.n3045 0.00158216
R10913 VSS VSS.n3043 0.00158216
R10914 VSS VSS.n3070 0.00158216
R10915 VSS VSS.n3068 0.00158216
R10916 VSS.n15 VSS 0.00158
R10917 VSS.n17 VSS 0.00158
R10918 VSS.n496 VSS 0.00157463
R10919 VSS.n2654 VSS 0.00157143
R10920 VSS.n1679 VSS 0.00156825
R10921 VSS.n1676 VSS 0.00156825
R10922 VSS.n2681 VSS 0.00156825
R10923 VSS.n2678 VSS 0.00156825
R10924 VSS.n2668 VSS 0.00156825
R10925 VSS.n2665 VSS 0.00156825
R10926 VSS.n951 VSS 0.00153746
R10927 VSS.n949 VSS 0.00153746
R10928 VSS.n2929 VSS 0.00153746
R10929 VSS VSS.n2934 0.00153746
R10930 VSS VSS.n3485 0.0015
R10931 VSS.n1703 VSS 0.0015
R10932 VSS VSS.n753 0.00149815
R10933 VSS VSS.n751 0.00149815
R10934 VSS.n2 VSS 0.00149448
R10935 VSS.n3487 VSS 0.00149448
R10936 VSS.n1701 VSS 0.00149448
R10937 VSS.n1697 VSS 0.00149448
R10938 VSS.n1737 VSS 0.00139776
R10939 VSS.n1740 VSS 0.00139776
R10940 VSS.n1752 VSS 0.00139776
R10941 VSS.n1756 VSS 0.00139776
R10942 VSS.n1770 VSS 0.00139552
R10943 VSS.n1776 VSS 0.00139552
R10944 VSS VSS.n1796 0.00139552
R10945 VSS VSS.n1794 0.00139552
R10946 VSS VSS.n573 0.00136539
R10947 VSS VSS.n854 0.00136539
R10948 VSS VSS.n231 0.00132569
R10949 VSS VSS.n317 0.00132569
R10950 VSS VSS.n226 0.00132569
R10951 VSS.n3220 VSS 0.00132569
R10952 VSS.n3218 VSS 0.00132569
R10953 VSS.n740 VSS 0.00130959
R10954 VSS VSS.n739 0.00130959
R10955 VSS.n736 VSS 0.00130959
R10956 VSS VSS.n735 0.00130959
R10957 VSS.n722 VSS 0.00130959
R10958 VSS VSS.n721 0.00130959
R10959 VSS.n718 VSS 0.00130959
R10960 VSS VSS.n717 0.00130959
R10961 VSS.n703 VSS 0.00130959
R10962 VSS VSS.n702 0.00130959
R10963 VSS.n699 VSS 0.00130959
R10964 VSS VSS.n698 0.00130959
R10965 VSS VSS.n2608 0.0013
R10966 VSS.n618 VSS 0.0013
R10967 VSS.n2603 VSS.n862 0.00129295
R10968 VSS VSS.n862 0.00129295
R10969 VSS.n631 VSS.n630 0.00129295
R10970 VSS.n630 VSS 0.00129295
R10971 VSS.n2413 VSS 0.0012563
R10972 VSS.n3268 VSS 0.0012563
R10973 VSS.n3253 VSS 0.0012563
R10974 VSS.n3245 VSS 0.0012563
R10975 VSS.n3235 VSS 0.0012563
R10976 VSS.n3243 VSS 0.0012563
R10977 VSS.n3251 VSS 0.0012563
R10978 VSS VSS.n3258 0.0012563
R10979 VSS.n3262 VSS 0.0012563
R10980 VSS VSS.n319 0.00124689
R10981 VSS VSS.n3072 0.0012438
R10982 VSS.n3038 VSS 0.00122144
R10983 VSS VSS.n3453 0.00122144
R10984 VSS.n3065 VSS 0.00122144
R10985 VSS.n3063 VSS 0.00122144
R10986 VSS VSS.n3024 0.00122
R10987 VSS VSS.n3030 0.00122
R10988 VSS.n3078 VSS 0.00118965
R10989 VSS VSS.n3092 0.00111785
R10990 VSS VSS.n3100 0.00111785
R10991 VSS VSS.n3108 0.00111785
R10992 VSS VSS.n3116 0.00111785
R10993 VSS.n3447 VSS 0.00111644
R10994 VSS VSS.n339 0.00103973
R10995 VSS.n747 VSS 0.00103973
R10996 VSS.n746 VSS 0.00103973
R10997 VSS VSS.n743 0.00103973
R10998 VSS.n731 VSS 0.00103973
R10999 VSS VSS.n730 0.00103973
R11000 VSS.n727 VSS 0.00103973
R11001 VSS VSS.n726 0.00103973
R11002 VSS.n713 VSS 0.00103973
R11003 VSS VSS.n710 0.00103973
R11004 VSS.n709 VSS 0.00103973
R11005 VSS VSS.n706 0.00103973
R11006 VSS.n1427 VSS.t501 0.00101932
R11007 VSS.n308 VSS 0.000983871
R11008 VSS.n3089 VSS 0.000954545
R11009 VSS VSS.n304 0.000945545
R11010 VSS.n3097 VSS 0.000945545
R11011 VSS.n233 VSS 0.000944444
R11012 VSS.n2604 VSS.n2603 0.000896476
R11013 VSS.n631 VSS.n625 0.000896476
R11014 VSS VSS.n1146 0.000894737
R11015 VSS VSS.n1154 0.000894737
R11016 VSS.n1163 VSS 0.000894737
R11017 VSS.n1138 VSS 0.000894737
R11018 VSS.n1184 VSS 0.000894737
R11019 VSS.n1191 VSS 0.000894737
R11020 VSS.n1195 VSS 0.000894737
R11021 VSS.n2940 VSS 0.000799003
R11022 VSS.n2945 VSS 0.000799003
R11023 VSS.n2948 VSS 0.000799003
R11024 VSS.n2952 VSS 0.000799003
R11025 VSS.n2957 VSS 0.000799003
R11026 VSS.n2961 VSS 0.000799003
R11027 VSS.n2963 VSS 0.000799003
R11028 VSS VSS.n3075 0.000799003
R11029 VSS.n3092 VSS.n305 0.00070595
R11030 VSS.n3094 VSS.n3093 0.00070595
R11031 VSS.n3096 VSS.n3095 0.00070595
R11032 VSS.n3100 VSS.n290 0.00070595
R11033 VSS.n3102 VSS.n3101 0.00070595
R11034 VSS.n3104 VSS.n3103 0.00070595
R11035 VSS.n3108 VSS.n289 0.00070595
R11036 VSS.n3110 VSS.n3109 0.00070595
R11037 VSS.n3112 VSS.n3111 0.00070595
R11038 VSS.n3116 VSS.n288 0.00070595
R11039 VSS.n3118 VSS.n3117 0.00070595
R11040 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n2 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t6 36.935
R11041 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n9 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t5 36.935
R11042 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n8 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t15 36.935
R11043 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n3 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t12 31.528
R11044 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n5 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t10 31.528
R11045 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n6 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t4 31.528
R11046 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n11 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t8 25.5364
R11047 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n2 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t9 18.1962
R11048 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n9 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t7 18.1962
R11049 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n8 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t3 18.1962
R11050 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n3 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t14 15.3826
R11051 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n5 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t13 15.3826
R11052 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n6 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t11 15.3826
R11053 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n11 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t2 14.0749
R11054 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n6 7.63631
R11055 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n3 6.86134
R11056 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n7 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 6.23913
R11057 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n5 8.03067
R11058 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n4 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 5.01116
R11059 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n0 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 4.5005
R11060 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n10 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 3.25197
R11061 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n7 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 2.91397
R11062 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n1 2.52047
R11063 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n12 2.3025
R11064 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n10 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 2.25107
R11065 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 2.24713
R11066 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n2 2.13398
R11067 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n8 2.12175
R11068 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n9 2.12075
R11069 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n0 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n7 1.69271
R11070 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n11 1.42706
R11071 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n12 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n4 1.32654
R11072 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n4 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 1.12056
R11073 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n0 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n10 1.02402
R11074 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n12 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n0 0.557773
R11075 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.n2 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.t8 36.935
R11076 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.n3 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.t5 31.4332
R11077 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.n5 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.t4 29.8135
R11078 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.n5 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.t3 27.8352
R11079 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.n2 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.t6 18.1962
R11080 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.n3 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.t7 15.3826
R11081 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.t2 7.09905
R11082 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.n3 6.86029
R11083 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.n4 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 5.01077
R11084 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.n6 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 3.41843
R11085 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.n1 3.25053
R11086 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.n1 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.t0 2.2755
R11087 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.n1 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.n0 2.2755
R11088 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.n6 2.2505
R11089 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.n2 2.13459
R11090 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.n5 1.74998
R11091 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.n6 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.n4 1.50381
R11092 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.n4 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 1.12067
R11093 VDD99.n286 VDD99.t341 2529.02
R11094 VDD99.n292 VDD99 2301.38
R11095 VDD99.n265 VDD99 2301.38
R11096 VDD99.n293 VDD99.n292 1842.37
R11097 VDD99.n266 VDD99.n265 1842.37
R11098 VDD99.n296 VDD99.t261 1403.56
R11099 VDD99.n298 VDD99.t56 1242.86
R11100 VDD99.n289 VDD99.t75 1105.93
R11101 VDD99.t345 VDD99.n283 1011.51
R11102 VDD99.t292 VDD99.n269 857.144
R11103 VDD99.t176 VDD99.n273 857.144
R11104 VDD99.n292 VDD99.t143 812.681
R11105 VDD99.n265 VDD99.t409 812.681
R11106 VDD99.t3 VDD99.t58 765.152
R11107 VDD99.t395 VDD99.t198 765.152
R11108 VDD99.t438 VDD99.t416 765.152
R11109 VDD99.t245 VDD99.t356 765.152
R11110 VDD99.t316 VDD99.t321 765.152
R11111 VDD99.t104 VDD99.t16 765.152
R11112 VDD99.t248 VDD99.t251 765.152
R11113 VDD99.t319 VDD99.t314 765.152
R11114 VDD99.t349 VDD99.t24 765.152
R11115 VDD99.t201 VDD99.t222 765.152
R11116 VDD99.t382 VDD99.t378 765.152
R11117 VDD99.t238 VDD99.t171 765.152
R11118 VDD99.t271 VDD99.t211 765.152
R11119 VDD99.t214 VDD99.t507 765.152
R11120 VDD99.t401 VDD99.t326 765.152
R11121 VDD99.t208 VDD99.t63 765.152
R11122 VDD99.t505 VDD99.t217 765.152
R11123 VDD99.t264 VDD99.t6 765.152
R11124 VDD99.t225 VDD99.t228 765.152
R11125 VDD99.t380 VDD99.t385 765.152
R11126 VDD99.t421 VDD99.t290 765.152
R11127 VDD99.t0 VDD99.t328 765.152
R11128 VDD99.t393 VDD99.t196 765.152
R11129 VDD99.t448 VDD99.t391 765.152
R11130 VDD99.t411 VDD99.t435 765.152
R11131 VDD99.t330 VDD99.t190 765.152
R11132 VDD99.t284 VDD99.t282 765.152
R11133 VDD99.t308 VDD99.t81 765.152
R11134 VDD99.t193 VDD99.t332 765.152
R11135 VDD99.t335 VDD99.t280 765.152
R11136 VDD99.t466 VDD99.t403 765.152
R11137 VDD99.t296 VDD99.t145 765.152
R11138 VDD99.t253 VDD99.t35 765.152
R11139 VDD99.t240 VDD99.t117 765.152
R11140 VDD99.t293 VDD99.t147 765.152
R11141 VDD99.t13 VDD99.t33 765.152
R11142 VDD99.t92 VDD99.t235 765.152
R11143 VDD99.t90 VDD99.t95 765.152
R11144 VDD99.t65 VDD99.t29 765.152
R11145 VDD99.t311 VDD99.t452 765.152
R11146 VDD99.t98 VDD99.t87 765.152
R11147 VDD99.t230 VDD99.t31 765.152
R11148 VDD99.t482 VDD99.t273 765.152
R11149 VDD99.t302 VDD99.t110 765.152
R11150 VDD99.t305 VDD99.t276 765.152
R11151 VDD99.t60 VDD99.t474 765.152
R11152 VDD99.t299 VDD99.t112 765.152
R11153 VDD99.t26 VDD99.t278 765.152
R11154 VDD99.n290 VDD99.t71 581.375
R11155 VDD99 VDD99.n290 572.967
R11156 VDD99.n485 VDD99.t11 480.199
R11157 VDD99.t261 VDD99.t158 461.096
R11158 VDD99.t261 VDD99.t138 461.096
R11159 VDD99.t140 VDD99.t423 461.096
R11160 VDD99.t351 VDD99.t431 461.096
R11161 VDD99 VDD99.n431 429.187
R11162 VDD99 VDD99.n399 429.187
R11163 VDD99 VDD99.n416 429.187
R11164 VDD99.n478 VDD99 427.092
R11165 VDD99 VDD99.n18 426.699
R11166 VDD99 VDD99.n122 426.699
R11167 VDD99 VDD99.n7 426.699
R11168 VDD99 VDD99.n245 426.699
R11169 VDD99.n137 VDD99 424.618
R11170 VDD99 VDD99.n260 424.618
R11171 VDD99.n283 VDD99.t343 420.793
R11172 VDD99.n136 VDD99 418.495
R11173 VDD99 VDD99.n255 418.495
R11174 VDD99.n431 VDD99.t462 386.365
R11175 VDD99.n462 VDD99.t20 386.365
R11176 VDD99.n416 VDD99.t387 386.365
R11177 VDD99.n399 VDD99.t399 386.365
R11178 VDD99.n18 VDD99.t471 386.365
R11179 VDD99.n122 VDD99.t84 386.365
R11180 VDD99.n7 VDD99.t485 386.365
R11181 VDD99.n245 VDD99.t457 386.365
R11182 VDD99.n136 VDD99.t77 378.788
R11183 VDD99.t428 VDD99.n466 375
R11184 VDD99.n463 VDD99.n462 368.159
R11185 VDD99.n292 VDD99.t140 351.586
R11186 VDD99.n265 VDD99.t351 351.586
R11187 VDD99.n466 VDD99.n464 343.137
R11188 VDD99.t8 VDD99.n136 322.223
R11189 VDD99.t406 VDD99.n255 322.223
R11190 VDD99.t120 VDD99.n137 320.635
R11191 VDD99.n260 VDD99.t477 320.635
R11192 VDD99.t205 VDD99.n478 306.118
R11193 VDD99.t187 VDD99.t438 303.031
R11194 VDD99.t162 VDD99.t104 303.031
R11195 VDD99.t365 VDD99.t319 303.031
R11196 VDD99.t184 VDD99.t349 303.031
R11197 VDD99.t171 VDD99.t181 303.031
R11198 VDD99.t326 VDD99.t165 303.031
R11199 VDD99.t371 VDD99.t505 303.031
R11200 VDD99.t150 VDD99.t264 303.031
R11201 VDD99.t362 VDD99.t380 303.031
R11202 VDD99.t168 VDD99.t421 303.031
R11203 VDD99.t368 VDD99.t393 303.031
R11204 VDD99.t155 VDD99.t448 303.031
R11205 VDD99.t435 VDD99.t494 303.031
R11206 VDD99.t81 VDD99.t492 303.031
R11207 VDD99.t374 VDD99.t193 303.031
R11208 VDD99.t490 VDD99.t466 303.031
R11209 VDD99.t117 VDD99.t488 303.031
R11210 VDD99.t376 VDD99.t293 303.031
R11211 VDD99.t235 VDD99.t134 303.031
R11212 VDD99.t452 VDD99.t132 303.031
R11213 VDD99.t358 VDD99.t98 303.031
R11214 VDD99.t130 VDD99.t482 303.031
R11215 VDD99.t474 VDD99.t136 303.031
R11216 VDD99.t360 VDD99.t299 303.031
R11217 VDD99.n481 VDD99.n469 298.536
R11218 VDD99.n485 VDD99.n469 288
R11219 VDD99.n271 VDD99.n270 199.562
R11220 VDD99.n275 VDD99.n274 199.562
R11221 VDD99.n422 VDD99.t440 193.183
R11222 VDD99.n423 VDD99.t3 193.183
R11223 VDD99.n429 VDD99.t198 193.183
R11224 VDD99.n430 VDD99.t187 193.183
R11225 VDD99.n454 VDD99.t101 193.183
R11226 VDD99.n456 VDD99.t245 193.183
R11227 VDD99.n458 VDD99.t316 193.183
R11228 VDD99.n461 VDD99.t162 193.183
R11229 VDD99.n467 VDD99.t428 193.183
R11230 VDD99.n433 VDD99.t346 193.183
R11231 VDD99.n435 VDD99.t248 193.183
R11232 VDD99.n438 VDD99.t365 193.183
R11233 VDD99.n441 VDD99.t184 193.183
R11234 VDD99.n403 VDD99.t173 193.183
R11235 VDD99.n409 VDD99.t222 193.183
R11236 VDD99.n410 VDD99.t382 193.183
R11237 VDD99.n415 VDD99.t181 193.183
R11238 VDD99.n386 VDD99.t323 193.183
R11239 VDD99.n392 VDD99.t211 193.183
R11240 VDD99.n393 VDD99.t214 193.183
R11241 VDD99.n398 VDD99.t165 193.183
R11242 VDD99.n365 VDD99.t258 193.183
R11243 VDD99.n367 VDD99.t208 193.183
R11244 VDD99.n370 VDD99.t371 193.183
R11245 VDD99.n373 VDD99.t150 193.183
R11246 VDD99.n337 VDD99.t425 193.183
R11247 VDD99.n339 VDD99.t225 193.183
R11248 VDD99.n342 VDD99.t362 193.183
R11249 VDD99.n345 VDD99.t168 193.183
R11250 VDD99.n309 VDD99.t443 193.183
R11251 VDD99.n311 VDD99.t0 193.183
R11252 VDD99.n314 VDD99.t368 193.183
R11253 VDD99.n317 VDD99.t155 193.183
R11254 VDD99.n480 VDD99.t445 191.288
R11255 VDD99.t494 VDD99.n28 191.288
R11256 VDD99.n29 VDD99.t330 191.288
R11257 VDD99.t282 VDD99.n39 191.288
R11258 VDD99.n40 VDD99.t433 191.288
R11259 VDD99.t492 VDD99.n62 191.288
R11260 VDD99.n63 VDD99.t374 191.288
R11261 VDD99.t280 VDD99.n71 191.288
R11262 VDD99.n72 VDD99.t79 191.288
R11263 VDD99.n121 VDD99.t490 191.288
R11264 VDD99.n120 VDD99.t145 191.288
R11265 VDD99.t35 VDD99.n86 191.288
R11266 VDD99.n88 VDD99.t469 191.288
R11267 VDD99.t488 VDD99.n99 191.288
R11268 VDD99.n100 VDD99.t376 191.288
R11269 VDD99.t33 VDD99.n108 191.288
R11270 VDD99.n109 VDD99.t115 191.288
R11271 VDD99.n129 VDD99.t77 191.288
R11272 VDD99.t134 VDD99.n152 191.288
R11273 VDD99.n153 VDD99.t90 191.288
R11274 VDD99.t29 VDD99.n163 191.288
R11275 VDD99.n164 VDD99.t233 191.288
R11276 VDD99.t132 VDD99.n185 191.288
R11277 VDD99.n186 VDD99.t358 191.288
R11278 VDD99.t31 VDD99.n194 191.288
R11279 VDD99.n195 VDD99.t455 191.288
R11280 VDD99.n244 VDD99.t130 191.288
R11281 VDD99.n243 VDD99.t110 191.288
R11282 VDD99.t276 VDD99.n209 191.288
R11283 VDD99.n211 VDD99.t480 191.288
R11284 VDD99.t136 VDD99.n222 191.288
R11285 VDD99.n223 VDD99.t360 191.288
R11286 VDD99.t278 VDD99.n231 191.288
R11287 VDD99.n232 VDD99.t478 191.288
R11288 VDD99.n252 VDD99.t460 191.288
R11289 VDD99.t37 VDD99.t345 175.631
R11290 VDD99.n270 VDD99.t292 170.577
R11291 VDD99.n270 VDD99.t256 170.577
R11292 VDD99.n274 VDD99.t176 170.577
R11293 VDD99.n274 VDD99.t106 170.577
R11294 VDD99.t341 VDD99.n285 153.678
R11295 VDD99.t445 VDD99.t268 151.516
R11296 VDD99.n138 VDD99.t120 142.857
R11297 VDD99.t477 VDD99.n258 142.857
R11298 VDD99.n466 VDD99.t38 132.353
R11299 VDD99.n477 VDD99.t18 124.511
R11300 VDD99.n481 VDD99.n480 117.216
R11301 VDD99.n464 VDD99.n463 112.746
R11302 VDD99.n28 VDD99.t471 111.743
R11303 VDD99.n29 VDD99.t411 111.743
R11304 VDD99.n39 VDD99.t190 111.743
R11305 VDD99.n40 VDD99.t284 111.743
R11306 VDD99.n62 VDD99.t45 111.743
R11307 VDD99.n63 VDD99.t308 111.743
R11308 VDD99.n71 VDD99.t332 111.743
R11309 VDD99.n72 VDD99.t335 111.743
R11310 VDD99.t84 VDD99.n121 111.743
R11311 VDD99.t403 VDD99.n120 111.743
R11312 VDD99.n86 VDD99.t296 111.743
R11313 VDD99.n88 VDD99.t253 111.743
R11314 VDD99.n99 VDD99.t49 111.743
R11315 VDD99.n100 VDD99.t240 111.743
R11316 VDD99.n108 VDD99.t147 111.743
R11317 VDD99.n109 VDD99.t13 111.743
R11318 VDD99.n129 VDD99.t496 111.743
R11319 VDD99.n152 VDD99.t485 111.743
R11320 VDD99.n153 VDD99.t92 111.743
R11321 VDD99.n163 VDD99.t95 111.743
R11322 VDD99.n164 VDD99.t65 111.743
R11323 VDD99.n185 VDD99.t41 111.743
R11324 VDD99.n186 VDD99.t311 111.743
R11325 VDD99.n194 VDD99.t87 111.743
R11326 VDD99.n195 VDD99.t230 111.743
R11327 VDD99.t457 VDD99.n244 111.743
R11328 VDD99.t273 VDD99.n243 111.743
R11329 VDD99.n209 VDD99.t302 111.743
R11330 VDD99.n211 VDD99.t305 111.743
R11331 VDD99.n222 VDD99.t53 111.743
R11332 VDD99.n223 VDD99.t60 111.743
R11333 VDD99.n231 VDD99.t112 111.743
R11334 VDD99.n232 VDD99.t26 111.743
R11335 VDD99.n252 VDD99.t124 111.743
R11336 VDD99.n138 VDD99.t8 111.112
R11337 VDD99.n258 VDD99.t406 111.112
R11338 VDD99.t58 VDD99.n422 109.849
R11339 VDD99.n423 VDD99.t395 109.849
R11340 VDD99.t416 VDD99.n429 109.849
R11341 VDD99.t462 VDD99.n430 109.849
R11342 VDD99.t356 VDD99.n454 109.849
R11343 VDD99.t321 VDD99.n456 109.849
R11344 VDD99.t16 VDD99.n458 109.849
R11345 VDD99.t20 VDD99.n461 109.849
R11346 VDD99.n467 VDD99.t266 109.849
R11347 VDD99.t251 VDD99.n433 109.849
R11348 VDD99.t314 VDD99.n435 109.849
R11349 VDD99.t24 VDD99.n438 109.849
R11350 VDD99.n441 VDD99.t22 109.849
R11351 VDD99.n403 VDD99.t201 109.849
R11352 VDD99.t378 VDD99.n409 109.849
R11353 VDD99.n410 VDD99.t238 109.849
R11354 VDD99.t387 VDD99.n415 109.849
R11355 VDD99.n386 VDD99.t271 109.849
R11356 VDD99.t507 VDD99.n392 109.849
R11357 VDD99.n393 VDD99.t401 109.849
R11358 VDD99.t399 VDD99.n398 109.849
R11359 VDD99.t63 VDD99.n365 109.849
R11360 VDD99.t217 VDD99.n367 109.849
R11361 VDD99.t6 VDD99.n370 109.849
R11362 VDD99.n373 VDD99.t397 109.849
R11363 VDD99.t228 VDD99.n337 109.849
R11364 VDD99.t385 VDD99.n339 109.849
R11365 VDD99.t290 VDD99.n342 109.849
R11366 VDD99.n345 VDD99.t389 109.849
R11367 VDD99.t328 VDD99.n309 109.849
R11368 VDD99.t196 VDD99.n311 109.849
R11369 VDD99.t391 VDD99.n314 109.849
R11370 VDD99.n317 VDD99.t464 109.849
R11371 VDD99.t268 VDD99.n476 96.5914
R11372 VDD99.n479 VDD99.n477 90.2261
R11373 VDD99.n290 VDD99.t414 80.0005
R11374 VDD99.n479 VDD99.t205 76.2337
R11375 VDD99.t56 VDD99 68.2053
R11376 VDD99.n283 VDD99 65.7064
R11377 VDD99.n18 VDD99.t502 62.1896
R11378 VDD99.n122 VDD99.t499 62.1896
R11379 VDD99.n7 VDD99.t127 62.1896
R11380 VDD99.n245 VDD99.t121 62.1896
R11381 VDD99.n298 VDD99.t450 61.9053
R11382 VDD99.n137 VDD99.t219 61.8817
R11383 VDD99.n260 VDD99.t338 61.8817
R11384 VDD99 VDD99.n463 61.0269
R11385 VDD99.n136 VDD99.t287 60.9761
R11386 VDD99.n255 VDD99.t68 60.9761
R11387 VDD99.n431 VDD99.t177 59.702
R11388 VDD99.n462 VDD99.t160 59.702
R11389 VDD99.n416 VDD99.t153 59.702
R11390 VDD99.n399 VDD99.t179 59.702
R11391 VDD99.n478 VDD99.t206 59.4064
R11392 VDD99.n286 VDD99.t75 55.0852
R11393 VDD99.t71 VDD99.n289 55.0852
R11394 VDD99.n476 VDD99.t418 54.9247
R11395 VDD99.n49 VDD99.t48 30.9379
R11396 VDD99.n173 VDD99.t52 30.9379
R11397 VDD99.n52 VDD99.t44 30.2877
R11398 VDD99.n176 VDD99.t40 30.2877
R11399 VDD99 VDD99.n518 25.8059
R11400 VDD99.n53 VDD99.t511 24.5101
R11401 VDD99.n49 VDD99.t510 24.5101
R11402 VDD99.n175 VDD99.t513 24.5101
R11403 VDD99.n173 VDD99.t515 24.5101
R11404 VDD99.n285 VDD99.t37 21.9544
R11405 VDD99.n480 VDD99.n479 20.147
R11406 VDD99.n281 VDD99.t72 14.0055
R11407 VDD99.n284 VDD99.t342 13.2223
R11408 VDD99.n287 VDD99.t76 12.3869
R11409 VDD99.n276 VDD99.t57 12.3869
R11410 VDD99.n281 VDD99.t415 10.1341
R11411 VDD99.n483 VDD99.n482 9.64171
R11412 VDD99.n517 VDD99.n516 8.64364
R11413 VDD99.n177 VDD99.n174 8.14131
R11414 VDD99.n51 VDD99.n50 8.14083
R11415 VDD99.n54 VDD99.n53 8.0005
R11416 VDD99.n175 VDD99.n172 8.0005
R11417 VDD99.n484 VDD99.n483 6.69176
R11418 VDD99 VDD99.n485 6.3005
R11419 VDD99.n487 VDD99.n469 6.3005
R11420 VDD99 VDD99.n481 6.3005
R11421 VDD99.n490 VDD99.n467 6.3005
R11422 VDD99 VDD99.n464 6.3005
R11423 VDD99.n442 VDD99.n441 6.3005
R11424 VDD99.n445 VDD99.n438 6.3005
R11425 VDD99.n448 VDD99.n435 6.3005
R11426 VDD99.n451 VDD99.n433 6.3005
R11427 VDD99.n504 VDD99.n454 6.3005
R11428 VDD99.n501 VDD99.n456 6.3005
R11429 VDD99.n498 VDD99.n458 6.3005
R11430 VDD99.n495 VDD99.n461 6.3005
R11431 VDD99.n374 VDD99.n373 6.3005
R11432 VDD99.n377 VDD99.n370 6.3005
R11433 VDD99.n380 VDD99.n367 6.3005
R11434 VDD99.n383 VDD99.n365 6.3005
R11435 VDD99.n387 VDD99.n386 6.3005
R11436 VDD99.n392 VDD99.n391 6.3005
R11437 VDD99.n394 VDD99.n393 6.3005
R11438 VDD99.n398 VDD99.n397 6.3005
R11439 VDD99.n346 VDD99.n345 6.3005
R11440 VDD99.n349 VDD99.n342 6.3005
R11441 VDD99.n352 VDD99.n339 6.3005
R11442 VDD99.n355 VDD99.n337 6.3005
R11443 VDD99.n404 VDD99.n403 6.3005
R11444 VDD99.n409 VDD99.n408 6.3005
R11445 VDD99.n411 VDD99.n410 6.3005
R11446 VDD99.n415 VDD99.n414 6.3005
R11447 VDD99.n318 VDD99.n317 6.3005
R11448 VDD99.n321 VDD99.n314 6.3005
R11449 VDD99.n324 VDD99.n311 6.3005
R11450 VDD99.n327 VDD99.n309 6.3005
R11451 VDD99.n422 VDD99.n421 6.3005
R11452 VDD99.n424 VDD99.n423 6.3005
R11453 VDD99.n429 VDD99.n428 6.3005
R11454 VDD99.n509 VDD99.n430 6.3005
R11455 VDD99.n285 VDD99.n284 6.3005
R11456 VDD99.n289 VDD99.n288 6.3005
R11457 VDD99 VDD99.n286 6.3005
R11458 VDD99.n299 VDD99.n298 6.3005
R11459 VDD99.n269 VDD99 6.3005
R11460 VDD99.n273 VDD99 6.3005
R11461 VDD99.n28 VDD99.n27 6.3005
R11462 VDD99.n30 VDD99.n29 6.3005
R11463 VDD99.n39 VDD99.n38 6.3005
R11464 VDD99.n41 VDD99.n40 6.3005
R11465 VDD99.n62 VDD99.n61 6.3005
R11466 VDD99.n64 VDD99.n63 6.3005
R11467 VDD99.n71 VDD99.n70 6.3005
R11468 VDD99.n73 VDD99.n72 6.3005
R11469 VDD99.n99 VDD99.n98 6.3005
R11470 VDD99.n101 VDD99.n100 6.3005
R11471 VDD99.n108 VDD99.n107 6.3005
R11472 VDD99.n110 VDD99.n109 6.3005
R11473 VDD99.n120 VDD99.n119 6.3005
R11474 VDD99.n116 VDD99.n86 6.3005
R11475 VDD99.n113 VDD99.n88 6.3005
R11476 VDD99.n121 VDD99.n78 6.3005
R11477 VDD99.n130 VDD99.n129 6.3005
R11478 VDD99.n139 VDD99.n138 6.3005
R11479 VDD99.n152 VDD99.n151 6.3005
R11480 VDD99.n154 VDD99.n153 6.3005
R11481 VDD99.n163 VDD99.n162 6.3005
R11482 VDD99.n165 VDD99.n164 6.3005
R11483 VDD99.n185 VDD99.n184 6.3005
R11484 VDD99.n187 VDD99.n186 6.3005
R11485 VDD99.n194 VDD99.n193 6.3005
R11486 VDD99.n196 VDD99.n195 6.3005
R11487 VDD99.n222 VDD99.n221 6.3005
R11488 VDD99.n224 VDD99.n223 6.3005
R11489 VDD99.n231 VDD99.n230 6.3005
R11490 VDD99.n233 VDD99.n232 6.3005
R11491 VDD99.n243 VDD99.n242 6.3005
R11492 VDD99.n239 VDD99.n209 6.3005
R11493 VDD99.n236 VDD99.n211 6.3005
R11494 VDD99.n244 VDD99.n201 6.3005
R11495 VDD99.n253 VDD99.n252 6.3005
R11496 VDD99.n521 VDD99.n258 6.3005
R11497 VDD99.n291 VDD99.t144 5.85907
R11498 VDD99.n135 VDD99.n132 5.85007
R11499 VDD99.n523 VDD99.n256 5.85007
R11500 VDD99.n511 VDD99.n510 5.69603
R11501 VDD99.n442 VDD99.t23 5.213
R11502 VDD99.n374 VDD99.t398 5.213
R11503 VDD99.n346 VDD99.t390 5.213
R11504 VDD99.n318 VDD99.t465 5.213
R11505 VDD99.n98 VDD99.n94 5.213
R11506 VDD99.n221 VDD99.n217 5.213
R11507 VDD99.n19 VDD99.n16 5.17567
R11508 VDD99.n36 VDD99.n35 5.17567
R11509 VDD99 VDD99.n17 5.16369
R11510 VDD99.n489 VDD99.t267 5.15377
R11511 VDD99.n491 VDD99.n465 5.13287
R11512 VDD99.n473 VDD99.n472 5.13287
R11513 VDD99.n474 VDD99.t420 5.13287
R11514 VDD99.n474 VDD99.t419 5.13287
R11515 VDD99.n494 VDD99.t21 5.13287
R11516 VDD99.n497 VDD99.t17 5.13287
R11517 VDD99.n499 VDD99.n457 5.13287
R11518 VDD99.n500 VDD99.t322 5.13287
R11519 VDD99.n502 VDD99.n455 5.13287
R11520 VDD99.n503 VDD99.t357 5.13287
R11521 VDD99.n505 VDD99.n453 5.13287
R11522 VDD99.n444 VDD99.t25 5.13287
R11523 VDD99.n447 VDD99.t315 5.13287
R11524 VDD99.n449 VDD99.n434 5.13287
R11525 VDD99.n450 VDD99.t252 5.13287
R11526 VDD99.n452 VDD99.n432 5.13287
R11527 VDD99.n357 VDD99.t400 5.13287
R11528 VDD99.n395 VDD99.t402 5.13287
R11529 VDD99.n361 VDD99.n360 5.13287
R11530 VDD99.n390 VDD99.t508 5.13287
R11531 VDD99.n389 VDD99.n362 5.13287
R11532 VDD99.n388 VDD99.t272 5.13287
R11533 VDD99.n385 VDD99.n363 5.13287
R11534 VDD99.n376 VDD99.t7 5.13287
R11535 VDD99.n379 VDD99.t218 5.13287
R11536 VDD99.n381 VDD99.n366 5.13287
R11537 VDD99.n382 VDD99.t64 5.13287
R11538 VDD99.n384 VDD99.n364 5.13287
R11539 VDD99.n348 VDD99.t291 5.13287
R11540 VDD99.n351 VDD99.t386 5.13287
R11541 VDD99.n353 VDD99.n338 5.13287
R11542 VDD99.n354 VDD99.t229 5.13287
R11543 VDD99.n356 VDD99.n336 5.13287
R11544 VDD99.n329 VDD99.t388 5.13287
R11545 VDD99.n412 VDD99.t239 5.13287
R11546 VDD99.n333 VDD99.n332 5.13287
R11547 VDD99.n407 VDD99.t379 5.13287
R11548 VDD99.n406 VDD99.n334 5.13287
R11549 VDD99.n405 VDD99.t202 5.13287
R11550 VDD99.n402 VDD99.n335 5.13287
R11551 VDD99.n508 VDD99.t463 5.13287
R11552 VDD99.n427 VDD99.t417 5.13287
R11553 VDD99.n426 VDD99.n304 5.13287
R11554 VDD99.n425 VDD99.t396 5.13287
R11555 VDD99.n306 VDD99.n305 5.13287
R11556 VDD99.n420 VDD99.t59 5.13287
R11557 VDD99.n419 VDD99.n307 5.13287
R11558 VDD99.n320 VDD99.t392 5.13287
R11559 VDD99.n323 VDD99.t197 5.13287
R11560 VDD99.n325 VDD99.n310 5.13287
R11561 VDD99.n326 VDD99.t329 5.13287
R11562 VDD99.n328 VDD99.n308 5.13287
R11563 VDD99.n294 VDD99.t424 5.13287
R11564 VDD99.n280 VDD99.n279 5.13287
R11565 VDD99.n297 VDD99.t139 5.13287
R11566 VDD99.n267 VDD99.t432 5.13287
R11567 VDD99.n263 VDD99.n262 5.13287
R11568 VDD99.n200 VDD99.n199 5.13287
R11569 VDD99.n159 VDD99.n158 5.13287
R11570 VDD99.n166 VDD99.t234 5.13287
R11571 VDD99.n77 VDD99.n76 5.13287
R11572 VDD99.n37 VDD99.t283 5.13287
R11573 VDD99.n32 VDD99.t331 5.13287
R11574 VDD99.n33 VDD99.n14 5.13287
R11575 VDD99.n23 VDD99.n22 5.13287
R11576 VDD99.n42 VDD99.t434 5.13287
R11577 VDD99.n47 VDD99.n46 5.13287
R11578 VDD99.n66 VDD99.n43 5.13287
R11579 VDD99.n69 VDD99.t281 5.13287
R11580 VDD99.n68 VDD99.n67 5.13287
R11581 VDD99.n74 VDD99.t80 5.13287
R11582 VDD99.n84 VDD99.n79 5.13287
R11583 VDD99.n118 VDD99.t146 5.13287
R11584 VDD99.n117 VDD99.n85 5.13287
R11585 VDD99.n115 VDD99.t36 5.13287
R11586 VDD99.n114 VDD99.n87 5.13287
R11587 VDD99.n112 VDD99.t470 5.13287
R11588 VDD99.n93 VDD99.n92 5.13287
R11589 VDD99.n103 VDD99.n89 5.13287
R11590 VDD99.n106 VDD99.t34 5.13287
R11591 VDD99.n105 VDD99.n104 5.13287
R11592 VDD99.n111 VDD99.t116 5.13287
R11593 VDD99.n128 VDD99.n11 5.13287
R11594 VDD99.n131 VDD99.t78 5.13287
R11595 VDD99.n5 VDD99.n4 5.13287
R11596 VDD99.n147 VDD99.n146 5.13287
R11597 VDD99.n155 VDD99.t91 5.13287
R11598 VDD99.n157 VDD99.n2 5.13287
R11599 VDD99.n161 VDD99.t30 5.13287
R11600 VDD99.n171 VDD99.n170 5.13287
R11601 VDD99.n189 VDD99.n167 5.13287
R11602 VDD99.n192 VDD99.t32 5.13287
R11603 VDD99.n191 VDD99.n190 5.13287
R11604 VDD99.n197 VDD99.t456 5.13287
R11605 VDD99.n207 VDD99.n202 5.13287
R11606 VDD99.n241 VDD99.t111 5.13287
R11607 VDD99.n240 VDD99.n208 5.13287
R11608 VDD99.n238 VDD99.t277 5.13287
R11609 VDD99.n237 VDD99.n210 5.13287
R11610 VDD99.n235 VDD99.t481 5.13287
R11611 VDD99.n216 VDD99.n215 5.13287
R11612 VDD99.n226 VDD99.n212 5.13287
R11613 VDD99.n229 VDD99.t279 5.13287
R11614 VDD99.n228 VDD99.n227 5.13287
R11615 VDD99.n234 VDD99.t479 5.13287
R11616 VDD99.n251 VDD99.n0 5.13287
R11617 VDD99.n254 VDD99.t461 5.13287
R11618 VDD99 VDD99.n515 5.13104
R11619 VDD99.n8 VDD99.n6 5.12213
R11620 VDD99 VDD99.t344 5.10424
R11621 VDD99.n482 VDD99.t19 5.09407
R11622 VDD99.n484 VDD99.t12 5.09407
R11623 VDD99.n468 VDD99.t207 5.09407
R11624 VDD99.n492 VDD99.t39 5.09407
R11625 VDD99.n493 VDD99.t161 5.09407
R11626 VDD99.n507 VDD99.t178 5.09407
R11627 VDD99.n400 VDD99.t180 5.09407
R11628 VDD99.n417 VDD99.t154 5.09407
R11629 VDD99.n264 VDD99.t410 5.09407
R11630 VDD99.n268 VDD99.t244 5.09407
R11631 VDD99.n272 VDD99.t109 5.09407
R11632 VDD99.n123 VDD99.n75 5.09407
R11633 VDD99.n10 VDD99.n9 5.09407
R11634 VDD99.n246 VDD99.n198 5.09407
R11635 VDD99.n261 VDD99.n259 5.09407
R11636 VDD99.n300 VDD99.t451 4.9655
R11637 VDD99.n57 VDD99.n56 4.8755
R11638 VDD99.n180 VDD99.n179 4.8755
R11639 VDD99.n271 VDD99.t257 4.40826
R11640 VDD99.n275 VDD99.t107 4.3915
R11641 VDD99.n269 VDD99.t243 4.26489
R11642 VDD99.n273 VDD99.t108 4.26489
R11643 VDD99.n134 VDD99.n133 4.12326
R11644 VDD99.n522 VDD99.n257 4.12326
R11645 VDD99.n486 VDD99.t74 4.11379
R11646 VDD99.n401 VDD99.n356 3.90405
R11647 VDD99.n520 VDD99.n519 3.26184
R11648 VDD99.n476 VDD99.n475 3.1505
R11649 VDD99.n518 VDD99.n517 3.00194
R11650 VDD99.n473 VDD99.n471 2.85787
R11651 VDD99.n496 VDD99.n460 2.85787
R11652 VDD99.n443 VDD99.n440 2.85787
R11653 VDD99.n446 VDD99.n437 2.85787
R11654 VDD99.n396 VDD99.n359 2.85787
R11655 VDD99.n375 VDD99.n372 2.85787
R11656 VDD99.n378 VDD99.n369 2.85787
R11657 VDD99.n347 VDD99.n344 2.85787
R11658 VDD99.n350 VDD99.n341 2.85787
R11659 VDD99.n413 VDD99.n331 2.85787
R11660 VDD99.n303 VDD99.n302 2.85787
R11661 VDD99.n319 VDD99.n316 2.85787
R11662 VDD99.n322 VDD99.n313 2.85787
R11663 VDD99.n295 VDD99.n278 2.85787
R11664 VDD99.n26 VDD99.n21 2.85787
R11665 VDD99.n60 VDD99.n59 2.85787
R11666 VDD99.n65 VDD99.n45 2.85787
R11667 VDD99.n83 VDD99.n81 2.85787
R11668 VDD99.n97 VDD99.n96 2.85787
R11669 VDD99.n102 VDD99.n91 2.85787
R11670 VDD99.n149 VDD99.n144 2.85787
R11671 VDD99.n183 VDD99.n182 2.85787
R11672 VDD99.n188 VDD99.n169 2.85787
R11673 VDD99.n206 VDD99.n204 2.85787
R11674 VDD99.n220 VDD99.n219 2.85787
R11675 VDD99.n225 VDD99.n214 2.85787
R11676 VDD99.n471 VDD99.t446 2.2755
R11677 VDD99.n471 VDD99.n470 2.2755
R11678 VDD99.n460 VDD99.t105 2.2755
R11679 VDD99.n460 VDD99.n459 2.2755
R11680 VDD99.n440 VDD99.t350 2.2755
R11681 VDD99.n440 VDD99.n439 2.2755
R11682 VDD99.n437 VDD99.t320 2.2755
R11683 VDD99.n437 VDD99.n436 2.2755
R11684 VDD99.n359 VDD99.t327 2.2755
R11685 VDD99.n359 VDD99.n358 2.2755
R11686 VDD99.n372 VDD99.t265 2.2755
R11687 VDD99.n372 VDD99.n371 2.2755
R11688 VDD99.n369 VDD99.t506 2.2755
R11689 VDD99.n369 VDD99.n368 2.2755
R11690 VDD99.n344 VDD99.t422 2.2755
R11691 VDD99.n344 VDD99.n343 2.2755
R11692 VDD99.n341 VDD99.t381 2.2755
R11693 VDD99.n341 VDD99.n340 2.2755
R11694 VDD99.n331 VDD99.t172 2.2755
R11695 VDD99.n331 VDD99.n330 2.2755
R11696 VDD99.n302 VDD99.t439 2.2755
R11697 VDD99.n302 VDD99.n301 2.2755
R11698 VDD99.n316 VDD99.t449 2.2755
R11699 VDD99.n316 VDD99.n315 2.2755
R11700 VDD99.n313 VDD99.t394 2.2755
R11701 VDD99.n313 VDD99.n312 2.2755
R11702 VDD99.n278 VDD99.t159 2.2755
R11703 VDD99.n278 VDD99.n277 2.2755
R11704 VDD99.n21 VDD99.t495 2.2755
R11705 VDD99.n21 VDD99.n20 2.2755
R11706 VDD99.n59 VDD99.t493 2.2755
R11707 VDD99.n59 VDD99.n58 2.2755
R11708 VDD99.n45 VDD99.t375 2.2755
R11709 VDD99.n45 VDD99.n44 2.2755
R11710 VDD99.n81 VDD99.t491 2.2755
R11711 VDD99.n81 VDD99.n80 2.2755
R11712 VDD99.n96 VDD99.t489 2.2755
R11713 VDD99.n96 VDD99.n95 2.2755
R11714 VDD99.n91 VDD99.t377 2.2755
R11715 VDD99.n91 VDD99.n90 2.2755
R11716 VDD99.n144 VDD99.t135 2.2755
R11717 VDD99.n144 VDD99.n143 2.2755
R11718 VDD99.n182 VDD99.t133 2.2755
R11719 VDD99.n182 VDD99.n181 2.2755
R11720 VDD99.n169 VDD99.t359 2.2755
R11721 VDD99.n169 VDD99.n168 2.2755
R11722 VDD99.n204 VDD99.t131 2.2755
R11723 VDD99.n204 VDD99.n203 2.2755
R11724 VDD99.n219 VDD99.t137 2.2755
R11725 VDD99.n219 VDD99.n218 2.2755
R11726 VDD99.n214 VDD99.t361 2.2755
R11727 VDD99.n214 VDD99.n213 2.2755
R11728 VDD99.n494 VDD99 2.25904
R11729 VDD99.n50 VDD99.n49 2.11346
R11730 VDD99.n174 VDD99.n173 2.11346
R11731 VDD99.n177 VDD99.n176 1.8236
R11732 VDD99.n52 VDD99.n51 1.82345
R11733 VDD99 VDD99.n200 1.81843
R11734 VDD99 VDD99.n77 1.81843
R11735 VDD99.n19 VDD99 1.79694
R11736 VDD99.n8 VDD99.n5 1.70466
R11737 VDD99.n518 VDD99 1.37046
R11738 VDD99.n112 VDD99.n111 1.16051
R11739 VDD99.n235 VDD99.n234 1.16051
R11740 VDD99.n247 VDD99.n197 1.0737
R11741 VDD99.n506 VDD99.n452 1.02928
R11742 VDD99.n418 VDD99.n328 1.02928
R11743 VDD99.n124 VDD99.n74 1.02347
R11744 VDD99.n385 VDD99.n384 0.881662
R11745 VDD99 VDD99.n297 0.786716
R11746 VDD99.n477 VDD99.t73 0.783764
R11747 VDD99.n24 VDD99.n19 0.682778
R11748 VDD99.n513 VDD99.n268 0.66512
R11749 VDD99.n512 VDD99.n272 0.634017
R11750 VDD99.n180 VDD99.n178 0.608132
R11751 VDD99.n141 VDD99.n8 0.601963
R11752 VDD99.n25 VDD99.n24 0.582756
R11753 VDD99.n36 VDD99.n12 0.582756
R11754 VDD99.n150 VDD99.n142 0.582756
R11755 VDD99.n148 VDD99.n145 0.582756
R11756 VDD99.n34 VDD99.n13 0.5405
R11757 VDD99.n31 VDD99.n15 0.5405
R11758 VDD99.n126 VDD99.n125 0.5405
R11759 VDD99.n156 VDD99.n3 0.5405
R11760 VDD99.n160 VDD99.n1 0.5405
R11761 VDD99.n249 VDD99.n248 0.5405
R11762 VDD99.n82 VDD99 0.468385
R11763 VDD99.n205 VDD99 0.468385
R11764 VDD99.n53 VDD99.n52 0.404541
R11765 VDD99.n176 VDD99.n175 0.404541
R11766 VDD99.n61 VDD99.n57 0.337997
R11767 VDD99.n184 VDD99.n180 0.337997
R11768 VDD99.n57 VDD99.n55 0.328132
R11769 VDD99.n447 VDD99.n446 0.233919
R11770 VDD99.n444 VDD99.n443 0.233919
R11771 VDD99.n379 VDD99.n378 0.233919
R11772 VDD99.n376 VDD99.n375 0.233919
R11773 VDD99.n351 VDD99.n350 0.233919
R11774 VDD99.n348 VDD99.n347 0.233919
R11775 VDD99.n323 VDD99.n322 0.233919
R11776 VDD99.n320 VDD99.n319 0.233919
R11777 VDD99.n60 VDD99.n47 0.233919
R11778 VDD99.n66 VDD99.n65 0.233919
R11779 VDD99.n97 VDD99.n93 0.233919
R11780 VDD99.n103 VDD99.n102 0.233919
R11781 VDD99.n183 VDD99.n171 0.233919
R11782 VDD99.n189 VDD99.n188 0.233919
R11783 VDD99.n220 VDD99.n216 0.233919
R11784 VDD99.n226 VDD99.n225 0.233919
R11785 VDD99 VDD99.n511 0.227487
R11786 VDD99.n488 VDD99.n487 0.224447
R11787 VDD99.n127 VDD99 0.223897
R11788 VDD99.n250 VDD99 0.223897
R11789 VDD99.n493 VDD99 0.205357
R11790 VDD99.n489 VDD99.n488 0.202146
R11791 VDD99.n519 VDD99 0.186599
R11792 VDD99.n250 VDD99.n249 0.178009
R11793 VDD99.n517 VDD99 0.17171
R11794 VDD99.n264 VDD99.n263 0.170231
R11795 VDD99.n507 VDD99.n506 0.167533
R11796 VDD99 VDD99.n329 0.160716
R11797 VDD99.n127 VDD99.n126 0.159769
R11798 VDD99.n508 VDD99 0.158984
R11799 VDD99 VDD99.n357 0.157289
R11800 VDD99.n418 VDD99.n417 0.155496
R11801 VDD99 VDD99.n282 0.154766
R11802 VDD99.n401 VDD99.n400 0.154581
R11803 VDD99.n450 VDD99.n449 0.141016
R11804 VDD99.n382 VDD99.n381 0.141016
R11805 VDD99.n354 VDD99.n353 0.141016
R11806 VDD99.n326 VDD99.n325 0.141016
R11807 VDD99.n33 VDD99.n32 0.141016
R11808 VDD99.n69 VDD99.n68 0.141016
R11809 VDD99.n106 VDD99.n105 0.141016
R11810 VDD99.n118 VDD99.n117 0.141016
R11811 VDD99.n115 VDD99.n114 0.141016
R11812 VDD99.n192 VDD99.n191 0.141016
R11813 VDD99.n229 VDD99.n228 0.141016
R11814 VDD99.n241 VDD99.n240 0.141016
R11815 VDD99.n238 VDD99.n237 0.141016
R11816 VDD99.n124 VDD99.n123 0.139745
R11817 VDD99.n247 VDD99.n246 0.139745
R11818 VDD99 VDD99.n140 0.138536
R11819 VDD99.n140 VDD99.n10 0.137219
R11820 VDD99.n520 VDD99.n261 0.137219
R11821 VDD99.n488 VDD99.n468 0.137126
R11822 VDD99.n402 VDD99.n401 0.131861
R11823 VDD99.n492 VDD99.n491 0.130567
R11824 VDD99.n514 VDD99.n267 0.129503
R11825 VDD99.n514 VDD99 0.12689
R11826 VDD99.n503 VDD99.n502 0.123551
R11827 VDD99.n500 VDD99.n499 0.123551
R11828 VDD99.n406 VDD99.n405 0.123551
R11829 VDD99.n407 VDD99.n333 0.123551
R11830 VDD99.n84 VDD99 0.123016
R11831 VDD99.n207 VDD99 0.123016
R11832 VDD99.n420 VDD99.n306 0.122176
R11833 VDD99.n426 VDD99.n425 0.122176
R11834 VDD99.n389 VDD99.n388 0.120831
R11835 VDD99.n390 VDD99.n361 0.120831
R11836 VDD99.n3 VDD99.n1 0.119765
R11837 VDD99.n506 VDD99.n505 0.116432
R11838 VDD99.n513 VDD99.n512 0.115201
R11839 VDD99.n419 VDD99.n418 0.115137
R11840 VDD99.n249 VDD99.n1 0.112148
R11841 VDD99 VDD99.n83 0.111403
R11842 VDD99.n149 VDD99 0.111403
R11843 VDD99 VDD99.n206 0.111403
R11844 VDD99.n37 VDD99.n36 0.109081
R11845 VDD99.n125 VDD99.n42 0.107919
R11846 VDD99.n50 VDD99 0.107393
R11847 VDD99.n174 VDD99 0.107393
R11848 VDD99.n38 VDD99.n37 0.107339
R11849 VDD99.n491 VDD99.n490 0.107339
R11850 VDD99.n452 VDD99.n451 0.107339
R11851 VDD99.n449 VDD99.n448 0.107339
R11852 VDD99.n384 VDD99.n383 0.107339
R11853 VDD99.n381 VDD99.n380 0.107339
R11854 VDD99.n356 VDD99.n355 0.107339
R11855 VDD99.n353 VDD99.n352 0.107339
R11856 VDD99.n328 VDD99.n327 0.107339
R11857 VDD99.n325 VDD99.n324 0.107339
R11858 VDD99.n266 VDD99.n263 0.107339
R11859 VDD99.n42 VDD99.n41 0.107339
R11860 VDD99.n70 VDD99.n69 0.107339
R11861 VDD99.n74 VDD99.n73 0.107339
R11862 VDD99.n107 VDD99.n106 0.107339
R11863 VDD99.n111 VDD99.n110 0.107339
R11864 VDD99.n119 VDD99.n118 0.107339
R11865 VDD99.n116 VDD99.n115 0.107339
R11866 VDD99.n113 VDD99.n112 0.107339
R11867 VDD99.n155 VDD99.n154 0.107339
R11868 VDD99.n162 VDD99.n161 0.107339
R11869 VDD99.n166 VDD99.n165 0.107339
R11870 VDD99.n193 VDD99.n192 0.107339
R11871 VDD99.n197 VDD99.n196 0.107339
R11872 VDD99.n230 VDD99.n229 0.107339
R11873 VDD99.n234 VDD99.n233 0.107339
R11874 VDD99.n242 VDD99.n241 0.107339
R11875 VDD99.n239 VDD99.n238 0.107339
R11876 VDD99.n236 VDD99.n235 0.107339
R11877 VDD99.n13 VDD99.n12 0.107337
R11878 VDD99.n497 VDD99 0.10728
R11879 VDD99 VDD99.n412 0.10728
R11880 VDD99 VDD99.n26 0.106758
R11881 VDD99 VDD99.n60 0.106758
R11882 VDD99.n65 VDD99 0.106758
R11883 VDD99 VDD99.n97 0.106758
R11884 VDD99.n102 VDD99 0.106758
R11885 VDD99 VDD99.n183 0.106758
R11886 VDD99.n188 VDD99 0.106758
R11887 VDD99 VDD99.n220 0.106758
R11888 VDD99.n225 VDD99 0.106758
R11889 VDD99.n446 VDD99 0.106177
R11890 VDD99.n443 VDD99 0.106177
R11891 VDD99.n378 VDD99 0.106177
R11892 VDD99.n375 VDD99 0.106177
R11893 VDD99.n350 VDD99 0.106177
R11894 VDD99.n347 VDD99 0.106177
R11895 VDD99.n322 VDD99 0.106177
R11896 VDD99.n319 VDD99 0.106177
R11897 VDD99.n427 VDD99 0.106087
R11898 VDD99 VDD99.n395 0.10492
R11899 VDD99.n145 VDD99.n3 0.10413
R11900 VDD99.n157 VDD99.n156 0.100371
R11901 VDD99.n172 VDD99 0.100075
R11902 VDD99.n141 VDD99 0.09952
R11903 VDD99 VDD99.n496 0.0981271
R11904 VDD99.n413 VDD99 0.0981271
R11905 VDD99 VDD99.n303 0.0970363
R11906 VDD99.n126 VDD99.n12 0.0967138
R11907 VDD99.n513 VDD99.n271 0.096125
R11908 VDD99.n396 VDD99 0.0959696
R11909 VDD99.n145 VDD99.n142 0.0947094
R11910 VDD99.n505 VDD99.n504 0.0940593
R11911 VDD99.n502 VDD99.n501 0.0940593
R11912 VDD99.n499 VDD99.n498 0.0940593
R11913 VDD99.n404 VDD99.n402 0.0940593
R11914 VDD99.n408 VDD99.n406 0.0940593
R11915 VDD99.n411 VDD99.n333 0.0940593
R11916 VDD99.n496 VDD99 0.0930424
R11917 VDD99 VDD99.n413 0.0930424
R11918 VDD99.n421 VDD99.n419 0.093014
R11919 VDD99.n424 VDD99.n306 0.093014
R11920 VDD99.n428 VDD99.n426 0.093014
R11921 VDD99.n387 VDD99.n385 0.0919917
R11922 VDD99.n391 VDD99.n389 0.0919917
R11923 VDD99.n394 VDD99.n361 0.0919917
R11924 VDD99 VDD99.n396 0.0909972
R11925 VDD99.n512 VDD99.n275 0.0905
R11926 VDD99.n248 VDD99.n247 0.089386
R11927 VDD99.n160 VDD99.n159 0.082371
R11928 VDD99.n26 VDD99.n25 0.0817903
R11929 VDD99.n142 VDD99.n141 0.08148
R11930 VDD99.n24 VDD99.n15 0.0808786
R11931 VDD99.n15 VDD99.n13 0.0808786
R11932 VDD99.n445 VDD99.n444 0.080629
R11933 VDD99.n377 VDD99.n376 0.080629
R11934 VDD99.n349 VDD99.n348 0.080629
R11935 VDD99.n321 VDD99.n320 0.080629
R11936 VDD99.n64 VDD99.n47 0.080629
R11937 VDD99.n101 VDD99.n93 0.080629
R11938 VDD99.n187 VDD99.n171 0.080629
R11939 VDD99.n224 VDD99.n216 0.080629
R11940 VDD99 VDD99.n450 0.0794677
R11941 VDD99 VDD99.n447 0.0794677
R11942 VDD99 VDD99.n382 0.0794677
R11943 VDD99 VDD99.n379 0.0794677
R11944 VDD99 VDD99.n354 0.0794677
R11945 VDD99 VDD99.n351 0.0794677
R11946 VDD99 VDD99.n326 0.0794677
R11947 VDD99 VDD99.n323 0.0794677
R11948 VDD99.n23 VDD99 0.0788871
R11949 VDD99 VDD99.n66 0.0788871
R11950 VDD99.n68 VDD99 0.0788871
R11951 VDD99 VDD99.n103 0.0788871
R11952 VDD99.n105 VDD99 0.0788871
R11953 VDD99 VDD99.n84 0.0788871
R11954 VDD99.n117 VDD99 0.0788871
R11955 VDD99.n114 VDD99 0.0788871
R11956 VDD99.n147 VDD99 0.0788871
R11957 VDD99 VDD99.n157 0.0788871
R11958 VDD99.n159 VDD99 0.0788871
R11959 VDD99 VDD99.n189 0.0788871
R11960 VDD99.n191 VDD99 0.0788871
R11961 VDD99 VDD99.n226 0.0788871
R11962 VDD99.n228 VDD99 0.0788871
R11963 VDD99 VDD99.n207 0.0788871
R11964 VDD99.n240 VDD99 0.0788871
R11965 VDD99.n237 VDD99 0.0788871
R11966 VDD99 VDD99.n282 0.0786971
R11967 VDD99.n267 VDD99 0.0759839
R11968 VDD99.n519 VDD99.n514 0.0753624
R11969 VDD99.n482 VDD99 0.0709717
R11970 VDD99 VDD99.n468 0.0709717
R11971 VDD99 VDD99.n493 0.0709717
R11972 VDD99 VDD99.n264 0.0709717
R11973 VDD99 VDD99.n268 0.0709717
R11974 VDD99 VDD99.n272 0.0709717
R11975 VDD99.n495 VDD99.n494 0.0706695
R11976 VDD99.n414 VDD99.n329 0.0706695
R11977 VDD99.n123 VDD99 0.0701226
R11978 VDD99 VDD99.n10 0.0701226
R11979 VDD99.n246 VDD99 0.0701226
R11980 VDD99.n261 VDD99 0.0701226
R11981 VDD99.n291 VDD99 0.0700788
R11982 VDD99.n509 VDD99.n508 0.0698855
R11983 VDD99 VDD99.n503 0.0696525
R11984 VDD99 VDD99.n500 0.0696525
R11985 VDD99 VDD99.n497 0.0696525
R11986 VDD99.n405 VDD99 0.0696525
R11987 VDD99 VDD99.n407 0.0696525
R11988 VDD99.n412 VDD99 0.0696525
R11989 VDD99.n397 VDD99.n357 0.0691188
R11990 VDD99.n48 VDD99 0.0690714
R11991 VDD99 VDD99.n420 0.0688799
R11992 VDD99.n425 VDD99 0.0688799
R11993 VDD99 VDD99.n427 0.0688799
R11994 VDD99.n388 VDD99 0.0681243
R11995 VDD99 VDD99.n390 0.0681243
R11996 VDD99.n395 VDD99 0.0681243
R11997 VDD99.n150 VDD99.n149 0.0649516
R11998 VDD99.n140 VDD99.n139 0.0617883
R11999 VDD99.n521 VDD99.n520 0.0617883
R12000 VDD99.n135 VDD99.n134 0.0608681
R12001 VDD99.n523 VDD99.n522 0.0608681
R12002 VDD99.n295 VDD99.n294 0.0598378
R12003 VDD99 VDD99.n131 0.0592117
R12004 VDD99 VDD99.n254 0.0592117
R12005 VDD99.n32 VDD99.n31 0.0591452
R12006 VDD99.n161 VDD99.n160 0.0591452
R12007 VDD99.n25 VDD99.n23 0.0574032
R12008 VDD99.n82 VDD99.n77 0.0556613
R12009 VDD99.n205 VDD99.n200 0.0556613
R12010 VDD99 VDD99.n486 0.0555633
R12011 VDD99 VDD99.n489 0.0550806
R12012 VDD99.n248 VDD99.n166 0.0550806
R12013 VDD99 VDD99.n473 0.0533387
R12014 VDD99.n510 VDD99.n303 0.0532933
R12015 VDD99.n31 VDD99.n30 0.0486936
R12016 VDD99.n55 VDD99.n48 0.0471071
R12017 VDD99 VDD99.n34 0.0452097
R12018 VDD99 VDD99.n492 0.043431
R12019 VDD99.n83 VDD99.n82 0.0417258
R12020 VDD99.n206 VDD99.n205 0.0417258
R12021 VDD99.n156 VDD99.n155 0.0411452
R12022 VDD99 VDD99.n281 0.041
R12023 VDD99.n417 VDD99 0.0404465
R12024 VDD99 VDD99.n507 0.0400238
R12025 VDD99.n400 VDD99 0.0396099
R12026 VDD99.n510 VDD99 0.0392151
R12027 VDD99.n54 VDD99.n51 0.0387493
R12028 VDD99 VDD99.n474 0.0382419
R12029 VDD99.n55 VDD99.n54 0.0358571
R12030 VDD99.n178 VDD99.n177 0.0344878
R12031 VDD99.n483 VDD99.n473 0.0344677
R12032 VDD99.n131 VDD99.n130 0.034365
R12033 VDD99.n254 VDD99.n253 0.034365
R12034 VDD99.n34 VDD99.n33 0.0341774
R12035 VDD99 VDD99.n280 0.0333767
R12036 VDD99.n288 VDD99.n287 0.0327683
R12037 VDD99 VDD99.n484 0.032019
R12038 VDD99.n125 VDD99.n124 0.0292131
R12039 VDD99.n287 VDD99 0.028378
R12040 VDD99.n150 VDD99.n5 0.0277903
R12041 VDD99.n134 VDD99 0.0270031
R12042 VDD99.n522 VDD99 0.0270031
R12043 VDD99.n148 VDD99.n147 0.0254677
R12044 VDD99.n299 VDD99.n276 0.0254153
R12045 VDD99 VDD99.n128 0.0242423
R12046 VDD99 VDD99.n251 0.0242423
R12047 VDD99.n128 VDD99.n127 0.0235061
R12048 VDD99.n251 VDD99.n250 0.0235061
R12049 VDD99 VDD99.n276 0.0220254
R12050 VDD99.n82 VDD99.n78 0.0206923
R12051 VDD99.n205 VDD99.n201 0.0206923
R12052 VDD99.n151 VDD99.n150 0.0197073
R12053 VDD99.n293 VDD99.n280 0.0194041
R12054 VDD99 VDD99.n295 0.0192629
R12055 VDD99.n36 VDD99 0.0155968
R12056 VDD99.n300 VDD99 0.0147732
R12057 VDD99.n297 VDD99.n296 0.0147268
R12058 VDD99.n294 VDD99 0.0138562
R12059 VDD99 VDD99.n282 0.0127264
R12060 VDD99.n512 VDD99 0.0120325
R12061 VDD99.n178 VDD99.n172 0.0119894
R12062 VDD99.n511 VDD99.n300 0.0112532
R12063 VDD99.n48 VDD99 0.00907143
R12064 VDD99.n8 VDD99 0.00708537
R12065 VDD99.n27 VDD99.n19 0.0068871
R12066 VDD99.n25 VDD99 0.00653659
R12067 VDD99.n486 VDD99 0.00543671
R12068 VDD99.n490 VDD99 0.00514516
R12069 VDD99 VDD99.n266 0.00514516
R12070 VDD99 VDD99.n513 0.00501948
R12071 VDD99 VDD99.n281 0.00368293
R12072 VDD99.n487 VDD99 0.00315823
R12073 VDD99.n475 VDD99 0.00282258
R12074 VDD99 VDD99.n148 0.00282258
R12075 VDD99.n38 VDD99 0.00224194
R12076 VDD99.n30 VDD99 0.00224194
R12077 VDD99.n41 VDD99 0.00224194
R12078 VDD99.n70 VDD99 0.00224194
R12079 VDD99.n73 VDD99 0.00224194
R12080 VDD99.n107 VDD99 0.00224194
R12081 VDD99.n110 VDD99 0.00224194
R12082 VDD99.n119 VDD99 0.00224194
R12083 VDD99 VDD99.n116 0.00224194
R12084 VDD99 VDD99.n113 0.00224194
R12085 VDD99.n154 VDD99 0.00224194
R12086 VDD99.n162 VDD99 0.00224194
R12087 VDD99.n165 VDD99 0.00224194
R12088 VDD99.n193 VDD99 0.00224194
R12089 VDD99.n196 VDD99 0.00224194
R12090 VDD99.n230 VDD99 0.00224194
R12091 VDD99.n233 VDD99 0.00224194
R12092 VDD99.n242 VDD99 0.00224194
R12093 VDD99 VDD99.n239 0.00224194
R12094 VDD99 VDD99.n236 0.00224194
R12095 VDD99.n130 VDD99 0.00215644
R12096 VDD99.n253 VDD99 0.00215644
R12097 VDD99.n139 VDD99 0.00178834
R12098 VDD99 VDD99.n521 0.00178834
R12099 VDD99.n451 VDD99 0.00166129
R12100 VDD99.n448 VDD99 0.00166129
R12101 VDD99 VDD99.n445 0.00166129
R12102 VDD99 VDD99.n442 0.00166129
R12103 VDD99.n383 VDD99 0.00166129
R12104 VDD99.n380 VDD99 0.00166129
R12105 VDD99 VDD99.n377 0.00166129
R12106 VDD99 VDD99.n374 0.00166129
R12107 VDD99.n355 VDD99 0.00166129
R12108 VDD99.n352 VDD99 0.00166129
R12109 VDD99 VDD99.n349 0.00166129
R12110 VDD99 VDD99.n346 0.00166129
R12111 VDD99.n327 VDD99 0.00166129
R12112 VDD99.n324 VDD99 0.00166129
R12113 VDD99 VDD99.n321 0.00166129
R12114 VDD99 VDD99.n318 0.00166129
R12115 VDD99.n504 VDD99 0.00151695
R12116 VDD99.n501 VDD99 0.00151695
R12117 VDD99.n498 VDD99 0.00151695
R12118 VDD99 VDD99.n495 0.00151695
R12119 VDD99 VDD99.n404 0.00151695
R12120 VDD99.n408 VDD99 0.00151695
R12121 VDD99 VDD99.n411 0.00151695
R12122 VDD99.n414 VDD99 0.00151695
R12123 VDD99.n421 VDD99 0.00150559
R12124 VDD99 VDD99.n424 0.00150559
R12125 VDD99.n428 VDD99 0.00150559
R12126 VDD99 VDD99.n509 0.00150559
R12127 VDD99 VDD99.n387 0.00149448
R12128 VDD99.n391 VDD99 0.00149448
R12129 VDD99 VDD99.n394 0.00149448
R12130 VDD99.n397 VDD99 0.00149448
R12131 VDD99 VDD99.n293 0.00132192
R12132 VDD99.n475 VDD99 0.00108064
R12133 VDD99.n27 VDD99 0.00108064
R12134 VDD99.n61 VDD99 0.00108064
R12135 VDD99 VDD99.n64 0.00108064
R12136 VDD99.n98 VDD99 0.00108064
R12137 VDD99 VDD99.n101 0.00108064
R12138 VDD99.n184 VDD99 0.00108064
R12139 VDD99 VDD99.n187 0.00108064
R12140 VDD99.n221 VDD99 0.00108064
R12141 VDD99 VDD99.n224 0.00108064
R12142 VDD99.n78 VDD99 0.00107692
R12143 VDD99.n201 VDD99 0.00107692
R12144 VDD99.n151 VDD99 0.00104878
R12145 VDD99.n284 VDD99 0.00100943
R12146 VDD99 VDD99.n135 0.000868098
R12147 VDD99 VDD99.n523 0.000868098
R12148 VDD99.n288 VDD99 0.000719512
R12149 VDD99.n296 VDD99 0.000706186
R12150 VDD99 VDD99.n291 0.000705479
R12151 VDD99 VDD99.n299 0.000669492
R12152 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n4 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t9 36.935
R12153 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n13 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t6 36.935
R12154 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n12 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t10 36.935
R12155 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n5 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t15 31.528
R12156 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n6 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t13 31.528
R12157 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n9 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t4 31.4332
R12158 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n11 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t5 25.5364
R12159 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n4 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t11 18.1962
R12160 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n13 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t7 18.1962
R12161 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n12 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t14 18.1962
R12162 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n9 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t8 15.3826
R12163 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n5 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t3 15.3826
R12164 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n6 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t16 15.3826
R12165 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n11 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t12 14.0749
R12166 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n5 7.63417
R12167 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n6 7.62076
R12168 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t1 7.09905
R12169 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n9 6.86029
R12170 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n8 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n7 6.65668
R12171 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n7 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 5.46205
R12172 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n7 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 4.73586
R12173 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n10 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n8 3.41968
R12174 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n3 3.25053
R12175 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n3 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t2 2.2755
R12176 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n3 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n2 2.2755
R12177 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n4 2.13459
R12178 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n13 2.13151
R12179 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 2.63808
R12180 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n12 2.13042
R12181 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n8 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 1.5916
R12182 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n10 1.49033
R12183 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n11 1.43689
R12184 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n0 1.22411
R12185 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n10 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 1.12067
R12186 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n0 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 1.12013
R12187 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n1 1.11863
R12188 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n0 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n1 0.927577
R12189 VDD100.n433 VDD100.n94 190685
R12190 VDD100.n433 VDD100.t470 83097.6
R12191 VDD100.n330 VDD100.t359 29077.7
R12192 VDD100.n398 VDD100.n397 11185.2
R12193 VDD100.n357 VDD100.n356 11185.2
R12194 VDD100.t390 VDD100.n88 1105.93
R12195 VDD100.n334 VDD100.t121 1105.93
R12196 VDD100.t301 VDD100.t111 961.905
R12197 VDD100.t410 VDD100.t330 961.905
R12198 VDD100.t466 VDD100.t270 961.905
R12199 VDD100.t125 VDD100.t163 961.905
R12200 VDD100.t264 VDD100.t328 961.905
R12201 VDD100.t198 VDD100.t46 961.905
R12202 VDD100.t3 VDD100.t322 765.152
R12203 VDD100.t0 VDD100.t113 765.152
R12204 VDD100.t17 VDD100.t129 765.152
R12205 VDD100.t6 VDD100.t325 765.152
R12206 VDD100.t338 VDD100.t115 765.152
R12207 VDD100.t401 VDD100.t28 765.152
R12208 VDD100.t57 VDD100.t51 765.152
R12209 VDD100.t157 VDD100.t249 765.152
R12210 VDD100.t25 VDD100.t144 765.152
R12211 VDD100.t53 VDD100.t55 765.152
R12212 VDD100.t311 VDD100.t196 765.152
R12213 VDD100.t267 VDD100.t44 765.152
R12214 VDD100.t119 VDD100.t20 765.152
R12215 VDD100.t216 VDD100.t293 765.152
R12216 VDD100.t200 VDD100.t11 765.152
R12217 VDD100.t141 VDD100.t262 765.152
R12218 VDD100.t332 VDD100.t363 765.152
R12219 VDD100.t347 VDD100.t319 765.152
R12220 VDD100.t186 VDD100.t399 765.152
R12221 VDD100.t354 VDD100.t350 765.152
R12222 VDD100.t135 VDD100.t437 765.152
R12223 VDD100.t34 VDD100.t289 765.152
R12224 VDD100.t387 VDD100.t194 765.152
R12225 VDD100.t295 VDD100.t415 765.152
R12226 VDD100.t189 VDD100.t396 765.152
R12227 VDD100.t277 VDD100.t352 765.152
R12228 VDD100.t234 VDD100.t254 765.152
R12229 VDD100.t138 VDD100.t259 765.152
R12230 VDD100.t393 VDD100.t365 765.152
R12231 VDD100.t463 VDD100.t146 765.152
R12232 VDD100.t151 VDD100.t39 765.152
R12233 VDD100.t179 VDD100.t106 765.152
R12234 VDD100.t298 VDD100.t62 765.152
R12235 VDD100.t309 VDD100.t272 765.152
R12236 VDD100.t443 VDD100.t335 765.152
R12237 VDD100.t148 VDD100.t229 765.152
R12238 VDD100.t286 VDD100.t31 765.152
R12239 VDD100.t432 VDD100.t192 765.152
R12240 VDD100.n397 VDD100.t153 676.191
R12241 VDD100.n356 VDD100.t117 676.191
R12242 VDD100.t274 VDD100.n94 669.048
R12243 VDD100.t159 VDD100.t161 645.307
R12244 VDD100.t280 VDD100.t304 642.843
R12245 VDD100.n433 VDD100.n90 525.424
R12246 VDD100.n331 VDD100.n330 525.424
R12247 VDD100.n398 VDD100.t247 485.714
R12248 VDD100.n357 VDD100.t69 485.714
R12249 VDD100 VDD100.n185 429.187
R12250 VDD100 VDD100.n340 427.092
R12251 VDD100.n346 VDD100 427.092
R12252 VDD100 VDD100.n246 426.699
R12253 VDD100 VDD100.n258 426.699
R12254 VDD100 VDD100.n478 426.699
R12255 VDD100.t461 VDD100.n398 426.44
R12256 VDD100.t171 VDD100.n357 426.44
R12257 VDD100 VDD100.n335 425.019
R12258 VDD100 VDD100.n79 424.618
R12259 VDD100 VDD100.n83 424.618
R12260 VDD100 VDD100.n87 422.557
R12261 VDD100.n478 VDD100.t14 386.365
R12262 VDD100.t224 VDD100.n79 386.365
R12263 VDD100.t239 VDD100.n83 386.365
R12264 VDD100.n185 VDD100.t155 386.365
R12265 VDD100.n346 VDD100.t214 386.365
R12266 VDD100.n340 VDD100.t456 386.365
R12267 VDD100.t132 VDD100.n246 386.365
R12268 VDD100.n258 VDD100.t65 386.365
R12269 VDD100.t470 VDD100.t410 380.952
R12270 VDD100.t163 VDD100.t453 380.952
R12271 VDD100.t46 VDD100.t168 380.952
R12272 VDD100.n79 VDD100.t222 378.788
R12273 VDD100.n83 VDD100.t430 378.788
R12274 VDD100.n87 VDD100.t232 378.788
R12275 VDD100.t211 VDD100.n346 378.788
R12276 VDD100.n340 VDD100.t173 378.788
R12277 VDD100.n335 VDD100.t208 378.788
R12278 VDD100.t403 VDD100.t341 303.031
R12279 VDD100.t322 VDD100.t375 303.031
R12280 VDD100.t129 VDD100.t245 303.031
R12281 VDD100.t249 VDD100.t448 303.031
R12282 VDD100.t369 VDD100.t53 303.031
R12283 VDD100.t440 VDD100.t311 303.031
R12284 VDD100.t379 VDD100.t119 303.031
R12285 VDD100.t181 VDD100.t216 303.031
R12286 VDD100.t359 VDD100.t200 303.031
R12287 VDD100.t319 VDD100.t257 303.031
R12288 VDD100.t437 VDD100.t420 303.031
R12289 VDD100.t415 VDD100.t237 303.031
R12290 VDD100.t385 VDD100.t189 303.031
R12291 VDD100.t254 VDD100.t357 303.031
R12292 VDD100.t367 VDD100.t138 303.031
R12293 VDD100.t382 VDD100.t151 303.031
R12294 VDD100.t445 VDD100.t179 303.031
R12295 VDD100.t372 VDD100.t309 303.031
R12296 VDD100.t473 VDD100.t443 303.031
R12297 VDD100.t229 VDD100.t422 303.031
R12298 VDD100.t377 VDD100.t286 303.031
R12299 VDD100.t307 VDD100.n94 292.858
R12300 VDD100.n397 VDD100.t36 285.714
R12301 VDD100.n356 VDD100.t22 285.714
R12302 VDD100.n425 VDD100.t412 242.857
R12303 VDD100.n426 VDD100.t301 242.857
R12304 VDD100.n432 VDD100.t274 242.857
R12305 VDD100.n384 VDD100.t165 242.857
R12306 VDD100.n385 VDD100.t466 242.857
R12307 VDD100.t36 VDD100.n396 242.857
R12308 VDD100.t453 VDD100.n395 242.857
R12309 VDD100.n212 VDD100.t48 242.857
R12310 VDD100.n213 VDD100.t264 242.857
R12311 VDD100.t22 VDD100.n355 242.857
R12312 VDD100.t168 VDD100.n354 242.857
R12313 VDD100.n172 VDD100.t251 193.183
R12314 VDD100.n178 VDD100.t28 193.183
R12315 VDD100.n179 VDD100.t57 193.183
R12316 VDD100.n184 VDD100.t448 193.183
R12317 VDD100.n117 VDD100.t314 193.183
R12318 VDD100.n119 VDD100.t25 193.183
R12319 VDD100.n122 VDD100.t369 193.183
R12320 VDD100.n125 VDD100.t440 193.183
R12321 VDD100.n188 VDD100.t205 193.183
R12322 VDD100.n190 VDD100.t267 193.183
R12323 VDD100.n193 VDD100.t379 193.183
R12324 VDD100.n196 VDD100.t181 193.183
R12325 VDD100.n347 VDD100.t211 193.183
R12326 VDD100.n345 VDD100.t173 193.183
R12327 VDD100.n339 VDD100.t208 193.183
R12328 VDD100.n360 VDD100.t176 193.183
R12329 VDD100.n362 VDD100.t463 193.183
R12330 VDD100.n365 VDD100.t382 193.183
R12331 VDD100.n368 VDD100.t445 193.183
R12332 VDD100.n401 VDD100.t458 193.183
R12333 VDD100.n403 VDD100.t298 193.183
R12334 VDD100.n406 VDD100.t372 193.183
R12335 VDD100.n409 VDD100.t473 193.183
R12336 VDD100.n33 VDD100.t403 191.288
R12337 VDD100.t375 VDD100.n38 191.288
R12338 VDD100.t113 VDD100.n42 191.288
R12339 VDD100.n44 VDD100.t344 191.288
R12340 VDD100.t245 VDD100.n486 191.288
R12341 VDD100.n487 VDD100.t6 191.288
R12342 VDD100.t115 VDD100.n495 191.288
R12343 VDD100.n496 VDD100.t127 191.288
R12344 VDD100.t222 VDD100.n77 191.288
R12345 VDD100.t430 VDD100.n81 191.288
R12346 VDD100.t232 VDD100.n85 191.288
R12347 VDD100.n329 VDD100.t262 191.288
R12348 VDD100.t363 VDD100.n242 191.288
R12349 VDD100.n244 VDD100.t203 191.288
R12350 VDD100.t257 VDD100.n248 191.288
R12351 VDD100.t399 VDD100.n252 191.288
R12352 VDD100.t350 VDD100.n254 191.288
R12353 VDD100.n256 VDD100.t317 191.288
R12354 VDD100.t420 VDD100.n463 191.288
R12355 VDD100.n464 VDD100.t34 191.288
R12356 VDD100.t194 VDD100.n472 191.288
R12357 VDD100.n473 VDD100.t435 191.288
R12358 VDD100.t237 VDD100.n270 191.288
R12359 VDD100.n271 VDD100.t385 191.288
R12360 VDD100.t352 VDD100.n279 191.288
R12361 VDD100.n280 VDD100.t418 191.288
R12362 VDD100.t357 VDD100.n307 191.288
R12363 VDD100.n308 VDD100.t367 191.288
R12364 VDD100.t365 VDD100.n316 191.288
R12365 VDD100.n317 VDD100.t408 191.288
R12366 VDD100.t422 VDD100.n58 191.288
R12367 VDD100.n59 VDD100.t377 191.288
R12368 VDD100.t192 VDD100.n67 191.288
R12369 VDD100.n68 VDD100.t227 191.288
R12370 VDD100.t111 VDD100.n425 138.095
R12371 VDD100.n426 VDD100.t307 138.095
R12372 VDD100.t330 VDD100.n432 138.095
R12373 VDD100.t270 VDD100.n384 138.095
R12374 VDD100.n385 VDD100.t153 138.095
R12375 VDD100.n396 VDD100.t125 138.095
R12376 VDD100.n395 VDD100.t247 138.095
R12377 VDD100.t328 VDD100.n212 138.095
R12378 VDD100.n213 VDD100.t117 138.095
R12379 VDD100.n355 VDD100.t198 138.095
R12380 VDD100.n354 VDD100.t69 138.095
R12381 VDD100.t346 VDD100.t337 120.755
R12382 VDD100.t292 VDD100.t313 120.755
R12383 VDD100.n33 VDD100.t90 111.743
R12384 VDD100.n38 VDD100.t8 111.743
R12385 VDD100.n42 VDD100.t3 111.743
R12386 VDD100.n44 VDD100.t0 111.743
R12387 VDD100.n486 VDD100.t14 111.743
R12388 VDD100.n487 VDD100.t17 111.743
R12389 VDD100.n495 VDD100.t325 111.743
R12390 VDD100.n496 VDD100.t338 111.743
R12391 VDD100.n77 VDD100.t427 111.743
R12392 VDD100.n81 VDD100.t224 111.743
R12393 VDD100.n85 VDD100.t239 111.743
R12394 VDD100.t11 VDD100.n329 111.743
R12395 VDD100.n242 VDD100.t141 111.743
R12396 VDD100.n244 VDD100.t332 111.743
R12397 VDD100.n248 VDD100.t132 111.743
R12398 VDD100.n252 VDD100.t347 111.743
R12399 VDD100.n254 VDD100.t186 111.743
R12400 VDD100.n256 VDD100.t354 111.743
R12401 VDD100.n463 VDD100.t65 111.743
R12402 VDD100.n464 VDD100.t135 111.743
R12403 VDD100.n472 VDD100.t289 111.743
R12404 VDD100.n473 VDD100.t387 111.743
R12405 VDD100.n270 VDD100.t72 111.743
R12406 VDD100.n271 VDD100.t295 111.743
R12407 VDD100.n279 VDD100.t396 111.743
R12408 VDD100.n280 VDD100.t277 111.743
R12409 VDD100.n307 VDD100.t76 111.743
R12410 VDD100.n308 VDD100.t234 111.743
R12411 VDD100.n316 VDD100.t259 111.743
R12412 VDD100.n317 VDD100.t393 111.743
R12413 VDD100.n58 VDD100.t103 111.743
R12414 VDD100.n59 VDD100.t148 111.743
R12415 VDD100.n67 VDD100.t31 111.743
R12416 VDD100.n68 VDD100.t432 111.743
R12417 VDD100.n172 VDD100.t401 109.849
R12418 VDD100.t51 VDD100.n178 109.849
R12419 VDD100.n179 VDD100.t157 109.849
R12420 VDD100.t155 VDD100.n184 109.849
R12421 VDD100.t144 VDD100.n117 109.849
R12422 VDD100.t55 VDD100.n119 109.849
R12423 VDD100.t196 VDD100.n122 109.849
R12424 VDD100.n125 VDD100.t94 109.849
R12425 VDD100.t44 VDD100.n188 109.849
R12426 VDD100.t20 VDD100.n190 109.849
R12427 VDD100.t293 VDD100.n193 109.849
R12428 VDD100.n196 VDD100.t83 109.849
R12429 VDD100.n347 VDD100.t184 109.849
R12430 VDD100.t214 VDD100.n345 109.849
R12431 VDD100.t456 VDD100.n339 109.849
R12432 VDD100.t146 VDD100.n360 109.849
R12433 VDD100.t39 VDD100.n362 109.849
R12434 VDD100.t106 VDD100.n365 109.849
R12435 VDD100.n368 VDD100.t97 109.849
R12436 VDD100.t62 VDD100.n401 109.849
R12437 VDD100.t272 VDD100.n403 109.849
R12438 VDD100.t335 VDD100.n406 109.849
R12439 VDD100.n409 VDD100.t80 109.849
R12440 VDD100.n436 VDD100.t108 105.66
R12441 VDD100.n230 VDD100.t123 105.66
R12442 VDD100.t108 VDD100.t100 63.3967
R12443 VDD100.t123 VDD100.t86 63.3967
R12444 VDD100.n478 VDD100.t405 62.1896
R12445 VDD100.n246 VDD100.t242 62.1896
R12446 VDD100.n258 VDD100.t424 62.1896
R12447 VDD100.n79 VDD100.t41 61.8817
R12448 VDD100.n83 VDD100.t283 61.8817
R12449 VDD100.t304 VDD100.n87 61.5769
R12450 VDD100.n185 VDD100.t451 59.702
R12451 VDD100.n346 VDD100.t218 59.4064
R12452 VDD100.n340 VDD100.t60 59.4064
R12453 VDD100.n335 VDD100.t159 59.1138
R12454 VDD100.n88 VDD100.t280 55.0852
R12455 VDD100.n90 VDD100.t390 55.0852
R12456 VDD100.n331 VDD100.t121 55.0852
R12457 VDD100.t161 VDD100.n334 55.0852
R12458 VDD100.n434 VDD100.n433 45.2835
R12459 VDD100.n235 VDD100.t86 44.5288
R12460 VDD100.n330 VDD100.n235 44.5288
R12461 VDD100.t100 VDD100.n434 43.7741
R12462 VDD100.n0 VDD100.t89 30.9379
R12463 VDD100.n3 VDD100.t71 30.9379
R12464 VDD100.n126 VDD100.t93 30.9379
R12465 VDD100.n128 VDD100.t96 30.9379
R12466 VDD100.n149 VDD100.t68 30.721
R12467 VDD100.n21 VDD100.t64 30.7204
R12468 VDD100.n9 VDD100.t85 30.7203
R12469 VDD100.n139 VDD100.t99 30.7203
R12470 VDD100.n146 VDD100.t82 30.3459
R12471 VDD100.n15 VDD100.t75 30.2877
R12472 VDD100.n25 VDD100.t102 30.2877
R12473 VDD100.n134 VDD100.t79 30.0062
R12474 VDD100.n25 VDD100.t477 24.9141
R12475 VDD100.n146 VDD100.t485 24.8618
R12476 VDD100.n0 VDD100.t483 24.5101
R12477 VDD100.n14 VDD100.t489 24.5101
R12478 VDD100.n3 VDD100.t492 24.5101
R12479 VDD100.n126 VDD100.t480 24.5101
R12480 VDD100.n128 VDD100.t479 24.5101
R12481 VDD100.n149 VDD100.t490 24.4816
R12482 VDD100.n139 VDD100.t478 24.4814
R12483 VDD100.n9 VDD100.t487 24.4814
R12484 VDD100.n21 VDD100.t481 24.4813
R12485 VDD100.n136 VDD100.t486 24.4392
R12486 VDD100.t337 VDD100.n436 15.0948
R12487 VDD100.n230 VDD100.t292 15.0948
R12488 VDD100 VDD100.t461 10.5649
R12489 VDD100 VDD100.t171 10.5649
R12490 VDD100.n501 VDD100.n500 8.64671
R12491 VDD100.n136 VDD100.n135 8.0005
R12492 VDD100 VDD100.t346 7.80993
R12493 VDD100.t313 VDD100 7.80993
R12494 VDD100.n29 VDD100.n28 6.39761
R12495 VDD100.n156 VDD100.n155 6.39748
R12496 VDD100.n436 VDD100 6.30126
R12497 VDD100 VDD100.n230 6.30126
R12498 VDD100.n160 VDD100.n125 6.3005
R12499 VDD100.n163 VDD100.n122 6.3005
R12500 VDD100.n166 VDD100.n119 6.3005
R12501 VDD100.n169 VDD100.n117 6.3005
R12502 VDD100.n184 VDD100.n183 6.3005
R12503 VDD100.n180 VDD100.n179 6.3005
R12504 VDD100.n178 VDD100.n177 6.3005
R12505 VDD100.n173 VDD100.n172 6.3005
R12506 VDD100.n197 VDD100.n196 6.3005
R12507 VDD100.n200 VDD100.n193 6.3005
R12508 VDD100.n203 VDD100.n190 6.3005
R12509 VDD100.n206 VDD100.n188 6.3005
R12510 VDD100.n270 VDD100.n269 6.3005
R12511 VDD100.n272 VDD100.n271 6.3005
R12512 VDD100.n279 VDD100.n278 6.3005
R12513 VDD100.n281 VDD100.n280 6.3005
R12514 VDD100.n294 VDD100.n248 6.3005
R12515 VDD100.n291 VDD100.n252 6.3005
R12516 VDD100.n288 VDD100.n254 6.3005
R12517 VDD100.n285 VDD100.n256 6.3005
R12518 VDD100.n307 VDD100.n306 6.3005
R12519 VDD100.n309 VDD100.n308 6.3005
R12520 VDD100.n316 VDD100.n315 6.3005
R12521 VDD100.n318 VDD100.n317 6.3005
R12522 VDD100.n329 VDD100.n328 6.3005
R12523 VDD100.n325 VDD100.n242 6.3005
R12524 VDD100.n322 VDD100.n244 6.3005
R12525 VDD100.n235 VDD100.n234 6.3005
R12526 VDD100 VDD100.n331 6.3005
R12527 VDD100.n334 VDD100.n333 6.3005
R12528 VDD100.n339 VDD100.n338 6.3005
R12529 VDD100.n345 VDD100.n344 6.3005
R12530 VDD100.n348 VDD100.n347 6.3005
R12531 VDD100.n354 VDD100.n353 6.3005
R12532 VDD100.n355 VDD100.n217 6.3005
R12533 VDD100.n214 VDD100.n213 6.3005
R12534 VDD100.n212 VDD100.n211 6.3005
R12535 VDD100.n369 VDD100.n368 6.3005
R12536 VDD100.n372 VDD100.n365 6.3005
R12537 VDD100.n375 VDD100.n362 6.3005
R12538 VDD100.n378 VDD100.n360 6.3005
R12539 VDD100.n395 VDD100.n394 6.3005
R12540 VDD100.n396 VDD100.n389 6.3005
R12541 VDD100.n386 VDD100.n385 6.3005
R12542 VDD100.n384 VDD100.n383 6.3005
R12543 VDD100.n410 VDD100.n409 6.3005
R12544 VDD100.n413 VDD100.n406 6.3005
R12545 VDD100.n416 VDD100.n403 6.3005
R12546 VDD100.n419 VDD100.n401 6.3005
R12547 VDD100.n432 VDD100.n431 6.3005
R12548 VDD100.n427 VDD100.n426 6.3005
R12549 VDD100.n425 VDD100.n424 6.3005
R12550 VDD100.n440 VDD100.n434 6.3005
R12551 VDD100 VDD100.n90 6.3005
R12552 VDD100.n443 VDD100.n88 6.3005
R12553 VDD100.n448 VDD100.n85 6.3005
R12554 VDD100.n452 VDD100.n81 6.3005
R12555 VDD100.n456 VDD100.n77 6.3005
R12556 VDD100.n463 VDD100.n462 6.3005
R12557 VDD100.n465 VDD100.n464 6.3005
R12558 VDD100.n472 VDD100.n471 6.3005
R12559 VDD100.n474 VDD100.n473 6.3005
R12560 VDD100.n58 VDD100.n57 6.3005
R12561 VDD100.n60 VDD100.n59 6.3005
R12562 VDD100.n67 VDD100.n66 6.3005
R12563 VDD100.n69 VDD100.n68 6.3005
R12564 VDD100.n486 VDD100.n485 6.3005
R12565 VDD100.n488 VDD100.n487 6.3005
R12566 VDD100.n495 VDD100.n494 6.3005
R12567 VDD100.n497 VDD100.n496 6.3005
R12568 VDD100.n34 VDD100.n33 6.3005
R12569 VDD100.n510 VDD100.n38 6.3005
R12570 VDD100.n507 VDD100.n42 6.3005
R12571 VDD100.n504 VDD100.n44 6.3005
R12572 VDD100.n18 VDD100.n17 5.30733
R12573 VDD100.n145 VDD100.n144 5.30657
R12574 VDD100.n197 VDD100.t84 5.213
R12575 VDD100.n269 VDD100.n265 5.213
R12576 VDD100.n306 VDD100.n302 5.213
R12577 VDD100.n369 VDD100.t98 5.213
R12578 VDD100.n410 VDD100.t81 5.213
R12579 VDD100.n57 VDD100.n53 5.213
R12580 VDD100 VDD100.t469 5.16454
R12581 VDD100 VDD100.n229 5.16369
R12582 VDD100.n226 VDD100.t162 5.14212
R12583 VDD100.n445 VDD100.n444 5.14212
R12584 VDD100.n511 VDD100.n37 5.13287
R12585 VDD100.n508 VDD100.n41 5.13287
R12586 VDD100.n506 VDD100.t114 5.13287
R12587 VDD100.n505 VDD100.n43 5.13287
R12588 VDD100.n503 VDD100.t345 5.13287
R12589 VDD100.n73 VDD100.n72 5.13287
R12590 VDD100.n459 VDD100.n458 5.13287
R12591 VDD100.n466 VDD100.t35 5.13287
R12592 VDD100.n467 VDD100.n71 5.13287
R12593 VDD100.n470 VDD100.t195 5.13287
R12594 VDD100.n469 VDD100.n468 5.13287
R12595 VDD100.n475 VDD100.t436 5.13287
R12596 VDD100.n438 VDD100.t101 5.13287
R12597 VDD100.n109 VDD100.t156 5.13287
R12598 VDD100.n181 VDD100.t158 5.13287
R12599 VDD100.n113 VDD100.n112 5.13287
R12600 VDD100.n176 VDD100.t52 5.13287
R12601 VDD100.n175 VDD100.n114 5.13287
R12602 VDD100.n174 VDD100.t402 5.13287
R12603 VDD100.n171 VDD100.n115 5.13287
R12604 VDD100.n162 VDD100.t197 5.13287
R12605 VDD100.n165 VDD100.t56 5.13287
R12606 VDD100.n167 VDD100.n118 5.13287
R12607 VDD100.n168 VDD100.t145 5.13287
R12608 VDD100.n170 VDD100.n116 5.13287
R12609 VDD100.n199 VDD100.t294 5.13287
R12610 VDD100.n202 VDD100.t21 5.13287
R12611 VDD100.n204 VDD100.n189 5.13287
R12612 VDD100.n205 VDD100.t45 5.13287
R12613 VDD100.n207 VDD100.n187 5.13287
R12614 VDD100.n232 VDD100.n228 5.13287
R12615 VDD100.n264 VDD100.n263 5.13287
R12616 VDD100.n274 VDD100.n260 5.13287
R12617 VDD100.n277 VDD100.t353 5.13287
R12618 VDD100.n276 VDD100.n275 5.13287
R12619 VDD100.n282 VDD100.t419 5.13287
R12620 VDD100.n295 VDD100.n247 5.13287
R12621 VDD100.n292 VDD100.n251 5.13287
R12622 VDD100.n290 VDD100.t400 5.13287
R12623 VDD100.n289 VDD100.n253 5.13287
R12624 VDD100.n287 VDD100.t351 5.13287
R12625 VDD100.n286 VDD100.n255 5.13287
R12626 VDD100.n284 VDD100.t318 5.13287
R12627 VDD100.n301 VDD100.n300 5.13287
R12628 VDD100.n311 VDD100.n297 5.13287
R12629 VDD100.n314 VDD100.t366 5.13287
R12630 VDD100.n313 VDD100.n312 5.13287
R12631 VDD100.n319 VDD100.t409 5.13287
R12632 VDD100.n240 VDD100.n236 5.13287
R12633 VDD100.n327 VDD100.t263 5.13287
R12634 VDD100.n326 VDD100.n241 5.13287
R12635 VDD100.n324 VDD100.t364 5.13287
R12636 VDD100.n323 VDD100.n243 5.13287
R12637 VDD100.n321 VDD100.t204 5.13287
R12638 VDD100.n224 VDD100.t457 5.13287
R12639 VDD100.n337 VDD100.n225 5.13287
R12640 VDD100.n343 VDD100.t215 5.13287
R12641 VDD100.n342 VDD100.n223 5.13287
R12642 VDD100.n349 VDD100.t185 5.13287
R12643 VDD100.n221 VDD100.n220 5.13287
R12644 VDD100.n104 VDD100.t70 5.13287
R12645 VDD100.n350 VDD100.t199 5.13287
R12646 VDD100.n216 VDD100.n105 5.13287
R12647 VDD100.n215 VDD100.t118 5.13287
R12648 VDD100.n107 VDD100.n106 5.13287
R12649 VDD100.n210 VDD100.t329 5.13287
R12650 VDD100.n209 VDD100.n108 5.13287
R12651 VDD100.n371 VDD100.t107 5.13287
R12652 VDD100.n374 VDD100.t40 5.13287
R12653 VDD100.n376 VDD100.n361 5.13287
R12654 VDD100.n377 VDD100.t147 5.13287
R12655 VDD100.n379 VDD100.n359 5.13287
R12656 VDD100.n99 VDD100.t248 5.13287
R12657 VDD100.n392 VDD100.t126 5.13287
R12658 VDD100.n388 VDD100.n100 5.13287
R12659 VDD100.n387 VDD100.t154 5.13287
R12660 VDD100.n102 VDD100.n101 5.13287
R12661 VDD100.n382 VDD100.t271 5.13287
R12662 VDD100.n381 VDD100.n103 5.13287
R12663 VDD100.n412 VDD100.t336 5.13287
R12664 VDD100.n415 VDD100.t273 5.13287
R12665 VDD100.n417 VDD100.n402 5.13287
R12666 VDD100.n418 VDD100.t63 5.13287
R12667 VDD100.n420 VDD100.n400 5.13287
R12668 VDD100.n430 VDD100.t331 5.13287
R12669 VDD100.n429 VDD100.n95 5.13287
R12670 VDD100.n428 VDD100.t308 5.13287
R12671 VDD100.n97 VDD100.n96 5.13287
R12672 VDD100.n423 VDD100.t112 5.13287
R12673 VDD100.n422 VDD100.n98 5.13287
R12674 VDD100.n449 VDD100.n84 5.13287
R12675 VDD100.n447 VDD100.t233 5.13287
R12676 VDD100.n453 VDD100.n80 5.13287
R12677 VDD100.n451 VDD100.t431 5.13287
R12678 VDD100.n457 VDD100.n76 5.13287
R12679 VDD100.n455 VDD100.t223 5.13287
R12680 VDD100.n52 VDD100.n51 5.13287
R12681 VDD100.n62 VDD100.n48 5.13287
R12682 VDD100.n65 VDD100.t193 5.13287
R12683 VDD100.n64 VDD100.n63 5.13287
R12684 VDD100.n70 VDD100.t228 5.13287
R12685 VDD100.n479 VDD100.n46 5.13287
R12686 VDD100.n483 VDD100.n482 5.13287
R12687 VDD100.n489 VDD100.t7 5.13287
R12688 VDD100.n490 VDD100.n45 5.13287
R12689 VDD100.n493 VDD100.t116 5.13287
R12690 VDD100.n492 VDD100.n491 5.13287
R12691 VDD100.n498 VDD100.t128 5.13287
R12692 VDD100 VDD100.n499 5.1189
R12693 VDD100.n332 VDD100.t122 5.09693
R12694 VDD100.n442 VDD100.n89 5.09693
R12695 VDD100.n186 VDD100.t452 5.09407
R12696 VDD100.n259 VDD100.n257 5.09407
R12697 VDD100.n296 VDD100.n245 5.09407
R12698 VDD100.n336 VDD100.t160 5.09407
R12699 VDD100.n341 VDD100.t61 5.09407
R12700 VDD100.n222 VDD100.t219 5.09407
R12701 VDD100.n358 VDD100.t172 5.09407
R12702 VDD100.n399 VDD100.t462 5.09407
R12703 VDD100.n446 VDD100.n86 5.09407
R12704 VDD100.n450 VDD100.n82 5.09407
R12705 VDD100.n454 VDD100.n78 5.09407
R12706 VDD100.n477 VDD100.n47 5.09407
R12707 VDD100.n32 VDD100.n31 4.8755
R12708 VDD100.n159 VDD100.t95 4.8755
R12709 VDD100.n28 VDD100.n18 4.84121
R12710 VDD100.n155 VDD100.n145 4.84121
R12711 VDD100.n137 VDD100.n136 4.5005
R12712 VDD100.n140 VDD100.n138 4.5005
R12713 VDD100.n141 VDD100.n138 4.5005
R12714 VDD100.n129 VDD100.n127 4.5005
R12715 VDD100.n130 VDD100.n127 4.5005
R12716 VDD100.n150 VDD100.n148 4.5005
R12717 VDD100.n151 VDD100.n148 4.5005
R12718 VDD100.n437 VDD100 4.40201
R12719 VDD100.n231 VDD100 4.40201
R12720 VDD100.n502 VDD100 4.04877
R12721 VDD100 VDD100.n501 3.99616
R12722 VDD100.n439 VDD100.n435 3.94862
R12723 VDD100.n233 VDD100.t124 3.94862
R12724 VDD100.n134 VDD100.n133 3.61662
R12725 VDD100.n231 VDD100 3.52487
R12726 VDD100.n437 VDD100 3.47987
R12727 VDD100.n29 VDD100.n0 2.88198
R12728 VDD100.n156 VDD100.n126 2.88182
R12729 VDD100.n239 VDD100.n238 2.88011
R12730 VDD100.n93 VDD100.n92 2.87966
R12731 VDD100.n512 VDD100.n36 2.85787
R12732 VDD100.n509 VDD100.n40 2.85787
R12733 VDD100.n461 VDD100.n75 2.85787
R12734 VDD100.n182 VDD100.n111 2.85787
R12735 VDD100.n161 VDD100.n124 2.85787
R12736 VDD100.n164 VDD100.n121 2.85787
R12737 VDD100.n198 VDD100.n195 2.85787
R12738 VDD100.n201 VDD100.n192 2.85787
R12739 VDD100.n268 VDD100.n267 2.85787
R12740 VDD100.n273 VDD100.n262 2.85787
R12741 VDD100.n293 VDD100.n250 2.85787
R12742 VDD100.n305 VDD100.n304 2.85787
R12743 VDD100.n310 VDD100.n299 2.85787
R12744 VDD100.n352 VDD100.n219 2.85787
R12745 VDD100.n370 VDD100.n367 2.85787
R12746 VDD100.n373 VDD100.n364 2.85787
R12747 VDD100.n393 VDD100.n391 2.85787
R12748 VDD100.n411 VDD100.n408 2.85787
R12749 VDD100.n414 VDD100.n405 2.85787
R12750 VDD100.n56 VDD100.n55 2.85787
R12751 VDD100.n61 VDD100.n50 2.85787
R12752 VDD100.n484 VDD100.n481 2.85787
R12753 VDD100.n36 VDD100.t404 2.2755
R12754 VDD100.n36 VDD100.n35 2.2755
R12755 VDD100.n40 VDD100.t376 2.2755
R12756 VDD100.n40 VDD100.n39 2.2755
R12757 VDD100.n75 VDD100.t421 2.2755
R12758 VDD100.n75 VDD100.n74 2.2755
R12759 VDD100.n92 VDD100.t411 2.2755
R12760 VDD100.n92 VDD100.n91 2.2755
R12761 VDD100.n111 VDD100.t250 2.2755
R12762 VDD100.n111 VDD100.n110 2.2755
R12763 VDD100.n124 VDD100.t312 2.2755
R12764 VDD100.n124 VDD100.n123 2.2755
R12765 VDD100.n121 VDD100.t54 2.2755
R12766 VDD100.n121 VDD100.n120 2.2755
R12767 VDD100.n195 VDD100.t217 2.2755
R12768 VDD100.n195 VDD100.n194 2.2755
R12769 VDD100.n192 VDD100.t120 2.2755
R12770 VDD100.n192 VDD100.n191 2.2755
R12771 VDD100.n238 VDD100.t360 2.2755
R12772 VDD100.n238 VDD100.n237 2.2755
R12773 VDD100.n267 VDD100.t238 2.2755
R12774 VDD100.n267 VDD100.n266 2.2755
R12775 VDD100.n262 VDD100.t386 2.2755
R12776 VDD100.n262 VDD100.n261 2.2755
R12777 VDD100.n250 VDD100.t258 2.2755
R12778 VDD100.n250 VDD100.n249 2.2755
R12779 VDD100.n304 VDD100.t358 2.2755
R12780 VDD100.n304 VDD100.n303 2.2755
R12781 VDD100.n299 VDD100.t368 2.2755
R12782 VDD100.n299 VDD100.n298 2.2755
R12783 VDD100.n219 VDD100.t47 2.2755
R12784 VDD100.n219 VDD100.n218 2.2755
R12785 VDD100.n367 VDD100.t180 2.2755
R12786 VDD100.n367 VDD100.n366 2.2755
R12787 VDD100.n364 VDD100.t152 2.2755
R12788 VDD100.n364 VDD100.n363 2.2755
R12789 VDD100.n391 VDD100.t164 2.2755
R12790 VDD100.n391 VDD100.n390 2.2755
R12791 VDD100.n408 VDD100.t444 2.2755
R12792 VDD100.n408 VDD100.n407 2.2755
R12793 VDD100.n405 VDD100.t310 2.2755
R12794 VDD100.n405 VDD100.n404 2.2755
R12795 VDD100.n55 VDD100.t423 2.2755
R12796 VDD100.n55 VDD100.n54 2.2755
R12797 VDD100.n50 VDD100.t378 2.2755
R12798 VDD100.n50 VDD100.n49 2.2755
R12799 VDD100.n481 VDD100.t246 2.2755
R12800 VDD100.n481 VDD100.n480 2.2755
R12801 VDD100.n12 VDD100.n11 2.2439
R12802 VDD100.n24 VDD100.n23 2.2439
R12803 VDD100.n143 VDD100.n142 2.2439
R12804 VDD100.n153 VDD100.n152 2.2439
R12805 VDD100.n6 VDD100.n5 2.24362
R12806 VDD100.n132 VDD100.n131 2.24362
R12807 VDD100.n4 VDD100.n3 2.12269
R12808 VDD100.n129 VDD100.n128 2.12257
R12809 VDD100.n16 VDD100.n15 1.82213
R12810 VDD100.n26 VDD100.n25 1.82213
R12811 VDD100 VDD100.n73 1.81843
R12812 VDD100 VDD100.n295 1.81843
R12813 VDD100 VDD100.n449 1.81843
R12814 VDD100 VDD100.n453 1.81843
R12815 VDD100.n479 VDD100 1.81843
R12816 VDD100.n147 VDD100.n146 1.81789
R12817 VDD100 VDD100.n109 1.77285
R12818 VDD100 VDD100.n224 1.77285
R12819 VDD100.n343 VDD100 1.77285
R12820 VDD100 VDD100.n104 1.77285
R12821 VDD100 VDD100.n99 1.77285
R12822 VDD100.n144 VDD100.n143 1.62565
R12823 VDD100.n154 VDD100.n153 1.62565
R12824 VDD100.n27 VDD100.n24 1.6239
R12825 VDD100.n17 VDD100.n12 1.6239
R12826 VDD100.n22 VDD100.n21 1.39892
R12827 VDD100.n10 VDD100.n9 1.3985
R12828 VDD100.n150 VDD100.n149 1.39782
R12829 VDD100.n140 VDD100.n139 1.39728
R12830 VDD100.n171 VDD100.n170 1.16167
R12831 VDD100.n17 VDD100.n16 1.12224
R12832 VDD100.n144 VDD100.n137 1.12171
R12833 VDD100.n154 VDD100.n147 1.12171
R12834 VDD100.n27 VDD100.n26 1.12167
R12835 VDD100.n502 VDD100.n498 1.12044
R12836 VDD100.n208 VDD100.n207 1.07428
R12837 VDD100.n380 VDD100.n379 1.07428
R12838 VDD100.n421 VDD100.n420 1.07428
R12839 VDD100.n283 VDD100.n282 1.0737
R12840 VDD100.n320 VDD100.n319 1.0737
R12841 VDD100.n476 VDD100.n70 1.0737
R12842 VDD100.n136 VDD100.n134 0.840632
R12843 VDD100.n460 VDD100.n457 0.715235
R12844 VDD100.n32 VDD100.n30 0.603658
R12845 VDD100.n28 VDD100.n27 0.523557
R12846 VDD100.n155 VDD100.n154 0.5228
R12847 VDD100.n18 VDD100.n6 0.497812
R12848 VDD100.n145 VDD100.n132 0.497812
R12849 VDD100 VDD100.n349 0.434967
R12850 VDD100.n15 VDD100.n14 0.404541
R12851 VDD100 VDD100.n441 0.339236
R12852 VDD100 VDD100.n227 0.338387
R12853 VDD100.n34 VDD100.n32 0.337997
R12854 VDD100.n160 VDD100.n159 0.337997
R12855 VDD100 VDD100.n226 0.334577
R12856 VDD100 VDD100.n445 0.334577
R12857 VDD100.n159 VDD100.n158 0.333658
R12858 VDD100.n443 VDD100.n442 0.318198
R12859 VDD100.n333 VDD100.n332 0.317357
R12860 VDD100.n351 VDD100 0.280768
R12861 VDD100.n165 VDD100.n164 0.233919
R12862 VDD100.n162 VDD100.n161 0.233919
R12863 VDD100.n202 VDD100.n201 0.233919
R12864 VDD100.n199 VDD100.n198 0.233919
R12865 VDD100.n268 VDD100.n264 0.233919
R12866 VDD100.n274 VDD100.n273 0.233919
R12867 VDD100.n305 VDD100.n301 0.233919
R12868 VDD100.n311 VDD100.n310 0.233919
R12869 VDD100.n374 VDD100.n373 0.233919
R12870 VDD100.n371 VDD100.n370 0.233919
R12871 VDD100.n415 VDD100.n414 0.233919
R12872 VDD100.n412 VDD100.n411 0.233919
R12873 VDD100.n56 VDD100.n52 0.233919
R12874 VDD100.n62 VDD100.n61 0.233919
R12875 VDD100.n512 VDD100.n511 0.233919
R12876 VDD100.n509 VDD100.n508 0.233919
R12877 VDD100.n447 VDD100.n446 0.170499
R12878 VDD100.n451 VDD100.n450 0.170499
R12879 VDD100.n455 VDD100.n454 0.170499
R12880 VDD100.n337 VDD100.n336 0.170231
R12881 VDD100.n342 VDD100.n341 0.170231
R12882 VDD100.n222 VDD100.n221 0.170231
R12883 VDD100.n501 VDD100 0.166174
R12884 VDD100.n332 VDD100 0.147133
R12885 VDD100.n442 VDD100 0.146292
R12886 VDD100.n284 VDD100.n283 0.143967
R12887 VDD100.n321 VDD100.n320 0.143967
R12888 VDD100.n476 VDD100.n475 0.143967
R12889 VDD100.n209 VDD100.n208 0.143501
R12890 VDD100.n381 VDD100.n380 0.143501
R12891 VDD100.n422 VDD100.n421 0.143501
R12892 VDD100.n168 VDD100.n167 0.141016
R12893 VDD100.n175 VDD100.n174 0.141016
R12894 VDD100.n176 VDD100.n113 0.141016
R12895 VDD100.n205 VDD100.n204 0.141016
R12896 VDD100.n277 VDD100.n276 0.141016
R12897 VDD100.n290 VDD100.n289 0.141016
R12898 VDD100.n287 VDD100.n286 0.141016
R12899 VDD100.n314 VDD100.n313 0.141016
R12900 VDD100.n327 VDD100.n326 0.141016
R12901 VDD100.n324 VDD100.n323 0.141016
R12902 VDD100.n210 VDD100.n107 0.141016
R12903 VDD100.n216 VDD100.n215 0.141016
R12904 VDD100.n377 VDD100.n376 0.141016
R12905 VDD100.n382 VDD100.n102 0.141016
R12906 VDD100.n388 VDD100.n387 0.141016
R12907 VDD100.n418 VDD100.n417 0.141016
R12908 VDD100.n423 VDD100.n97 0.141016
R12909 VDD100.n429 VDD100.n428 0.141016
R12910 VDD100.n467 VDD100.n466 0.141016
R12911 VDD100.n470 VDD100.n469 0.141016
R12912 VDD100.n65 VDD100.n64 0.141016
R12913 VDD100.n490 VDD100.n489 0.141016
R12914 VDD100.n493 VDD100.n492 0.141016
R12915 VDD100.n506 VDD100.n505 0.141016
R12916 VDD100.n283 VDD100.n259 0.139745
R12917 VDD100.n477 VDD100.n476 0.139745
R12918 VDD100.n208 VDD100.n186 0.138896
R12919 VDD100.n380 VDD100.n358 0.138896
R12920 VDD100 VDD100.n296 0.128708
R12921 VDD100 VDD100.n399 0.127858
R12922 VDD100 VDD100.n292 0.123016
R12923 VDD100.n240 VDD100 0.123016
R12924 VDD100 VDD100.n483 0.123016
R12925 VDD100 VDD100.n181 0.122435
R12926 VDD100 VDD100.n392 0.122435
R12927 VDD100.n430 VDD100 0.122435
R12928 VDD100.n26 VDD100 0.112066
R12929 VDD100.n182 VDD100 0.111984
R12930 VDD100.n352 VDD100 0.111984
R12931 VDD100.n393 VDD100 0.111984
R12932 VDD100.n30 VDD100 0.111564
R12933 VDD100.n293 VDD100 0.111403
R12934 VDD100.n461 VDD100 0.111403
R12935 VDD100.n484 VDD100 0.111403
R12936 VDD100.n147 VDD100 0.110941
R12937 VDD100 VDD100.n93 0.108832
R12938 VDD100 VDD100.n239 0.108613
R12939 VDD100.n170 VDD100.n169 0.107339
R12940 VDD100.n167 VDD100.n166 0.107339
R12941 VDD100.n173 VDD100.n171 0.107339
R12942 VDD100.n177 VDD100.n175 0.107339
R12943 VDD100.n180 VDD100.n113 0.107339
R12944 VDD100.n207 VDD100.n206 0.107339
R12945 VDD100.n204 VDD100.n203 0.107339
R12946 VDD100.n278 VDD100.n277 0.107339
R12947 VDD100.n282 VDD100.n281 0.107339
R12948 VDD100.n291 VDD100.n290 0.107339
R12949 VDD100.n288 VDD100.n287 0.107339
R12950 VDD100.n285 VDD100.n284 0.107339
R12951 VDD100.n315 VDD100.n314 0.107339
R12952 VDD100.n319 VDD100.n318 0.107339
R12953 VDD100.n328 VDD100.n327 0.107339
R12954 VDD100.n325 VDD100.n324 0.107339
R12955 VDD100.n322 VDD100.n321 0.107339
R12956 VDD100.n338 VDD100.n337 0.107339
R12957 VDD100.n344 VDD100.n342 0.107339
R12958 VDD100.n348 VDD100.n221 0.107339
R12959 VDD100.n211 VDD100.n209 0.107339
R12960 VDD100.n214 VDD100.n107 0.107339
R12961 VDD100.n217 VDD100.n216 0.107339
R12962 VDD100.n379 VDD100.n378 0.107339
R12963 VDD100.n376 VDD100.n375 0.107339
R12964 VDD100.n383 VDD100.n381 0.107339
R12965 VDD100.n386 VDD100.n102 0.107339
R12966 VDD100.n389 VDD100.n388 0.107339
R12967 VDD100.n420 VDD100.n419 0.107339
R12968 VDD100.n417 VDD100.n416 0.107339
R12969 VDD100.n424 VDD100.n422 0.107339
R12970 VDD100.n427 VDD100.n97 0.107339
R12971 VDD100.n431 VDD100.n429 0.107339
R12972 VDD100.n448 VDD100.n447 0.107339
R12973 VDD100.n452 VDD100.n451 0.107339
R12974 VDD100.n456 VDD100.n455 0.107339
R12975 VDD100.n466 VDD100.n465 0.107339
R12976 VDD100.n471 VDD100.n470 0.107339
R12977 VDD100.n475 VDD100.n474 0.107339
R12978 VDD100.n66 VDD100.n65 0.107339
R12979 VDD100.n70 VDD100.n69 0.107339
R12980 VDD100.n489 VDD100.n488 0.107339
R12981 VDD100.n494 VDD100.n493 0.107339
R12982 VDD100.n498 VDD100.n497 0.107339
R12983 VDD100.n507 VDD100.n506 0.107339
R12984 VDD100.n504 VDD100.n503 0.107339
R12985 VDD100 VDD100.n268 0.106758
R12986 VDD100.n273 VDD100 0.106758
R12987 VDD100 VDD100.n293 0.106758
R12988 VDD100 VDD100.n305 0.106758
R12989 VDD100.n310 VDD100 0.106758
R12990 VDD100 VDD100.n461 0.106758
R12991 VDD100 VDD100.n56 0.106758
R12992 VDD100.n61 VDD100 0.106758
R12993 VDD100 VDD100.n484 0.106758
R12994 VDD100 VDD100.n512 0.106758
R12995 VDD100 VDD100.n509 0.106758
R12996 VDD100.n164 VDD100 0.106177
R12997 VDD100.n161 VDD100 0.106177
R12998 VDD100 VDD100.n182 0.106177
R12999 VDD100.n201 VDD100 0.106177
R13000 VDD100.n198 VDD100 0.106177
R13001 VDD100 VDD100.n352 0.106177
R13002 VDD100.n373 VDD100 0.106177
R13003 VDD100.n370 VDD100 0.106177
R13004 VDD100 VDD100.n393 0.106177
R13005 VDD100.n414 VDD100 0.106177
R13006 VDD100.n411 VDD100 0.106177
R13007 VDD100.n13 VDD100 0.0850665
R13008 VDD100.n135 VDD100 0.0839415
R13009 VDD100 VDD100.n460 0.0829516
R13010 VDD100 VDD100.n351 0.082371
R13011 VDD100.n8 VDD100 0.0816915
R13012 VDD100.n141 VDD100 0.0816915
R13013 VDD100.n163 VDD100.n162 0.080629
R13014 VDD100.n183 VDD100.n109 0.080629
R13015 VDD100.n200 VDD100.n199 0.080629
R13016 VDD100.n272 VDD100.n264 0.080629
R13017 VDD100.n295 VDD100.n294 0.080629
R13018 VDD100.n309 VDD100.n301 0.080629
R13019 VDD100.n353 VDD100.n104 0.080629
R13020 VDD100.n372 VDD100.n371 0.080629
R13021 VDD100.n394 VDD100.n99 0.080629
R13022 VDD100.n413 VDD100.n412 0.080629
R13023 VDD100.n462 VDD100.n73 0.080629
R13024 VDD100.n60 VDD100.n52 0.080629
R13025 VDD100.n485 VDD100.n479 0.080629
R13026 VDD100.n511 VDD100.n510 0.080629
R13027 VDD100.n20 VDD100 0.0805665
R13028 VDD100.n151 VDD100 0.0805665
R13029 VDD100 VDD100.n168 0.0794677
R13030 VDD100 VDD100.n165 0.0794677
R13031 VDD100.n174 VDD100 0.0794677
R13032 VDD100 VDD100.n176 0.0794677
R13033 VDD100.n181 VDD100 0.0794677
R13034 VDD100 VDD100.n205 0.0794677
R13035 VDD100 VDD100.n202 0.0794677
R13036 VDD100 VDD100.n210 0.0794677
R13037 VDD100.n215 VDD100 0.0794677
R13038 VDD100.n350 VDD100 0.0794677
R13039 VDD100 VDD100.n377 0.0794677
R13040 VDD100 VDD100.n374 0.0794677
R13041 VDD100 VDD100.n382 0.0794677
R13042 VDD100.n387 VDD100 0.0794677
R13043 VDD100.n392 VDD100 0.0794677
R13044 VDD100 VDD100.n418 0.0794677
R13045 VDD100 VDD100.n415 0.0794677
R13046 VDD100 VDD100.n423 0.0794677
R13047 VDD100.n428 VDD100 0.0794677
R13048 VDD100 VDD100.n430 0.0794677
R13049 VDD100 VDD100.n226 0.0794623
R13050 VDD100.n445 VDD100 0.0794623
R13051 VDD100 VDD100.n274 0.0788871
R13052 VDD100.n276 VDD100 0.0788871
R13053 VDD100.n292 VDD100 0.0788871
R13054 VDD100.n289 VDD100 0.0788871
R13055 VDD100.n286 VDD100 0.0788871
R13056 VDD100 VDD100.n311 0.0788871
R13057 VDD100.n313 VDD100 0.0788871
R13058 VDD100 VDD100.n240 0.0788871
R13059 VDD100.n326 VDD100 0.0788871
R13060 VDD100.n323 VDD100 0.0788871
R13061 VDD100.n459 VDD100 0.0788871
R13062 VDD100 VDD100.n467 0.0788871
R13063 VDD100.n469 VDD100 0.0788871
R13064 VDD100 VDD100.n62 0.0788871
R13065 VDD100.n64 VDD100 0.0788871
R13066 VDD100.n483 VDD100 0.0788871
R13067 VDD100 VDD100.n490 0.0788871
R13068 VDD100.n492 VDD100 0.0788871
R13069 VDD100.n508 VDD100 0.0788871
R13070 VDD100.n505 VDD100 0.0788871
R13071 VDD100 VDD100.n224 0.0759839
R13072 VDD100 VDD100.n343 0.0759839
R13073 VDD100.n349 VDD100 0.0759839
R13074 VDD100.n449 VDD100 0.0754032
R13075 VDD100.n453 VDD100 0.0754032
R13076 VDD100.n457 VDD100 0.0754032
R13077 VDD100.n2 VDD100 0.0749415
R13078 VDD100.n130 VDD100 0.0738165
R13079 VDD100.n158 VDD100.n156 0.0725
R13080 VDD100.n186 VDD100 0.0709717
R13081 VDD100.n336 VDD100 0.0709717
R13082 VDD100.n341 VDD100 0.0709717
R13083 VDD100 VDD100.n222 0.0709717
R13084 VDD100.n358 VDD100 0.0709717
R13085 VDD100.n399 VDD100 0.0709717
R13086 VDD100.n259 VDD100 0.0701226
R13087 VDD100.n296 VDD100 0.0701226
R13088 VDD100.n446 VDD100 0.0701226
R13089 VDD100.n450 VDD100 0.0701226
R13090 VDD100.n454 VDD100 0.0701226
R13091 VDD100 VDD100.n477 0.0701226
R13092 VDD100.n157 VDD100 0.0700455
R13093 VDD100 VDD100.n227 0.0491131
R13094 VDD100.n441 VDD100 0.0487847
R13095 VDD100.n158 VDD100.n157 0.0455
R13096 VDD100.n232 VDD100.n231 0.0409015
R13097 VDD100.n438 VDD100.n437 0.040573
R13098 VDD100.n351 VDD100.n350 0.0405645
R13099 VDD100.n460 VDD100.n459 0.0405645
R13100 VDD100.n503 VDD100.n502 0.0405645
R13101 VDD100.n30 VDD100.n29 0.0344889
R13102 VDD100.n11 VDD100.n8 0.0275
R13103 VDD100.n16 VDD100.n13 0.0275
R13104 VDD100.n142 VDD100.n141 0.0275
R13105 VDD100.n135 VDD100.n133 0.0275
R13106 VDD100.n23 VDD100.n20 0.026375
R13107 VDD100.n152 VDD100.n151 0.026375
R13108 VDD100.n12 VDD100.n7 0.025705
R13109 VDD100.n24 VDD100.n19 0.025705
R13110 VDD100.n143 VDD100.n138 0.025705
R13111 VDD100.n153 VDD100.n148 0.025705
R13112 VDD100.n233 VDD100.n232 0.025135
R13113 VDD100.n439 VDD100.n438 0.025135
R13114 VDD100.n234 VDD100.n233 0.0211934
R13115 VDD100.n440 VDD100.n439 0.0211934
R13116 VDD100.n131 VDD100.n130 0.02075
R13117 VDD100.n5 VDD100.n2 0.019625
R13118 VDD100.n6 VDD100.n1 0.0169383
R13119 VDD100.n132 VDD100.n127 0.0169383
R13120 VDD100.n441 VDD100.n93 0.0132147
R13121 VDD100.n239 VDD100.n227 0.0131133
R13122 VDD100.n320 VDD100 0.0115377
R13123 VDD100.n421 VDD100 0.0115377
R13124 VDD100.n5 VDD100.n4 0.010625
R13125 VDD100.n131 VDD100.n129 0.0095
R13126 VDD100 VDD100.n448 0.00572581
R13127 VDD100 VDD100.n452 0.00572581
R13128 VDD100 VDD100.n456 0.00572581
R13129 VDD100.n338 VDD100 0.00514516
R13130 VDD100.n344 VDD100 0.00514516
R13131 VDD100 VDD100.n348 0.00514516
R13132 VDD100.n157 VDD100 0.00459091
R13133 VDD100.n23 VDD100.n22 0.003875
R13134 VDD100.n152 VDD100.n150 0.003875
R13135 VDD100.n11 VDD100.n10 0.00275
R13136 VDD100.n142 VDD100.n140 0.00275
R13137 VDD100.n278 VDD100 0.00224194
R13138 VDD100.n281 VDD100 0.00224194
R13139 VDD100 VDD100.n291 0.00224194
R13140 VDD100 VDD100.n288 0.00224194
R13141 VDD100 VDD100.n285 0.00224194
R13142 VDD100.n315 VDD100 0.00224194
R13143 VDD100.n318 VDD100 0.00224194
R13144 VDD100.n328 VDD100 0.00224194
R13145 VDD100 VDD100.n325 0.00224194
R13146 VDD100 VDD100.n322 0.00224194
R13147 VDD100.n465 VDD100 0.00224194
R13148 VDD100.n471 VDD100 0.00224194
R13149 VDD100.n474 VDD100 0.00224194
R13150 VDD100.n66 VDD100 0.00224194
R13151 VDD100.n69 VDD100 0.00224194
R13152 VDD100.n488 VDD100 0.00224194
R13153 VDD100.n494 VDD100 0.00224194
R13154 VDD100.n497 VDD100 0.00224194
R13155 VDD100 VDD100.n507 0.00224194
R13156 VDD100 VDD100.n504 0.00224194
R13157 VDD100.n333 VDD100 0.00219811
R13158 VDD100 VDD100.n443 0.00219811
R13159 VDD100.n169 VDD100 0.00166129
R13160 VDD100.n166 VDD100 0.00166129
R13161 VDD100 VDD100.n163 0.00166129
R13162 VDD100 VDD100.n160 0.00166129
R13163 VDD100 VDD100.n173 0.00166129
R13164 VDD100.n177 VDD100 0.00166129
R13165 VDD100 VDD100.n180 0.00166129
R13166 VDD100.n183 VDD100 0.00166129
R13167 VDD100.n206 VDD100 0.00166129
R13168 VDD100.n203 VDD100 0.00166129
R13169 VDD100 VDD100.n200 0.00166129
R13170 VDD100 VDD100.n197 0.00166129
R13171 VDD100.n211 VDD100 0.00166129
R13172 VDD100 VDD100.n214 0.00166129
R13173 VDD100 VDD100.n217 0.00166129
R13174 VDD100.n353 VDD100 0.00166129
R13175 VDD100.n378 VDD100 0.00166129
R13176 VDD100.n375 VDD100 0.00166129
R13177 VDD100 VDD100.n372 0.00166129
R13178 VDD100 VDD100.n369 0.00166129
R13179 VDD100.n383 VDD100 0.00166129
R13180 VDD100 VDD100.n386 0.00166129
R13181 VDD100 VDD100.n389 0.00166129
R13182 VDD100.n394 VDD100 0.00166129
R13183 VDD100.n419 VDD100 0.00166129
R13184 VDD100.n416 VDD100 0.00166129
R13185 VDD100 VDD100.n413 0.00166129
R13186 VDD100 VDD100.n410 0.00166129
R13187 VDD100.n424 VDD100 0.00166129
R13188 VDD100 VDD100.n427 0.00166129
R13189 VDD100.n431 VDD100 0.00166129
R13190 VDD100.n137 VDD100.n133 0.001625
R13191 VDD100 VDD100.n440 0.00115693
R13192 VDD100.n269 VDD100 0.00108064
R13193 VDD100 VDD100.n272 0.00108064
R13194 VDD100.n294 VDD100 0.00108064
R13195 VDD100.n306 VDD100 0.00108064
R13196 VDD100 VDD100.n309 0.00108064
R13197 VDD100.n462 VDD100 0.00108064
R13198 VDD100.n57 VDD100 0.00108064
R13199 VDD100 VDD100.n60 0.00108064
R13200 VDD100.n485 VDD100 0.00108064
R13201 VDD100 VDD100.n34 0.00108064
R13202 VDD100.n510 VDD100 0.00108064
R13203 VDD100.n234 VDD100 0.000828467
R13204 F0.n39 F0.t12 36.935
R13205 F0.n46 F0.t16 36.935
R13206 F0.n55 F0.t7 36.935
R13207 F0.n51 F0.t1 36.7829
R13208 F0.n10 F0.t2 31.528
R13209 F0.n1 F0.t13 31.528
R13210 F0.n25 F0.t9 31.528
R13211 F0.n17 F0.t24 31.528
R13212 F0.n4 F0.t3 25.7638
R13213 F0.n34 F0.t23 25.7638
R13214 F0.n15 F0.t4 25.7638
R13215 F0.n20 F0.t19 25.7638
R13216 F0.n62 F0.t21 25.432
R13217 F0.n39 F0.t10 18.1962
R13218 F0.n46 F0.t15 18.1962
R13219 F0.n55 F0.t5 18.1962
R13220 F0.n49 F0.t0 17.281
R13221 F0.n10 F0.t8 15.3826
R13222 F0.n1 F0.t20 15.3826
R13223 F0.n25 F0.t17 15.3826
R13224 F0.n17 F0.t11 15.3826
R13225 F0.n4 F0.t18 13.2969
R13226 F0.n34 F0.t14 13.2969
R13227 F0.n15 F0.t6 13.2969
R13228 F0.n20 F0.t22 13.2969
R13229 F0.n61 F0.t25 12.4441
R13230 F0 F0.n69 11.7386
R13231 F0.n69 F0.n37 11.5868
R13232 F0.n39 F0 8.01615
R13233 F0.n51 F0 8.01336
R13234 F0.n46 F0 8.01224
R13235 F0.n18 F0.n17 7.6291
R13236 F0.n2 F0.n1 7.6289
R13237 F0.n12 F0.n10 7.62076
R13238 F0.n26 F0.n25 7.62076
R13239 F0 F0.n9 4.53443
R13240 F0.n24 F0 4.53443
R13241 F0.n13 F0 4.52853
R13242 F0.n6 F0 4.52833
R13243 F0.n36 F0 4.52833
R13244 F0.n30 F0 4.52833
R13245 F0.n22 F0 4.52833
R13246 F0.n57 F0 4.52643
R13247 F0.n63 F0.n62 4.5005
R13248 F0.n52 F0.n51 4.5005
R13249 F0.n50 F0.n49 3.62236
R13250 F0.n56 F0.n55 2.8805
R13251 F0.n40 F0.n39 2.8798
R13252 F0.n47 F0.n46 2.8789
R13253 F0 F0.n0 2.26791
R13254 F0.n35 F0.n33 2.25478
R13255 F0.n32 F0.n16 2.25386
R13256 F0.n31 F0.n16 2.2505
R13257 F0.n35 F0.n14 2.2505
R13258 F0.n65 F0.n64 2.2485
R13259 F0.n61 F0 2.20644
R13260 F0.n8 F0.n7 2.19776
R13261 F0.n28 F0.n23 2.19633
R13262 F0.n5 F0.n4 2.11815
R13263 F0.n35 F0.n34 2.11815
R13264 F0.n16 F0.n15 2.11815
R13265 F0.n21 F0.n20 2.11815
R13266 F0.n33 F0.n32 1.87738
R13267 F0.n58 F0.n57 1.79371
R13268 F0.n60 F0.n59 1.60479
R13269 F0.n59 F0.n58 1.59764
R13270 F0.n12 F0.n11 1.5005
R13271 F0.n27 F0.n26 1.5005
R13272 F0.n44 F0.n43 1.49986
R13273 F0.n30 F0.n29 1.31185
R13274 F0.n23 F0.n22 1.2853
R13275 F0.n7 F0.n6 1.28387
R13276 F0.n59 F0.n48 1.27535
R13277 F0.n58 F0.n53 1.2731
R13278 F0.n37 F0.n36 1.27101
R13279 F0.n67 F0.n60 1.20307
R13280 F0.n5 F0.n3 1.13046
R13281 F0.n21 F0.n19 1.13
R13282 F0.n57 F0.n54 1.12143
R13283 F0.n7 F0.n2 0.948428
R13284 F0.n23 F0.n18 0.948389
R13285 F0.n62 F0.n61 0.802693
R13286 F0.n69 F0.n68 0.5369
R13287 F0.n60 F0.n45 0.128961
R13288 F0.n18 F0 0.109321
R13289 F0.n2 F0 0.108522
R13290 F0 F0.n65 0.0902065
R13291 F0.n54 F0 0.0822111
R13292 F0.n9 F0 0.0780742
R13293 F0.n24 F0 0.0780197
R13294 F0.n66 F0 0.0612636
R13295 F0.n53 F0 0.0537005
R13296 F0.n48 F0 0.0533296
R13297 F0.n43 F0 0.0532041
R13298 F0.n37 F0.n13 0.0399145
R13299 F0.n12 F0.n9 0.0373852
R13300 F0.n26 F0.n24 0.0373852
R13301 F0.n13 F0.n8 0.0359098
R13302 F0.n29 F0.n28 0.0359098
R13303 F0.n65 F0.n38 0.0314769
R13304 F0.n22 F0.n19 0.0303837
R13305 F0.n6 F0.n3 0.0303834
R13306 F0.n31 F0.n30 0.0289694
R13307 F0.n36 F0.n14 0.0289694
R13308 F0.n45 F0.n44 0.0273966
R13309 F0.n48 F0.n47 0.021401
R13310 F0.n53 F0.n52 0.0173852
R13311 F0.n47 F0 0.017274
R13312 F0.n33 F0 0.0169815
R13313 F0.n32 F0 0.0160631
R13314 F0.n40 F0 0.0147725
R13315 F0.n67 F0.n66 0.0131
R13316 F0 F0.n56 0.0127034
R13317 F0.n42 F0.n41 0.0122391
R13318 F0.n56 F0.n54 0.0116287
R13319 F0.n64 F0.n63 0.0112609
R13320 F0 F0.n50 0.0107857
R13321 F0 F0.n12 0.00935246
R13322 F0.n43 F0.n42 0.00925458
R13323 F0.n52 F0.n50 0.00821429
R13324 F0.n63 F0 0.00734783
R13325 F0.n68 F0.n38 0.00692857
R13326 F0.n11 F0 0.00345082
R13327 F0.n27 F0 0.00345082
R13328 F0.n41 F0.n40 0.00287748
R13329 F0 F0.n31 0.00233673
R13330 F0 F0.n14 0.00233673
R13331 F0.n11 F0.n8 0.00197541
R13332 F0.n28 F0.n27 0.00197541
R13333 F0.n3 F0 0.00192201
R13334 F0.n19 F0 0.00192164
R13335 F0 F0.n5 0.00142783
R13336 F0 F0.n35 0.00142783
R13337 F0 F0.n16 0.00142783
R13338 F0 F0.n21 0.00142783
R13339 F0.n68 F0.n67 0.0014
R13340 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n19 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t11 36.935
R13341 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n18 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t10 36.935
R13342 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n22 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t15 36.935
R13343 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n21 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t18 36.935
R13344 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n13 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t5 36.935
R13345 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n15 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t20 31.4332
R13346 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n24 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t8 30.6613
R13347 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n20 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t17 25.4744
R13348 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n26 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t9 25.4744
R13349 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n24 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t12 21.6718
R13350 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n19 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t6 18.1962
R13351 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n18 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t7 18.1962
R13352 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n22 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t13 18.1962
R13353 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n21 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t16 18.1962
R13354 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n13 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t4 18.1962
R13355 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n15 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t19 15.3826
R13356 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n26 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t14 14.1417
R13357 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n20 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t3 14.1417
R13358 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n0 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n25 9.9005
R13359 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n12 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t0 7.09905
R13360 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n16 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n15 6.86029
R13361 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n17 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n14 5.01077
R13362 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n2 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n3 1.11863
R13363 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n4 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n5 1.11863
R13364 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n20 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n9 1.42995
R13365 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n0 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n1 1.11781
R13366 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n12 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n11 3.25053
R13367 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n11 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t2 2.2755
R13368 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n11 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n10 2.2755
R13369 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n28 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n27 2.2505
R13370 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n23 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n9 1.16587
R13371 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n14 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n13 2.13459
R13372 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n3 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n19 2.13265
R13373 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n5 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n22 2.13265
R13374 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n2 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n7 2.63776
R13375 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n4 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n8 2.63776
R13376 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n27 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n17 1.52773
R13377 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n18 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n7 2.13261
R13378 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n21 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n8 2.13281
R13379 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n1 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n26 1.42999
R13380 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n6 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n24 1.41101
R13381 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n17 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n16 1.12067
R13382 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n25 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n23 0.286289
R13383 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n1 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 0.196008
R13384 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n9 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 0.196051
R13385 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n28 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n12 0.0905
R13386 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n16 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 0.0857632
R13387 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n28 0.0834687
R13388 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n6 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 0.104828
R13389 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n14 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 0.0800273
R13390 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n8 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 0.0771461
R13391 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n7 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 0.0771461
R13392 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n5 0.077103
R13393 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n3 0.077103
R13394 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n27 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 0.0289903
R13395 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n25 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n6 7.13895
R13396 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n0 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n2 1.18681
R13397 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n23 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n4 0.938524
R13398 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n0 0.680217
R13399 VDD110.t16 VDD110.n374 57397.6
R13400 VDD110.t10 VDD110.n413 57397.6
R13401 VDD110.t22 VDD110.n232 57397.6
R13402 VDD110.n18 VDD110.t62 2529.02
R13403 VDD110.n24 VDD110 2301.38
R13404 VDD110.n525 VDD110 2301.38
R13405 VDD110.n25 VDD110.n24 1842.37
R13406 VDD110.n526 VDD110.n525 1842.37
R13407 VDD110.n28 VDD110.t329 1403.56
R13408 VDD110.n30 VDD110.t31 1242.86
R13409 VDD110.n263 VDD110.t302 1105.93
R13410 VDD110.n21 VDD110.t171 1105.93
R13411 VDD110.t89 VDD110.n15 1011.51
R13412 VDD110.t127 VDD110.t344 961.905
R13413 VDD110.t360 VDD110.t225 961.905
R13414 VDD110.t38 VDD110.t265 961.905
R13415 VDD110.t142 VDD110.t182 961.905
R13416 VDD110.t81 VDD110.t5 961.905
R13417 VDD110.t205 VDD110.t33 961.905
R13418 VDD110.n374 VDD110.t259 864.287
R13419 VDD110.n413 VDD110.t380 864.287
R13420 VDD110.n232 VDD110.t337 864.287
R13421 VDD110.t168 VDD110.n1 857.144
R13422 VDD110.t454 VDD110.n5 857.144
R13423 VDD110.n24 VDD110.t116 812.681
R13424 VDD110.n525 VDD110.t96 812.681
R13425 VDD110.t299 VDD110.t415 765.152
R13426 VDD110.t276 VDD110.t269 765.152
R13427 VDD110.t439 VDD110.t284 765.152
R13428 VDD110.t256 VDD110.t68 765.152
R13429 VDD110.t135 VDD110.t66 765.152
R13430 VDD110.t178 VDD110.t180 765.152
R13431 VDD110.t227 VDD110.t78 765.152
R13432 VDD110.t339 VDD110.t425 765.152
R13433 VDD110.t7 VDD110.t200 765.152
R13434 VDD110.t35 VDD110.t104 765.152
R13435 VDD110.t385 VDD110.t382 765.152
R13436 VDD110.t161 VDD110.t106 765.152
R13437 VDD110.t133 VDD110.t130 765.152
R13438 VDD110.t261 VDD110.t108 765.152
R13439 VDD110.t58 VDD110.t346 765.152
R13440 VDD110.t376 VDD110.t373 765.152
R13441 VDD110.t0 VDD110.t366 765.152
R13442 VDD110.t114 VDD110.t191 765.152
R13443 VDD110.t370 VDD110.t193 765.152
R13444 VDD110.t368 VDD110.t3 765.152
R13445 VDD110.t417 VDD110.t102 765.152
R13446 VDD110.t253 VDD110.t443 765.152
R13447 VDD110.t64 VDD110.t138 765.152
R13448 VDD110.t87 VDD110.t98 765.152
R13449 VDD110.t60 VDD110.t306 765.152
R13450 VDD110.t286 VDD110.t125 765.152
R13451 VDD110.t413 VDD110.t455 765.152
R13452 VDD110.t166 VDD110.t236 765.152
R13453 VDD110.t449 VDD110.t316 765.152
R13454 VDD110.t378 VDD110.t335 765.152
R13455 VDD110.t233 VDD110.t121 765.152
R13456 VDD110.t314 VDD110.t452 765.152
R13457 VDD110.t318 VDD110.t282 765.152
R13458 VDD110.t309 VDD110.t312 765.152
R13459 VDD110.t123 VDD110.t289 765.152
R13460 VDD110.t48 VDD110.t231 765.152
R13461 VDD110.t296 VDD110.t29 765.152
R13462 VDD110.t274 VDD110.t272 765.152
R13463 VDD110.t429 VDD110.t119 765.152
R13464 VDD110.n260 VDD110.t304 747.159
R13465 VDD110.t251 VDD110.t229 642.843
R13466 VDD110.n22 VDD110.t169 581.375
R13467 VDD110 VDD110.n22 572.967
R13468 VDD110.n493 VDD110.t364 480.199
R13469 VDD110.t329 VDD110.t475 461.096
R13470 VDD110.t329 VDD110.t291 461.096
R13471 VDD110.t293 VDD110.t43 461.096
R13472 VDD110.t93 VDD110.t41 461.096
R13473 VDD110 VDD110.n163 429.187
R13474 VDD110 VDD110.n131 429.187
R13475 VDD110 VDD110.n148 429.187
R13476 VDD110 VDD110.n477 426.699
R13477 VDD110 VDD110.n450 426.699
R13478 VDD110 VDD110.n403 426.699
R13479 VDD110 VDD110.n363 426.699
R13480 VDD110.n275 VDD110 424.618
R13481 VDD110 VDD110.n269 424.618
R13482 VDD110 VDD110.n264 422.557
R13483 VDD110.n486 VDD110.n485 421.611
R13484 VDD110.n15 VDD110.t247 420.793
R13485 VDD110.n163 VDD110.t447 386.365
R13486 VDD110.n194 VDD110.t239 386.365
R13487 VDD110.n477 VDD110.t19 386.365
R13488 VDD110.n450 VDD110.t189 386.365
R13489 VDD110.n403 VDD110.t25 386.365
R13490 VDD110.n363 VDD110.t112 386.365
R13491 VDD110.n275 VDD110.t362 386.365
R13492 VDD110.n269 VDD110.t218 386.365
R13493 VDD110.n148 VDD110.t243 386.365
R13494 VDD110.n131 VDD110.t278 386.365
R13495 VDD110.t110 VDD110.t410 380.952
R13496 VDD110.t155 VDD110.t360 380.952
R13497 VDD110.t387 VDD110.t395 380.952
R13498 VDD110.t212 VDD110.t142 380.952
R13499 VDD110.t423 VDD110.t398 380.952
R13500 VDD110.t73 VDD110.t205 380.952
R13501 VDD110.t354 VDD110.n275 378.788
R13502 VDD110.n269 VDD110.t147 378.788
R13503 VDD110.n264 VDD110.t357 378.788
R13504 VDD110.t53 VDD110.n198 375
R13505 VDD110.n195 VDD110.n194 368.159
R13506 VDD110.n24 VDD110.t293 351.586
R13507 VDD110.n525 VDD110.t93 351.586
R13508 VDD110.n198 VDD110.n196 343.137
R13509 VDD110.t163 VDD110.n486 306.118
R13510 VDD110.t484 VDD110.t439 303.031
R13511 VDD110.t472 VDD110.t178 303.031
R13512 VDD110.t200 VDD110.t70 303.031
R13513 VDD110.t202 VDD110.t161 303.031
R13514 VDD110.t346 VDD110.t144 303.031
R13515 VDD110.t191 VDD110.t215 303.031
R13516 VDD110.t404 VDD110.t368 303.031
R13517 VDD110.t220 VDD110.t417 303.031
R13518 VDD110.t401 VDD110.t64 303.031
R13519 VDD110.t460 VDD110.t87 303.031
R13520 VDD110.t455 VDD110.t463 303.031
R13521 VDD110.t335 VDD110.t479 303.031
R13522 VDD110.t392 VDD110.t314 303.031
R13523 VDD110.t466 VDD110.t318 303.031
R13524 VDD110.t389 VDD110.t123 303.031
R13525 VDD110.t491 VDD110.t48 303.031
R13526 VDD110.t407 VDD110.t274 303.031
R13527 VDD110.t469 VDD110.t429 303.031
R13528 VDD110.n489 VDD110.n201 298.536
R13529 VDD110.n493 VDD110.n201 288
R13530 VDD110.n366 VDD110.t351 242.857
R13531 VDD110.n368 VDD110.t127 242.857
R13532 VDD110.t410 VDD110.n371 242.857
R13533 VDD110.n375 VDD110.t155 242.857
R13534 VDD110.n405 VDD110.t150 242.857
R13535 VDD110.n407 VDD110.t38 242.857
R13536 VDD110.t395 VDD110.n410 242.857
R13537 VDD110.n414 VDD110.t212 242.857
R13538 VDD110.n224 VDD110.t209 242.857
R13539 VDD110.n226 VDD110.t81 242.857
R13540 VDD110.t398 VDD110.n229 242.857
R13541 VDD110.n233 VDD110.t73 242.857
R13542 VDD110.n3 VDD110.n2 199.562
R13543 VDD110.n7 VDD110.n6 199.562
R13544 VDD110.n154 VDD110.t436 193.183
R13545 VDD110.n155 VDD110.t299 193.183
R13546 VDD110.n161 VDD110.t269 193.183
R13547 VDD110.n162 VDD110.t484 193.183
R13548 VDD110.n186 VDD110.t173 193.183
R13549 VDD110.n188 VDD110.t256 193.183
R13550 VDD110.n190 VDD110.t135 193.183
R13551 VDD110.n193 VDD110.t472 193.183
R13552 VDD110.n199 VDD110.t53 193.183
R13553 VDD110.n459 VDD110.t197 193.183
R13554 VDD110.n465 VDD110.t78 193.183
R13555 VDD110.n466 VDD110.t339 193.183
R13556 VDD110.n476 VDD110.t70 193.183
R13557 VDD110.n437 VDD110.t158 193.183
R13558 VDD110.n438 VDD110.t35 193.183
R13559 VDD110.n448 VDD110.t382 193.183
R13560 VDD110.n449 VDD110.t202 193.183
R13561 VDD110.n389 VDD110.t348 193.183
R13562 VDD110.n395 VDD110.t130 193.183
R13563 VDD110.n396 VDD110.t261 193.183
R13564 VDD110.n402 VDD110.t144 193.183
R13565 VDD110.n350 VDD110.t186 193.183
R13566 VDD110.n356 VDD110.t373 193.183
R13567 VDD110.n357 VDD110.t0 193.183
R13568 VDD110.n362 VDD110.t215 193.183
R13569 VDD110.n295 VDD110.t420 193.183
R13570 VDD110.n297 VDD110.t370 193.183
R13571 VDD110.n300 VDD110.t404 193.183
R13572 VDD110.n303 VDD110.t220 193.183
R13573 VDD110.n276 VDD110.t354 193.183
R13574 VDD110.n274 VDD110.t147 193.183
R13575 VDD110.n268 VDD110.t357 193.183
R13576 VDD110.n165 VDD110.t90 193.183
R13577 VDD110.n167 VDD110.t253 193.183
R13578 VDD110.n170 VDD110.t401 193.183
R13579 VDD110.n173 VDD110.t460 193.183
R13580 VDD110.n135 VDD110.t457 193.183
R13581 VDD110.n141 VDD110.t306 193.183
R13582 VDD110.n142 VDD110.t286 193.183
R13583 VDD110.n147 VDD110.t463 193.183
R13584 VDD110.n118 VDD110.t332 193.183
R13585 VDD110.n124 VDD110.t236 193.183
R13586 VDD110.n125 VDD110.t449 193.183
R13587 VDD110.n130 VDD110.t479 193.183
R13588 VDD110.n97 VDD110.t326 193.183
R13589 VDD110.n99 VDD110.t233 193.183
R13590 VDD110.n102 VDD110.t392 193.183
R13591 VDD110.n105 VDD110.t466 193.183
R13592 VDD110.n69 VDD110.t50 193.183
R13593 VDD110.n71 VDD110.t309 193.183
R13594 VDD110.n74 VDD110.t389 193.183
R13595 VDD110.n77 VDD110.t491 193.183
R13596 VDD110.n41 VDD110.t431 193.183
R13597 VDD110.n43 VDD110.t296 193.183
R13598 VDD110.n46 VDD110.t407 193.183
R13599 VDD110.n49 VDD110.t469 193.183
R13600 VDD110.n488 VDD110.t434 191.288
R13601 VDD110.t264 VDD110.t419 175.631
R13602 VDD110.t118 VDD110.t89 175.631
R13603 VDD110.n2 VDD110.t168 170.577
R13604 VDD110.n2 VDD110.t324 170.577
R13605 VDD110.n6 VDD110.t454 170.577
R13606 VDD110.n6 VDD110.t176 170.577
R13607 VDD110.t304 VDD110.n259 153.678
R13608 VDD110.t62 VDD110.n17 153.678
R13609 VDD110.t434 VDD110.t84 151.516
R13610 VDD110.t344 VDD110.n366 138.095
R13611 VDD110.t259 VDD110.n368 138.095
R13612 VDD110.t225 VDD110.n371 138.095
R13613 VDD110.n375 VDD110.t16 138.095
R13614 VDD110.t265 VDD110.n405 138.095
R13615 VDD110.t380 VDD110.n407 138.095
R13616 VDD110.t182 VDD110.n410 138.095
R13617 VDD110.n414 VDD110.t10 138.095
R13618 VDD110.t5 VDD110.n224 138.095
R13619 VDD110.t337 VDD110.n226 138.095
R13620 VDD110.t33 VDD110.n229 138.095
R13621 VDD110.n233 VDD110.t22 138.095
R13622 VDD110.n198 VDD110.t56 132.353
R13623 VDD110.n209 VDD110.t195 124.511
R13624 VDD110.n489 VDD110.n488 117.216
R13625 VDD110.n196 VDD110.n195 112.746
R13626 VDD110.t415 VDD110.n154 109.849
R13627 VDD110.n155 VDD110.t276 109.849
R13628 VDD110.t284 VDD110.n161 109.849
R13629 VDD110.t447 VDD110.n162 109.849
R13630 VDD110.t68 VDD110.n186 109.849
R13631 VDD110.t66 VDD110.n188 109.849
R13632 VDD110.t180 VDD110.n190 109.849
R13633 VDD110.t239 VDD110.n193 109.849
R13634 VDD110.n199 VDD110.t320 109.849
R13635 VDD110.n459 VDD110.t227 109.849
R13636 VDD110.t425 VDD110.n465 109.849
R13637 VDD110.n466 VDD110.t7 109.849
R13638 VDD110.t19 VDD110.n476 109.849
R13639 VDD110.t104 VDD110.n437 109.849
R13640 VDD110.n438 VDD110.t385 109.849
R13641 VDD110.t106 VDD110.n448 109.849
R13642 VDD110.t189 VDD110.n449 109.849
R13643 VDD110.n389 VDD110.t133 109.849
R13644 VDD110.t108 VDD110.n395 109.849
R13645 VDD110.n396 VDD110.t58 109.849
R13646 VDD110.t25 VDD110.n402 109.849
R13647 VDD110.n350 VDD110.t376 109.849
R13648 VDD110.t366 VDD110.n356 109.849
R13649 VDD110.n357 VDD110.t114 109.849
R13650 VDD110.t112 VDD110.n362 109.849
R13651 VDD110.t193 VDD110.n295 109.849
R13652 VDD110.t3 VDD110.n297 109.849
R13653 VDD110.t102 VDD110.n300 109.849
R13654 VDD110.n303 VDD110.t13 109.849
R13655 VDD110.n276 VDD110.t153 109.849
R13656 VDD110.t362 VDD110.n274 109.849
R13657 VDD110.t218 VDD110.n268 109.849
R13658 VDD110.t443 VDD110.n165 109.849
R13659 VDD110.t138 VDD110.n167 109.849
R13660 VDD110.t98 VDD110.n170 109.849
R13661 VDD110.n173 VDD110.t241 109.849
R13662 VDD110.n135 VDD110.t60 109.849
R13663 VDD110.t125 VDD110.n141 109.849
R13664 VDD110.n142 VDD110.t413 109.849
R13665 VDD110.t243 VDD110.n147 109.849
R13666 VDD110.n118 VDD110.t166 109.849
R13667 VDD110.t316 VDD110.n124 109.849
R13668 VDD110.n125 VDD110.t378 109.849
R13669 VDD110.t278 VDD110.n130 109.849
R13670 VDD110.t121 VDD110.n97 109.849
R13671 VDD110.t452 VDD110.n99 109.849
R13672 VDD110.t282 VDD110.n102 109.849
R13673 VDD110.n105 VDD110.t280 109.849
R13674 VDD110.t312 VDD110.n69 109.849
R13675 VDD110.t289 VDD110.n71 109.849
R13676 VDD110.t231 VDD110.n74 109.849
R13677 VDD110.n77 VDD110.t245 109.849
R13678 VDD110.t29 VDD110.n41 109.849
R13679 VDD110.t272 VDD110.n43 109.849
R13680 VDD110.t119 VDD110.n46 109.849
R13681 VDD110.n49 VDD110.t445 109.849
R13682 VDD110.n374 VDD110.t110 97.6195
R13683 VDD110.n413 VDD110.t387 97.6195
R13684 VDD110.n232 VDD110.t423 97.6195
R13685 VDD110.t84 VDD110.n208 96.5914
R13686 VDD110.n487 VDD110.n209 90.2261
R13687 VDD110.n22 VDD110.t249 80.0005
R13688 VDD110.n487 VDD110.t163 76.2337
R13689 VDD110.t31 VDD110 68.2053
R13690 VDD110.n15 VDD110 65.7064
R13691 VDD110.n477 VDD110.t76 62.1896
R13692 VDD110.n450 VDD110.t223 62.1896
R13693 VDD110.n403 VDD110.t140 62.1896
R13694 VDD110.n363 VDD110.t207 62.1896
R13695 VDD110.n30 VDD110.t427 61.9053
R13696 VDD110.n275 VDD110.t267 61.8817
R13697 VDD110.n269 VDD110.t100 61.8817
R13698 VDD110.n264 VDD110.t251 61.5769
R13699 VDD110 VDD110.n195 61.0269
R13700 VDD110.n163 VDD110.t482 59.702
R13701 VDD110.n194 VDD110.t489 59.702
R13702 VDD110.n148 VDD110.t487 59.702
R13703 VDD110.n131 VDD110.t477 59.702
R13704 VDD110.n486 VDD110.t164 59.4064
R13705 VDD110.n260 VDD110.t302 55.0852
R13706 VDD110.t229 VDD110.n263 55.0852
R13707 VDD110.n18 VDD110.t171 55.0852
R13708 VDD110.t169 VDD110.n21 55.0852
R13709 VDD110.n208 VDD110.t45 54.9247
R13710 VDD110.n333 VDD110.t12 30.9379
R13711 VDD110.n305 VDD110.t9 30.9379
R13712 VDD110.n324 VDD110.t24 30.7203
R13713 VDD110.n311 VDD110.t18 30.7203
R13714 VDD110.n329 VDD110.t15 30.2877
R13715 VDD110.n317 VDD110.t21 29.1661
R13716 VDD110.n329 VDD110.t497 24.9141
R13717 VDD110.n333 VDD110.t498 24.5101
R13718 VDD110.n319 VDD110.t495 24.5101
R13719 VDD110.n305 VDD110.t499 24.5101
R13720 VDD110.n311 VDD110.t496 24.4814
R13721 VDD110.n324 VDD110.t494 24.4814
R13722 VDD110.n259 VDD110.t264 21.9544
R13723 VDD110.n17 VDD110.t118 21.9544
R13724 VDD110.n488 VDD110.n487 20.147
R13725 VDD110 VDD110.n537 14.2941
R13726 VDD110.n13 VDD110.t170 14.0055
R13727 VDD110.n16 VDD110.t63 13.2223
R13728 VDD110.n261 VDD110.t303 12.3869
R13729 VDD110.n19 VDD110.t172 12.3869
R13730 VDD110.n8 VDD110.t32 12.3869
R13731 VDD110.n13 VDD110.t250 10.1341
R13732 VDD110.n491 VDD110.n490 9.64171
R13733 VDD110.n319 VDD110.n318 8.0005
R13734 VDD110.n317 VDD110.n316 8.0005
R13735 VDD110.n485 VDD110.n484 7.01458
R13736 VDD110.n492 VDD110.n491 6.69176
R13737 VDD110.n334 VDD110.n332 6.39748
R13738 VDD110.n259 VDD110 6.30126
R13739 VDD110.n534 VDD110.n533 6.3005
R13740 VDD110.n533 VDD110.n529 6.3005
R13741 VDD110 VDD110.n493 6.3005
R13742 VDD110.n495 VDD110.n201 6.3005
R13743 VDD110 VDD110.n489 6.3005
R13744 VDD110.n347 VDD110.n295 6.3005
R13745 VDD110.n344 VDD110.n297 6.3005
R13746 VDD110.n341 VDD110.n300 6.3005
R13747 VDD110.n338 VDD110.n303 6.3005
R13748 VDD110.n351 VDD110.n350 6.3005
R13749 VDD110.n356 VDD110.n355 6.3005
R13750 VDD110.n358 VDD110.n357 6.3005
R13751 VDD110.n362 VDD110.n361 6.3005
R13752 VDD110.n385 VDD110.n366 6.3005
R13753 VDD110.n382 VDD110.n368 6.3005
R13754 VDD110.n379 VDD110.n371 6.3005
R13755 VDD110.n376 VDD110.n375 6.3005
R13756 VDD110.n390 VDD110.n389 6.3005
R13757 VDD110.n395 VDD110.n394 6.3005
R13758 VDD110.n397 VDD110.n396 6.3005
R13759 VDD110 VDD110.n260 6.3005
R13760 VDD110.n263 VDD110.n262 6.3005
R13761 VDD110.n268 VDD110.n267 6.3005
R13762 VDD110.n274 VDD110.n273 6.3005
R13763 VDD110.n277 VDD110.n276 6.3005
R13764 VDD110.n402 VDD110.n401 6.3005
R13765 VDD110.n424 VDD110.n405 6.3005
R13766 VDD110.n421 VDD110.n407 6.3005
R13767 VDD110.n418 VDD110.n410 6.3005
R13768 VDD110.n415 VDD110.n414 6.3005
R13769 VDD110.n437 VDD110.n436 6.3005
R13770 VDD110.n439 VDD110.n438 6.3005
R13771 VDD110.n448 VDD110.n447 6.3005
R13772 VDD110.n449 VDD110.n246 6.3005
R13773 VDD110.n243 VDD110.n224 6.3005
R13774 VDD110.n240 VDD110.n226 6.3005
R13775 VDD110.n237 VDD110.n229 6.3005
R13776 VDD110.n234 VDD110.n233 6.3005
R13777 VDD110.n460 VDD110.n459 6.3005
R13778 VDD110.n465 VDD110.n464 6.3005
R13779 VDD110.n467 VDD110.n466 6.3005
R13780 VDD110.n476 VDD110.n475 6.3005
R13781 VDD110.n498 VDD110.n199 6.3005
R13782 VDD110 VDD110.n196 6.3005
R13783 VDD110.n174 VDD110.n173 6.3005
R13784 VDD110.n177 VDD110.n170 6.3005
R13785 VDD110.n180 VDD110.n167 6.3005
R13786 VDD110.n183 VDD110.n165 6.3005
R13787 VDD110.n512 VDD110.n186 6.3005
R13788 VDD110.n509 VDD110.n188 6.3005
R13789 VDD110.n506 VDD110.n190 6.3005
R13790 VDD110.n503 VDD110.n193 6.3005
R13791 VDD110.n106 VDD110.n105 6.3005
R13792 VDD110.n109 VDD110.n102 6.3005
R13793 VDD110.n112 VDD110.n99 6.3005
R13794 VDD110.n115 VDD110.n97 6.3005
R13795 VDD110.n119 VDD110.n118 6.3005
R13796 VDD110.n124 VDD110.n123 6.3005
R13797 VDD110.n126 VDD110.n125 6.3005
R13798 VDD110.n130 VDD110.n129 6.3005
R13799 VDD110.n78 VDD110.n77 6.3005
R13800 VDD110.n81 VDD110.n74 6.3005
R13801 VDD110.n84 VDD110.n71 6.3005
R13802 VDD110.n87 VDD110.n69 6.3005
R13803 VDD110.n136 VDD110.n135 6.3005
R13804 VDD110.n141 VDD110.n140 6.3005
R13805 VDD110.n143 VDD110.n142 6.3005
R13806 VDD110.n147 VDD110.n146 6.3005
R13807 VDD110.n50 VDD110.n49 6.3005
R13808 VDD110.n53 VDD110.n46 6.3005
R13809 VDD110.n56 VDD110.n43 6.3005
R13810 VDD110.n59 VDD110.n41 6.3005
R13811 VDD110.n154 VDD110.n153 6.3005
R13812 VDD110.n156 VDD110.n155 6.3005
R13813 VDD110.n161 VDD110.n160 6.3005
R13814 VDD110.n517 VDD110.n162 6.3005
R13815 VDD110.n17 VDD110.n16 6.3005
R13816 VDD110.n21 VDD110.n20 6.3005
R13817 VDD110 VDD110.n18 6.3005
R13818 VDD110.n31 VDD110.n30 6.3005
R13819 VDD110.n1 VDD110 6.3005
R13820 VDD110.n5 VDD110 6.3005
R13821 VDD110.n23 VDD110.t117 5.85907
R13822 VDD110.n519 VDD110.n518 5.69603
R13823 VDD110.n322 VDD110.n321 5.30733
R13824 VDD110.n376 VDD110.t17 5.213
R13825 VDD110.n415 VDD110.t11 5.213
R13826 VDD110.n234 VDD110.t23 5.213
R13827 VDD110.n174 VDD110.t242 5.213
R13828 VDD110.n106 VDD110.t281 5.213
R13829 VDD110.n78 VDD110.t246 5.213
R13830 VDD110.n50 VDD110.t446 5.213
R13831 VDD110.n398 VDD110.t59 5.16792
R13832 VDD110.n497 VDD110.t321 5.15377
R13833 VDD110.n499 VDD110.n197 5.13287
R13834 VDD110.n205 VDD110.n204 5.13287
R13835 VDD110.n206 VDD110.t47 5.13287
R13836 VDD110.n206 VDD110.t46 5.13287
R13837 VDD110.n348 VDD110.n294 5.13287
R13838 VDD110.n346 VDD110.t194 5.13287
R13839 VDD110.n345 VDD110.n296 5.13287
R13840 VDD110.n343 VDD110.t4 5.13287
R13841 VDD110.n340 VDD110.t103 5.13287
R13842 VDD110.n349 VDD110.n293 5.13287
R13843 VDD110.n352 VDD110.t377 5.13287
R13844 VDD110.n353 VDD110.n292 5.13287
R13845 VDD110.n354 VDD110.t367 5.13287
R13846 VDD110.n291 VDD110.n290 5.13287
R13847 VDD110.n359 VDD110.t115 5.13287
R13848 VDD110.n287 VDD110.t113 5.13287
R13849 VDD110.n386 VDD110.n365 5.13287
R13850 VDD110.n384 VDD110.t345 5.13287
R13851 VDD110.n383 VDD110.n367 5.13287
R13852 VDD110.n381 VDD110.t260 5.13287
R13853 VDD110.n378 VDD110.t226 5.13287
R13854 VDD110.n388 VDD110.n286 5.13287
R13855 VDD110.n391 VDD110.t134 5.13287
R13856 VDD110.n392 VDD110.n285 5.13287
R13857 VDD110.n393 VDD110.t109 5.13287
R13858 VDD110.n284 VDD110.n283 5.13287
R13859 VDD110.n280 VDD110.t26 5.13287
R13860 VDD110.n266 VDD110.n256 5.13287
R13861 VDD110.n255 VDD110.t219 5.13287
R13862 VDD110.n271 VDD110.n254 5.13287
R13863 VDD110.n272 VDD110.t363 5.13287
R13864 VDD110.n252 VDD110.n251 5.13287
R13865 VDD110.n278 VDD110.t154 5.13287
R13866 VDD110.n425 VDD110.n404 5.13287
R13867 VDD110.n423 VDD110.t266 5.13287
R13868 VDD110.n422 VDD110.n406 5.13287
R13869 VDD110.n420 VDD110.t381 5.13287
R13870 VDD110.n417 VDD110.t183 5.13287
R13871 VDD110.n250 VDD110.n249 5.13287
R13872 VDD110.n435 VDD110.t105 5.13287
R13873 VDD110.n434 VDD110.n433 5.13287
R13874 VDD110.n440 VDD110.t386 5.13287
R13875 VDD110.n441 VDD110.n247 5.13287
R13876 VDD110.n445 VDD110.t107 5.13287
R13877 VDD110.n452 VDD110.t190 5.13287
R13878 VDD110.n244 VDD110.n223 5.13287
R13879 VDD110.n242 VDD110.t6 5.13287
R13880 VDD110.n241 VDD110.n225 5.13287
R13881 VDD110.n239 VDD110.t338 5.13287
R13882 VDD110.n236 VDD110.t34 5.13287
R13883 VDD110.n458 VDD110.n222 5.13287
R13884 VDD110.n461 VDD110.t228 5.13287
R13885 VDD110.n463 VDD110.n221 5.13287
R13886 VDD110.n219 VDD110.t426 5.13287
R13887 VDD110.n468 VDD110.n220 5.13287
R13888 VDD110.n217 VDD110.t8 5.13287
R13889 VDD110.n214 VDD110.t20 5.13287
R13890 VDD110.n502 VDD110.t240 5.13287
R13891 VDD110.n505 VDD110.t181 5.13287
R13892 VDD110.n507 VDD110.n189 5.13287
R13893 VDD110.n508 VDD110.t67 5.13287
R13894 VDD110.n510 VDD110.n187 5.13287
R13895 VDD110.n511 VDD110.t69 5.13287
R13896 VDD110.n513 VDD110.n185 5.13287
R13897 VDD110.n176 VDD110.t99 5.13287
R13898 VDD110.n179 VDD110.t139 5.13287
R13899 VDD110.n181 VDD110.n166 5.13287
R13900 VDD110.n182 VDD110.t444 5.13287
R13901 VDD110.n184 VDD110.n164 5.13287
R13902 VDD110.n89 VDD110.t279 5.13287
R13903 VDD110.n127 VDD110.t379 5.13287
R13904 VDD110.n93 VDD110.n92 5.13287
R13905 VDD110.n122 VDD110.t317 5.13287
R13906 VDD110.n121 VDD110.n94 5.13287
R13907 VDD110.n120 VDD110.t167 5.13287
R13908 VDD110.n117 VDD110.n95 5.13287
R13909 VDD110.n108 VDD110.t283 5.13287
R13910 VDD110.n111 VDD110.t453 5.13287
R13911 VDD110.n113 VDD110.n98 5.13287
R13912 VDD110.n114 VDD110.t122 5.13287
R13913 VDD110.n116 VDD110.n96 5.13287
R13914 VDD110.n80 VDD110.t232 5.13287
R13915 VDD110.n83 VDD110.t290 5.13287
R13916 VDD110.n85 VDD110.n70 5.13287
R13917 VDD110.n86 VDD110.t313 5.13287
R13918 VDD110.n88 VDD110.n68 5.13287
R13919 VDD110.n61 VDD110.t244 5.13287
R13920 VDD110.n144 VDD110.t414 5.13287
R13921 VDD110.n65 VDD110.n64 5.13287
R13922 VDD110.n139 VDD110.t126 5.13287
R13923 VDD110.n138 VDD110.n66 5.13287
R13924 VDD110.n137 VDD110.t61 5.13287
R13925 VDD110.n134 VDD110.n67 5.13287
R13926 VDD110.n516 VDD110.t448 5.13287
R13927 VDD110.n159 VDD110.t285 5.13287
R13928 VDD110.n158 VDD110.n36 5.13287
R13929 VDD110.n157 VDD110.t277 5.13287
R13930 VDD110.n38 VDD110.n37 5.13287
R13931 VDD110.n152 VDD110.t416 5.13287
R13932 VDD110.n151 VDD110.n39 5.13287
R13933 VDD110.n52 VDD110.t120 5.13287
R13934 VDD110.n55 VDD110.t273 5.13287
R13935 VDD110.n57 VDD110.n42 5.13287
R13936 VDD110.n58 VDD110.t30 5.13287
R13937 VDD110.n60 VDD110.n40 5.13287
R13938 VDD110.n26 VDD110.t44 5.13287
R13939 VDD110.n12 VDD110.n11 5.13287
R13940 VDD110.n29 VDD110.t292 5.13287
R13941 VDD110.n527 VDD110.t42 5.13287
R13942 VDD110.n523 VDD110.n522 5.13287
R13943 VDD110 VDD110.n530 5.13104
R13944 VDD110 VDD110.t248 5.10424
R13945 VDD110.n257 VDD110.t230 5.09836
R13946 VDD110.n490 VDD110.t196 5.09407
R13947 VDD110.n492 VDD110.t365 5.09407
R13948 VDD110.n364 VDD110.t208 5.09407
R13949 VDD110.n265 VDD110.t252 5.09407
R13950 VDD110.n270 VDD110.t101 5.09407
R13951 VDD110.n253 VDD110.t268 5.09407
R13952 VDD110.n427 VDD110.t141 5.09407
R13953 VDD110.n451 VDD110.t224 5.09407
R13954 VDD110.n212 VDD110.t77 5.09407
R13955 VDD110.n210 VDD110.t165 5.09407
R13956 VDD110.n500 VDD110.t57 5.09407
R13957 VDD110.n501 VDD110.t490 5.09407
R13958 VDD110.n515 VDD110.t483 5.09407
R13959 VDD110.n132 VDD110.t478 5.09407
R13960 VDD110.n149 VDD110.t488 5.09407
R13961 VDD110.n524 VDD110.t97 5.09407
R13962 VDD110.n0 VDD110.t442 5.09407
R13963 VDD110.n4 VDD110.t343 5.09407
R13964 VDD110.n462 VDD110.n218 5.0055
R13965 VDD110.n446 VDD110.n245 5.0055
R13966 VDD110.n479 VDD110.n478 5.0005
R13967 VDD110.n474 VDD110.n213 5.0005
R13968 VDD110.n472 VDD110.n471 5.0005
R13969 VDD110.n430 VDD110.n248 4.9955
R13970 VDD110.n532 VDD110.n531 4.9917
R13971 VDD110.n470 VDD110.n469 4.9905
R13972 VDD110.n456 VDD110.n455 4.9905
R13973 VDD110.n432 VDD110.n431 4.9905
R13974 VDD110.n454 VDD110.n453 4.9855
R13975 VDD110.n429 VDD110.n428 4.9805
R13976 VDD110.n32 VDD110.t428 4.9655
R13977 VDD110.n485 VDD110 4.91611
R13978 VDD110.n337 VDD110.t14 4.8755
R13979 VDD110.n332 VDD110.n322 4.84121
R13980 VDD110.n481 VDD110.n480 4.7947
R13981 VDD110.n536 VDD110.n535 4.52523
R13982 VDD110.n312 VDD110.n310 4.5005
R13983 VDD110.n313 VDD110.n310 4.5005
R13984 VDD110.n306 VDD110.n304 4.5005
R13985 VDD110.n307 VDD110.n304 4.5005
R13986 VDD110.n325 VDD110.n323 4.5005
R13987 VDD110.n326 VDD110.n323 4.5005
R13988 VDD110.n482 VDD110.n200 4.5005
R13989 VDD110.n481 VDD110.n211 4.5005
R13990 VDD110.n3 VDD110.t325 4.40826
R13991 VDD110.n7 VDD110.t177 4.3915
R13992 VDD110.n1 VDD110.t441 4.26489
R13993 VDD110.n5 VDD110.t342 4.26489
R13994 VDD110.n494 VDD110.t28 4.11379
R13995 VDD110.n258 VDD110.t305 3.94862
R13996 VDD110.n133 VDD110.n88 3.90405
R13997 VDD110 VDD110.n258 3.6765
R13998 VDD110.n208 VDD110.n207 3.1505
R13999 VDD110.n334 VDD110.n333 2.88182
R14000 VDD110.n320 VDD110.n319 2.88074
R14001 VDD110.n205 VDD110.n203 2.85787
R14002 VDD110.n342 VDD110.n299 2.85787
R14003 VDD110.n339 VDD110.n302 2.85787
R14004 VDD110.n360 VDD110.n289 2.85787
R14005 VDD110.n380 VDD110.n370 2.85787
R14006 VDD110.n377 VDD110.n373 2.85787
R14007 VDD110.n400 VDD110.n282 2.85787
R14008 VDD110.n419 VDD110.n409 2.85787
R14009 VDD110.n416 VDD110.n412 2.85787
R14010 VDD110.n444 VDD110.n443 2.85787
R14011 VDD110.n238 VDD110.n228 2.85787
R14012 VDD110.n235 VDD110.n231 2.85787
R14013 VDD110.n473 VDD110.n216 2.85787
R14014 VDD110.n504 VDD110.n192 2.85787
R14015 VDD110.n175 VDD110.n172 2.85787
R14016 VDD110.n178 VDD110.n169 2.85787
R14017 VDD110.n128 VDD110.n91 2.85787
R14018 VDD110.n107 VDD110.n104 2.85787
R14019 VDD110.n110 VDD110.n101 2.85787
R14020 VDD110.n79 VDD110.n76 2.85787
R14021 VDD110.n82 VDD110.n73 2.85787
R14022 VDD110.n145 VDD110.n63 2.85787
R14023 VDD110.n35 VDD110.n34 2.85787
R14024 VDD110.n51 VDD110.n48 2.85787
R14025 VDD110.n54 VDD110.n45 2.85787
R14026 VDD110.n27 VDD110.n10 2.85787
R14027 VDD110.n480 VDD110.n479 2.65128
R14028 VDD110.n537 VDD110.n536 2.55589
R14029 VDD110.n538 VDD110 2.4235
R14030 VDD110.n203 VDD110.t435 2.2755
R14031 VDD110.n203 VDD110.n202 2.2755
R14032 VDD110.n299 VDD110.t369 2.2755
R14033 VDD110.n299 VDD110.n298 2.2755
R14034 VDD110.n302 VDD110.t418 2.2755
R14035 VDD110.n302 VDD110.n301 2.2755
R14036 VDD110.n289 VDD110.t192 2.2755
R14037 VDD110.n289 VDD110.n288 2.2755
R14038 VDD110.n370 VDD110.t111 2.2755
R14039 VDD110.n370 VDD110.n369 2.2755
R14040 VDD110.n373 VDD110.t361 2.2755
R14041 VDD110.n373 VDD110.n372 2.2755
R14042 VDD110.n282 VDD110.t347 2.2755
R14043 VDD110.n282 VDD110.n281 2.2755
R14044 VDD110.n409 VDD110.t388 2.2755
R14045 VDD110.n409 VDD110.n408 2.2755
R14046 VDD110.n412 VDD110.t143 2.2755
R14047 VDD110.n412 VDD110.n411 2.2755
R14048 VDD110.n443 VDD110.t162 2.2755
R14049 VDD110.n443 VDD110.n442 2.2755
R14050 VDD110.n228 VDD110.t424 2.2755
R14051 VDD110.n228 VDD110.n227 2.2755
R14052 VDD110.n231 VDD110.t206 2.2755
R14053 VDD110.n231 VDD110.n230 2.2755
R14054 VDD110.n216 VDD110.t201 2.2755
R14055 VDD110.n216 VDD110.n215 2.2755
R14056 VDD110.n192 VDD110.t179 2.2755
R14057 VDD110.n192 VDD110.n191 2.2755
R14058 VDD110.n172 VDD110.t88 2.2755
R14059 VDD110.n172 VDD110.n171 2.2755
R14060 VDD110.n169 VDD110.t65 2.2755
R14061 VDD110.n169 VDD110.n168 2.2755
R14062 VDD110.n91 VDD110.t336 2.2755
R14063 VDD110.n91 VDD110.n90 2.2755
R14064 VDD110.n104 VDD110.t319 2.2755
R14065 VDD110.n104 VDD110.n103 2.2755
R14066 VDD110.n101 VDD110.t315 2.2755
R14067 VDD110.n101 VDD110.n100 2.2755
R14068 VDD110.n76 VDD110.t49 2.2755
R14069 VDD110.n76 VDD110.n75 2.2755
R14070 VDD110.n73 VDD110.t124 2.2755
R14071 VDD110.n73 VDD110.n72 2.2755
R14072 VDD110.n63 VDD110.t456 2.2755
R14073 VDD110.n63 VDD110.n62 2.2755
R14074 VDD110.n34 VDD110.t440 2.2755
R14075 VDD110.n34 VDD110.n33 2.2755
R14076 VDD110.n48 VDD110.t430 2.2755
R14077 VDD110.n48 VDD110.n47 2.2755
R14078 VDD110.n45 VDD110.t275 2.2755
R14079 VDD110.n45 VDD110.n44 2.2755
R14080 VDD110.n10 VDD110.t476 2.2755
R14081 VDD110.n10 VDD110.n9 2.2755
R14082 VDD110.n502 VDD110 2.25904
R14083 VDD110.n315 VDD110.n314 2.2439
R14084 VDD110.n328 VDD110.n327 2.2439
R14085 VDD110.n309 VDD110.n308 2.24362
R14086 VDD110.n532 VDD110.n528 2.21368
R14087 VDD110.n306 VDD110.n305 2.12277
R14088 VDD110.n330 VDD110.n329 1.82213
R14089 VDD110 VDD110.n287 1.81785
R14090 VDD110.n319 VDD110.n317 1.77234
R14091 VDD110.n321 VDD110.n315 1.6239
R14092 VDD110.n331 VDD110.n328 1.6239
R14093 VDD110.n483 VDD110.n482 1.50339
R14094 VDD110.n325 VDD110.n324 1.39846
R14095 VDD110.n312 VDD110.n311 1.39728
R14096 VDD110.n537 VDD110 1.36829
R14097 VDD110.n349 VDD110.n348 1.16167
R14098 VDD110.n321 VDD110.n320 1.12314
R14099 VDD110.n331 VDD110.n330 1.12224
R14100 VDD110.n387 VDD110.n386 1.07428
R14101 VDD110.n514 VDD110.n184 1.02928
R14102 VDD110.n150 VDD110.n60 1.02928
R14103 VDD110.n426 VDD110.n425 1.01882
R14104 VDD110.n457 VDD110.n244 1.01882
R14105 VDD110.n117 VDD110.n116 0.881662
R14106 VDD110 VDD110.n29 0.819742
R14107 VDD110.n209 VDD110.t27 0.783764
R14108 VDD110.n533 VDD110.n532 0.707829
R14109 VDD110.n521 VDD110.n0 0.66512
R14110 VDD110.n536 VDD110.n528 0.654546
R14111 VDD110.n520 VDD110.n4 0.634017
R14112 VDD110.n332 VDD110.n331 0.52356
R14113 VDD110.n322 VDD110.n309 0.497812
R14114 VDD110.n338 VDD110.n337 0.337997
R14115 VDD110.n337 VDD110.n336 0.333658
R14116 VDD110 VDD110.n519 0.281196
R14117 VDD110.n399 VDD110.n279 0.25039
R14118 VDD110.n343 VDD110.n342 0.233919
R14119 VDD110.n340 VDD110.n339 0.233919
R14120 VDD110.n381 VDD110.n380 0.233919
R14121 VDD110.n378 VDD110.n377 0.233919
R14122 VDD110.n420 VDD110.n419 0.233919
R14123 VDD110.n417 VDD110.n416 0.233919
R14124 VDD110.n239 VDD110.n238 0.233919
R14125 VDD110.n236 VDD110.n235 0.233919
R14126 VDD110.n179 VDD110.n178 0.233919
R14127 VDD110.n176 VDD110.n175 0.233919
R14128 VDD110.n111 VDD110.n110 0.233919
R14129 VDD110.n108 VDD110.n107 0.233919
R14130 VDD110.n83 VDD110.n82 0.233919
R14131 VDD110.n80 VDD110.n79 0.233919
R14132 VDD110.n55 VDD110.n54 0.233919
R14133 VDD110.n52 VDD110.n51 0.233919
R14134 VDD110.n496 VDD110.n495 0.224447
R14135 VDD110.n501 VDD110 0.205357
R14136 VDD110.n497 VDD110.n496 0.202146
R14137 VDD110.n454 VDD110.n245 0.201676
R14138 VDD110.n429 VDD110.n279 0.200832
R14139 VDD110.n430 VDD110.n245 0.183147
R14140 VDD110.n480 VDD110.n212 0.182938
R14141 VDD110.n538 VDD110.n527 0.181055
R14142 VDD110.n431 VDD110.n429 0.1805
R14143 VDD110.n431 VDD110.n430 0.177853
R14144 VDD110.n524 VDD110.n523 0.170231
R14145 VDD110.n515 VDD110.n514 0.167533
R14146 VDD110.n455 VDD110.n218 0.167265
R14147 VDD110 VDD110.n258 0.16613
R14148 VDD110.n455 VDD110.n454 0.161971
R14149 VDD110 VDD110.n61 0.160716
R14150 VDD110.n516 VDD110 0.158984
R14151 VDD110 VDD110.n89 0.157289
R14152 VDD110.n150 VDD110.n149 0.155496
R14153 VDD110.n133 VDD110.n132 0.154581
R14154 VDD110.n534 VDD110 0.153049
R14155 VDD110.n470 VDD110.n218 0.151382
R14156 VDD110 VDD110.n14 0.149922
R14157 VDD110.n471 VDD110.n213 0.148735
R14158 VDD110.n471 VDD110.n470 0.146088
R14159 VDD110.n388 VDD110.n387 0.144547
R14160 VDD110.n521 VDD110.n520 0.142342
R14161 VDD110.n346 VDD110.n345 0.141016
R14162 VDD110.n353 VDD110.n352 0.141016
R14163 VDD110.n354 VDD110.n291 0.141016
R14164 VDD110.n384 VDD110.n383 0.141016
R14165 VDD110.n392 VDD110.n391 0.141016
R14166 VDD110.n393 VDD110.n284 0.141016
R14167 VDD110.n423 VDD110.n422 0.141016
R14168 VDD110.n242 VDD110.n241 0.141016
R14169 VDD110.n182 VDD110.n181 0.141016
R14170 VDD110.n114 VDD110.n113 0.141016
R14171 VDD110.n86 VDD110.n85 0.141016
R14172 VDD110.n58 VDD110.n57 0.141016
R14173 VDD110.n387 VDD110.n364 0.138896
R14174 VDD110.n134 VDD110.n133 0.131861
R14175 VDD110.n500 VDD110.n499 0.130567
R14176 VDD110.n511 VDD110.n510 0.123551
R14177 VDD110.n508 VDD110.n507 0.123551
R14178 VDD110.n138 VDD110.n137 0.123551
R14179 VDD110.n139 VDD110.n65 0.123551
R14180 VDD110 VDD110.n359 0.122435
R14181 VDD110.n479 VDD110.n213 0.122265
R14182 VDD110.n152 VDD110.n38 0.122176
R14183 VDD110.n158 VDD110.n157 0.122176
R14184 VDD110.n121 VDD110.n120 0.120831
R14185 VDD110.n122 VDD110.n93 0.120831
R14186 VDD110.n514 VDD110.n513 0.116432
R14187 VDD110.n151 VDD110.n150 0.115137
R14188 VDD110.n360 VDD110 0.111984
R14189 VDD110.n330 VDD110 0.110941
R14190 VDD110 VDD110.n14 0.107354
R14191 VDD110.n348 VDD110.n347 0.107339
R14192 VDD110.n345 VDD110.n344 0.107339
R14193 VDD110.n351 VDD110.n349 0.107339
R14194 VDD110.n355 VDD110.n353 0.107339
R14195 VDD110.n358 VDD110.n291 0.107339
R14196 VDD110.n386 VDD110.n385 0.107339
R14197 VDD110.n383 VDD110.n382 0.107339
R14198 VDD110.n390 VDD110.n388 0.107339
R14199 VDD110.n394 VDD110.n392 0.107339
R14200 VDD110.n397 VDD110.n284 0.107339
R14201 VDD110.n425 VDD110.n424 0.107339
R14202 VDD110.n422 VDD110.n421 0.107339
R14203 VDD110.n244 VDD110.n243 0.107339
R14204 VDD110.n241 VDD110.n240 0.107339
R14205 VDD110.n499 VDD110.n498 0.107339
R14206 VDD110.n184 VDD110.n183 0.107339
R14207 VDD110.n181 VDD110.n180 0.107339
R14208 VDD110.n116 VDD110.n115 0.107339
R14209 VDD110.n113 VDD110.n112 0.107339
R14210 VDD110.n88 VDD110.n87 0.107339
R14211 VDD110.n85 VDD110.n84 0.107339
R14212 VDD110.n60 VDD110.n59 0.107339
R14213 VDD110.n57 VDD110.n56 0.107339
R14214 VDD110.n526 VDD110.n523 0.107339
R14215 VDD110.n505 VDD110 0.10728
R14216 VDD110 VDD110.n144 0.10728
R14217 VDD110.n342 VDD110 0.106177
R14218 VDD110.n339 VDD110 0.106177
R14219 VDD110 VDD110.n360 0.106177
R14220 VDD110.n380 VDD110 0.106177
R14221 VDD110.n377 VDD110 0.106177
R14222 VDD110.n419 VDD110 0.106177
R14223 VDD110.n416 VDD110 0.106177
R14224 VDD110.n238 VDD110 0.106177
R14225 VDD110.n235 VDD110 0.106177
R14226 VDD110.n178 VDD110 0.106177
R14227 VDD110.n175 VDD110 0.106177
R14228 VDD110.n110 VDD110 0.106177
R14229 VDD110.n107 VDD110 0.106177
R14230 VDD110.n82 VDD110 0.106177
R14231 VDD110.n79 VDD110 0.106177
R14232 VDD110.n54 VDD110 0.106177
R14233 VDD110.n51 VDD110 0.106177
R14234 VDD110.n159 VDD110 0.106087
R14235 VDD110 VDD110.n538 0.105243
R14236 VDD110 VDD110.n127 0.10492
R14237 VDD110 VDD110.n504 0.0981271
R14238 VDD110.n145 VDD110 0.0981271
R14239 VDD110 VDD110.n35 0.0970363
R14240 VDD110.n521 VDD110.n3 0.096125
R14241 VDD110.n128 VDD110 0.0959696
R14242 VDD110.n23 VDD110 0.0956733
R14243 VDD110.n513 VDD110.n512 0.0940593
R14244 VDD110.n510 VDD110.n509 0.0940593
R14245 VDD110.n507 VDD110.n506 0.0940593
R14246 VDD110.n136 VDD110.n134 0.0940593
R14247 VDD110.n140 VDD110.n138 0.0940593
R14248 VDD110.n143 VDD110.n65 0.0940593
R14249 VDD110.n504 VDD110 0.0930424
R14250 VDD110 VDD110.n145 0.0930424
R14251 VDD110.n153 VDD110.n151 0.093014
R14252 VDD110.n156 VDD110.n38 0.093014
R14253 VDD110.n160 VDD110.n158 0.093014
R14254 VDD110.n119 VDD110.n117 0.0919917
R14255 VDD110.n123 VDD110.n121 0.0919917
R14256 VDD110.n126 VDD110.n93 0.0919917
R14257 VDD110 VDD110.n128 0.0909972
R14258 VDD110.n520 VDD110.n7 0.0905
R14259 VDD110 VDD110.n255 0.084523
R14260 VDD110.n272 VDD110 0.084523
R14261 VDD110 VDD110.n257 0.0842767
R14262 VDD110.n318 VDD110 0.0839415
R14263 VDD110.n279 VDD110.n278 0.0826283
R14264 VDD110.n496 VDD110.n200 0.0819374
R14265 VDD110.n27 VDD110.n26 0.0817097
R14266 VDD110.n313 VDD110 0.0816915
R14267 VDD110.n478 VDD110.n214 0.0816286
R14268 VDD110.n341 VDD110.n340 0.080629
R14269 VDD110.n361 VDD110.n287 0.080629
R14270 VDD110.n379 VDD110.n378 0.080629
R14271 VDD110.n418 VDD110.n417 0.080629
R14272 VDD110.n237 VDD110.n236 0.080629
R14273 VDD110.n177 VDD110.n176 0.080629
R14274 VDD110.n109 VDD110.n108 0.080629
R14275 VDD110.n81 VDD110.n80 0.080629
R14276 VDD110.n53 VDD110.n52 0.080629
R14277 VDD110.n326 VDD110 0.0805665
R14278 VDD110 VDD110.n346 0.0794677
R14279 VDD110 VDD110.n343 0.0794677
R14280 VDD110.n352 VDD110 0.0794677
R14281 VDD110 VDD110.n354 0.0794677
R14282 VDD110.n359 VDD110 0.0794677
R14283 VDD110 VDD110.n384 0.0794677
R14284 VDD110 VDD110.n381 0.0794677
R14285 VDD110.n391 VDD110 0.0794677
R14286 VDD110 VDD110.n393 0.0794677
R14287 VDD110 VDD110.n423 0.0794677
R14288 VDD110 VDD110.n420 0.0794677
R14289 VDD110 VDD110.n242 0.0794677
R14290 VDD110 VDD110.n239 0.0794677
R14291 VDD110 VDD110.n182 0.0794677
R14292 VDD110 VDD110.n179 0.0794677
R14293 VDD110 VDD110.n114 0.0794677
R14294 VDD110 VDD110.n111 0.0794677
R14295 VDD110 VDD110.n86 0.0794677
R14296 VDD110 VDD110.n83 0.0794677
R14297 VDD110 VDD110.n58 0.0794677
R14298 VDD110 VDD110.n55 0.0794677
R14299 VDD110.n398 VDD110 0.0765085
R14300 VDD110.n527 VDD110 0.0759839
R14301 VDD110.n307 VDD110 0.0738165
R14302 VDD110.n336 VDD110.n334 0.0725
R14303 VDD110.n490 VDD110 0.0709717
R14304 VDD110.n364 VDD110 0.0709717
R14305 VDD110.n210 VDD110 0.0709717
R14306 VDD110 VDD110.n501 0.0709717
R14307 VDD110 VDD110.n524 0.0709717
R14308 VDD110 VDD110.n0 0.0709717
R14309 VDD110 VDD110.n4 0.0709717
R14310 VDD110.n503 VDD110.n502 0.0706695
R14311 VDD110.n146 VDD110.n61 0.0706695
R14312 VDD110.n517 VDD110.n516 0.0698855
R14313 VDD110 VDD110.n511 0.0696525
R14314 VDD110 VDD110.n508 0.0696525
R14315 VDD110 VDD110.n505 0.0696525
R14316 VDD110.n137 VDD110 0.0696525
R14317 VDD110 VDD110.n139 0.0696525
R14318 VDD110.n144 VDD110 0.0696525
R14319 VDD110.n129 VDD110.n89 0.0691188
R14320 VDD110 VDD110.n152 0.0688799
R14321 VDD110.n157 VDD110 0.0688799
R14322 VDD110 VDD110.n159 0.0688799
R14323 VDD110.n120 VDD110 0.0681243
R14324 VDD110 VDD110.n122 0.0681243
R14325 VDD110.n127 VDD110 0.0681243
R14326 VDD110.n335 VDD110 0.0659545
R14327 VDD110.n435 VDD110.n434 0.0647478
R14328 VDD110.n441 VDD110.n440 0.0647478
R14329 VDD110.n266 VDD110.n265 0.0618169
R14330 VDD110.n271 VDD110.n270 0.0618169
R14331 VDD110.n253 VDD110.n252 0.0618169
R14332 VDD110.n426 VDD110.n250 0.0607039
R14333 VDD110.n458 VDD110.n457 0.0607039
R14334 VDD110.n262 VDD110.n261 0.0599607
R14335 VDD110.n469 VDD110.n468 0.0597035
R14336 VDD110.n463 VDD110.n462 0.0586416
R14337 VDD110.n445 VDD110 0.0562522
R14338 VDD110 VDD110.n13 0.0559424
R14339 VDD110 VDD110.n494 0.0555633
R14340 VDD110 VDD110.n497 0.0550806
R14341 VDD110.n427 VDD110.n426 0.0536232
R14342 VDD110 VDD110.n205 0.0533387
R14343 VDD110.n518 VDD110.n35 0.0532933
R14344 VDD110 VDD110.n472 0.0522699
R14345 VDD110.n261 VDD110 0.0518708
R14346 VDD110.n400 VDD110 0.0514734
R14347 VDD110 VDD110.n444 0.0514734
R14348 VDD110.n473 VDD110 0.0514734
R14349 VDD110.n447 VDD110.n441 0.0493496
R14350 VDD110.n460 VDD110.n458 0.0493496
R14351 VDD110.n464 VDD110.n463 0.0493496
R14352 VDD110.n468 VDD110.n467 0.0493496
R14353 VDD110 VDD110.n400 0.0488186
R14354 VDD110.n436 VDD110.n432 0.0488186
R14355 VDD110.n444 VDD110 0.0488186
R14356 VDD110.n267 VDD110.n266 0.0487799
R14357 VDD110.n273 VDD110.n271 0.0487799
R14358 VDD110.n277 VDD110.n252 0.0487799
R14359 VDD110.n428 VDD110.n280 0.046557
R14360 VDD110.n336 VDD110.n335 0.0455
R14361 VDD110.n20 VDD110.n19 0.0446736
R14362 VDD110 VDD110.n12 0.0444695
R14363 VDD110.n474 VDD110.n473 0.0437743
R14364 VDD110 VDD110.n500 0.043431
R14365 VDD110.n149 VDD110 0.0404465
R14366 VDD110 VDD110.n515 0.0400238
R14367 VDD110.n132 VDD110 0.0396099
R14368 VDD110.n428 VDD110 0.0394398
R14369 VDD110.n518 VDD110 0.0392151
R14370 VDD110.n451 VDD110 0.039182
R14371 VDD110.n19 VDD110 0.0386636
R14372 VDD110 VDD110.n206 0.0382419
R14373 VDD110.n452 VDD110 0.0377891
R14374 VDD110.n399 VDD110.n398 0.0371957
R14375 VDD110.n401 VDD110.n280 0.0371372
R14376 VDD110.n475 VDD110.n214 0.0371372
R14377 VDD110 VDD110.n435 0.0366062
R14378 VDD110.n440 VDD110 0.0366062
R14379 VDD110.n461 VDD110 0.0366062
R14380 VDD110 VDD110.n219 0.0366062
R14381 VDD110 VDD110.n217 0.0366062
R14382 VDD110 VDD110.n257 0.0350843
R14383 VDD110 VDD110.n255 0.0346108
R14384 VDD110 VDD110.n272 0.0346108
R14385 VDD110.n278 VDD110 0.0346108
R14386 VDD110.n491 VDD110.n205 0.0344677
R14387 VDD110.n484 VDD110.n210 0.0327642
R14388 VDD110 VDD110.n492 0.032019
R14389 VDD110.n31 VDD110.n8 0.0319625
R14390 VDD110.n434 VDD110.n248 0.0291726
R14391 VDD110 VDD110.n8 0.0276819
R14392 VDD110.n314 VDD110.n313 0.0275
R14393 VDD110.n318 VDD110.n316 0.0275
R14394 VDD110.n446 VDD110.n445 0.0265177
R14395 VDD110.n327 VDD110.n326 0.026375
R14396 VDD110.n25 VDD110.n12 0.0257824
R14397 VDD110.n315 VDD110.n310 0.025705
R14398 VDD110.n328 VDD110.n323 0.025705
R14399 VDD110 VDD110.n27 0.0256227
R14400 VDD110.n453 VDD110.n246 0.0233319
R14401 VDD110.n211 VDD110.n200 0.0225755
R14402 VDD110 VDD110.n427 0.021904
R14403 VDD110 VDD110.n451 0.021904
R14404 VDD110 VDD110.n212 0.021904
R14405 VDD110.n265 VDD110 0.0216615
R14406 VDD110.n270 VDD110 0.0216615
R14407 VDD110 VDD110.n253 0.0216615
R14408 VDD110 VDD110.n399 0.0214735
R14409 VDD110.n308 VDD110.n307 0.02075
R14410 VDD110.n439 VDD110.n248 0.020677
R14411 VDD110.n29 VDD110.n28 0.0195491
R14412 VDD110.n482 VDD110.n481 0.0193811
R14413 VDD110.n32 VDD110 0.0184587
R14414 VDD110.n26 VDD110 0.0183626
R14415 VDD110.n535 VDD110.n529 0.0177727
R14416 VDD110.n309 VDD110.n304 0.0169383
R14417 VDD110.n520 VDD110 0.0147612
R14418 VDD110.n453 VDD110.n452 0.0143053
R14419 VDD110.n519 VDD110.n32 0.0137976
R14420 VDD110 VDD110.n14 0.0127264
R14421 VDD110.n457 VDD110.n456 0.0126203
R14422 VDD110 VDD110.n446 0.0105885
R14423 VDD110.n308 VDD110.n306 0.0095
R14424 VDD110.n335 VDD110 0.00868182
R14425 VDD110.n462 VDD110.n461 0.00660619
R14426 VDD110 VDD110.n521 0.00608887
R14427 VDD110.n469 VDD110.n219 0.00554425
R14428 VDD110 VDD110.n474 0.00554425
R14429 VDD110.n494 VDD110 0.00543671
R14430 VDD110.n498 VDD110 0.00514516
R14431 VDD110 VDD110.n526 0.00514516
R14432 VDD110 VDD110.n13 0.00485726
R14433 VDD110.n472 VDD110.n217 0.0044823
R14434 VDD110.n478 VDD110 0.00436819
R14435 VDD110.n327 VDD110.n325 0.003875
R14436 VDD110.n495 VDD110 0.00315823
R14437 VDD110.n207 VDD110 0.00282258
R14438 VDD110.n456 VDD110 0.00282092
R14439 VDD110.n314 VDD110.n312 0.00275
R14440 VDD110.n267 VDD110 0.00259913
R14441 VDD110.n273 VDD110 0.00259913
R14442 VDD110 VDD110.n277 0.00259913
R14443 VDD110.n529 VDD110.n528 0.00231818
R14444 VDD110.n535 VDD110.n534 0.00231818
R14445 VDD110.n320 VDD110.n316 0.00171994
R14446 VDD110.n347 VDD110 0.00166129
R14447 VDD110.n344 VDD110 0.00166129
R14448 VDD110 VDD110.n341 0.00166129
R14449 VDD110 VDD110.n338 0.00166129
R14450 VDD110 VDD110.n351 0.00166129
R14451 VDD110.n355 VDD110 0.00166129
R14452 VDD110 VDD110.n358 0.00166129
R14453 VDD110.n361 VDD110 0.00166129
R14454 VDD110.n385 VDD110 0.00166129
R14455 VDD110.n382 VDD110 0.00166129
R14456 VDD110 VDD110.n379 0.00166129
R14457 VDD110 VDD110.n376 0.00166129
R14458 VDD110 VDD110.n390 0.00166129
R14459 VDD110.n394 VDD110 0.00166129
R14460 VDD110 VDD110.n397 0.00166129
R14461 VDD110.n424 VDD110 0.00166129
R14462 VDD110.n421 VDD110 0.00166129
R14463 VDD110 VDD110.n418 0.00166129
R14464 VDD110 VDD110.n415 0.00166129
R14465 VDD110.n243 VDD110 0.00166129
R14466 VDD110.n240 VDD110 0.00166129
R14467 VDD110 VDD110.n237 0.00166129
R14468 VDD110 VDD110.n234 0.00166129
R14469 VDD110.n183 VDD110 0.00166129
R14470 VDD110.n180 VDD110 0.00166129
R14471 VDD110 VDD110.n177 0.00166129
R14472 VDD110 VDD110.n174 0.00166129
R14473 VDD110.n115 VDD110 0.00166129
R14474 VDD110.n112 VDD110 0.00166129
R14475 VDD110 VDD110.n109 0.00166129
R14476 VDD110 VDD110.n106 0.00166129
R14477 VDD110.n87 VDD110 0.00166129
R14478 VDD110.n84 VDD110 0.00166129
R14479 VDD110 VDD110.n81 0.00166129
R14480 VDD110 VDD110.n78 0.00166129
R14481 VDD110.n59 VDD110 0.00166129
R14482 VDD110.n56 VDD110 0.00166129
R14483 VDD110 VDD110.n53 0.00166129
R14484 VDD110 VDD110.n50 0.00166129
R14485 VDD110 VDD110.n25 0.00159924
R14486 VDD110.n484 VDD110.n483 0.00156548
R14487 VDD110.n512 VDD110 0.00151695
R14488 VDD110.n509 VDD110 0.00151695
R14489 VDD110.n506 VDD110 0.00151695
R14490 VDD110 VDD110.n503 0.00151695
R14491 VDD110 VDD110.n136 0.00151695
R14492 VDD110.n140 VDD110 0.00151695
R14493 VDD110 VDD110.n143 0.00151695
R14494 VDD110.n146 VDD110 0.00151695
R14495 VDD110.n153 VDD110 0.00150559
R14496 VDD110 VDD110.n156 0.00150559
R14497 VDD110.n160 VDD110 0.00150559
R14498 VDD110 VDD110.n517 0.00150559
R14499 VDD110 VDD110.n119 0.00149448
R14500 VDD110.n123 VDD110 0.00149448
R14501 VDD110 VDD110.n126 0.00149448
R14502 VDD110.n129 VDD110 0.00149448
R14503 VDD110.n483 VDD110.n211 0.00128347
R14504 VDD110.n207 VDD110 0.00108064
R14505 VDD110.n401 VDD110 0.00103097
R14506 VDD110.n432 VDD110.n250 0.00103097
R14507 VDD110.n436 VDD110 0.00103097
R14508 VDD110 VDD110.n439 0.00103097
R14509 VDD110.n447 VDD110 0.00103097
R14510 VDD110 VDD110.n246 0.00103097
R14511 VDD110 VDD110.n460 0.00103097
R14512 VDD110.n464 VDD110 0.00103097
R14513 VDD110.n467 VDD110 0.00103097
R14514 VDD110.n475 VDD110 0.00103097
R14515 VDD110.n16 VDD110 0.00100943
R14516 VDD110.n262 VDD110 0.000904494
R14517 VDD110.n20 VDD110 0.000800501
R14518 VDD110.n28 VDD110 0.000776074
R14519 VDD110 VDD110.n23 0.000774809
R14520 VDD110 VDD110.n31 0.000714031
R14521 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n20 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t24 36.935
R14522 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n19 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t16 36.935
R14523 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n30 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t14 36.935
R14524 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n29 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t7 36.935
R14525 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n28 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t25 36.935
R14526 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n26 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t27 36.935
R14527 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n25 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t19 36.935
R14528 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n23 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t17 36.935
R14529 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n22 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t20 36.935
R14530 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n21 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t9 25.5364
R14531 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n27 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t22 25.5364
R14532 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n24 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t18 25.5364
R14533 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n31 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t5 25.5361
R14534 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n20 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t10 18.1962
R14535 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n19 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t2 18.1962
R14536 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n30 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t23 18.1962
R14537 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n29 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t15 18.1962
R14538 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n28 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t8 18.1962
R14539 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n26 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t12 18.1962
R14540 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n25 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t4 18.1962
R14541 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n23 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t3 18.1962
R14542 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n22 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t6 18.1962
R14543 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n27 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t13 14.0749
R14544 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n24 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t11 14.0749
R14545 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n21 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t26 14.0749
R14546 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n31 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t21 14.0734
R14547 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n18 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t0 9.33985
R14548 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n33 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3 5.77906
R14549 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n18 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t1 5.17836
R14550 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n35 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n34 5.11659
R14551 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n10 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n19 2.13042
R14552 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n3 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n2 1.11863
R14553 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n11 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n29 2.13042
R14554 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n5 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n4 1.11863
R14555 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n14 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n31 1.43628
R14556 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n0 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n32 4.94724
R14557 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n12 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n25 2.13042
R14558 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n7 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n6 1.11863
R14559 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n15 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n27 1.43559
R14560 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n13 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n22 2.13042
R14561 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n9 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n8 1.11863
R14562 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n16 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n24 1.43559
R14563 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n1 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n17 1.49204
R14564 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n36 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n35 4.5005
R14565 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n34 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3 4.43149
R14566 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n33 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n32 3.5258
R14567 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n32 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3 2.3355
R14568 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n3 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n20 2.13151
R14569 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n5 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n30 2.13151
R14570 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n7 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n26 2.13151
R14571 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n9 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n23 2.13151
R14572 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n2 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n10 2.63808
R14573 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n4 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n11 2.63808
R14574 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n6 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n12 2.63808
R14575 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n8 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n13 2.63808
R14576 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n16 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n8 2.10738
R14577 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n15 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n6 2.10738
R14578 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n14 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n4 2.10738
R14579 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n34 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n33 1.62556
R14580 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n17 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n21 1.42706
R14581 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n2 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n1 0.991659
R14582 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n36 0.1705
R14583 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n18 0.115328
R14584 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n0 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3 0.0684998
R14585 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n3 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3 0.0786548
R14586 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n10 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3 0.0807313
R14587 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n5 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3 0.0786548
R14588 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n11 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3 0.0807313
R14589 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n7 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3 0.0786548
R14590 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n12 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3 0.0807313
R14591 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n9 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3 0.0786548
R14592 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n13 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3 0.0807313
R14593 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n36 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n17 0.033
R14594 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n16 0.1953
R14595 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n15 0.1953
R14596 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n14 0.1953
R14597 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n35 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n1 0.0170403
R14598 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n0 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n28 2.14709
R14599 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t5 37.1986
R14600 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t3 31.528
R14601 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n3 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t6 30.6315
R14602 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n3 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t7 24.5953
R14603 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t4 17.6614
R14604 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n4 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 17.0516
R14605 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t8 15.3826
R14606 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n1 7.62751
R14607 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n5 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n4 3.28711
R14608 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n7 2.99416
R14609 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n4 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 2.81128
R14610 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n5 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 2.67866
R14611 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n7 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t0 2.2755
R14612 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n7 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n6 2.2755
R14613 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n5 2.2505
R14614 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n3 1.80496
R14615 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n2 1.43709
R14616 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n0 0.281955
R14617 VDD108.n157 VDD108.t407 107239
R14618 VDD108.n352 VDD108.t367 107239
R14619 VDD108.t34 VDD108.n260 57397.6
R14620 VDD108.n350 VDD108.n334 4006.3
R14621 VDD108.n155 VDD108.n139 4006.3
R14622 VDD108.n157 VDD108.n137 3116.02
R14623 VDD108.n352 VDD108.n332 3116.02
R14624 VDD108.n156 VDD108.n137 2331.49
R14625 VDD108.n351 VDD108.n332 2331.49
R14626 VDD108.n156 VDD108.n155 1668.51
R14627 VDD108.n351 VDD108.n350 1668.51
R14628 VDD108.t171 VDD108.t410 1164.27
R14629 VDD108.t231 VDD108.t333 1164.27
R14630 VDD108.t44 VDD108.t369 1164.27
R14631 VDD108.t7 VDD108.t68 1164.27
R14632 VDD108.t317 VDD108.n156 1046.11
R14633 VDD108.t277 VDD108.n351 1046.11
R14634 VDD108.t47 VDD108.t153 961.905
R14635 VDD108.t288 VDD108.t161 961.905
R14636 VDD108.n260 VDD108.t83 864.287
R14637 VDD108.t434 VDD108.t240 765.152
R14638 VDD108.t258 VDD108.t253 765.152
R14639 VDD108.t426 VDD108.t174 765.152
R14640 VDD108.t303 VDD108.t282 765.152
R14641 VDD108.t206 VDD108.t200 765.152
R14642 VDD108.t198 VDD108.t196 765.152
R14643 VDD108.t285 VDD108.t60 765.152
R14644 VDD108.t202 VDD108.t204 765.152
R14645 VDD108.t212 VDD108.t55 765.152
R14646 VDD108.t126 VDD108.t123 765.152
R14647 VDD108.t129 VDD108.t138 765.152
R14648 VDD108.t155 VDD108.t244 765.152
R14649 VDD108.t163 VDD108.t106 765.152
R14650 VDD108.t168 VDD108.t234 765.152
R14651 VDD108.t140 VDD108.t72 765.152
R14652 VDD108.t116 VDD108.t150 765.152
R14653 VDD108.t166 VDD108.t237 765.152
R14654 VDD108.t76 VDD108.t74 765.152
R14655 VDD108.t50 VDD108.t53 765.152
R14656 VDD108.t85 VDD108.t79 765.152
R14657 VDD108.t363 VDD108.t365 765.152
R14658 VDD108.t179 VDD108.t260 765.152
R14659 VDD108.t263 VDD108.t280 765.152
R14660 VDD108.t326 VDD108.t70 765.152
R14661 VDD108.t393 VDD108.t191 765.152
R14662 VDD108.t189 VDD108.t274 765.152
R14663 VDD108.t227 VDD108.t358 765.152
R14664 VDD108.t396 VDD108.t146 765.152
R14665 VDD108.t187 VDD108.t272 765.152
R14666 VDD108.t62 VDD108.t301 765.152
R14667 VDD108.t404 VDD108.t269 765.152
R14668 VDD108.t315 VDD108.t323 765.152
R14669 VDD108.t331 VDD108.t335 765.152
R14670 VDD108.t298 VDD108.t214 765.152
R14671 VDD108.t132 VDD108.t135 765.152
R14672 VDD108.t184 VDD108.t242 765.152
R14673 VDD108.t431 VDD108.t249 765.152
R14674 VDD108.t256 VDD108.t251 765.152
R14675 VDD108.t424 VDD108.t329 765.152
R14676 VDD108.t444 VDD108.t37 461.096
R14677 VDD108.t410 VDD108.t444 461.096
R14678 VDD108.t356 VDD108.t171 461.096
R14679 VDD108.t320 VDD108.t356 461.096
R14680 VDD108.t333 VDD108.t317 461.096
R14681 VDD108.t407 VDD108.t231 461.096
R14682 VDD108.t376 VDD108.t41 461.096
R14683 VDD108.t369 VDD108.t376 461.096
R14684 VDD108.t347 VDD108.t44 461.096
R14685 VDD108.t266 VDD108.t347 461.096
R14686 VDD108.t68 VDD108.t277 461.096
R14687 VDD108.t367 VDD108.t7 461.096
R14688 VDD108 VDD108.n196 429.187
R14689 VDD108.n325 VDD108 429.187
R14690 VDD108 VDD108.n108 429.187
R14691 VDD108 VDD108.n64 429.187
R14692 VDD108 VDD108.n442 429.187
R14693 VDD108 VDD108.n462 429.187
R14694 VDD108 VDD108.n301 427.092
R14695 VDD108 VDD108.n119 427.092
R14696 VDD108 VDD108.n303 426.699
R14697 VDD108 VDD108.n373 426.699
R14698 VDD108 VDD108.n192 424.618
R14699 VDD108 VDD108.n292 420.935
R14700 VDD108 VDD108.n115 420.935
R14701 VDD108.n208 VDD108 418.495
R14702 VDD108.n442 VDD108.t11 386.365
R14703 VDD108.t399 VDD108.n64 386.365
R14704 VDD108.n196 VDD108.t176 386.365
R14705 VDD108.n303 VDD108.t229 386.365
R14706 VDD108.t113 VDD108.n325 386.365
R14707 VDD108.n373 VDD108.t290 386.365
R14708 VDD108.t219 VDD108.n108 386.365
R14709 VDD108.t81 VDD108.t349 380.952
R14710 VDD108.t103 VDD108.t288 380.952
R14711 VDD108.t292 VDD108.n208 378.788
R14712 VDD108.n292 VDD108.t111 378.788
R14713 VDD108.n115 VDD108.t222 378.788
R14714 VDD108.n208 VDD108.t0 322.223
R14715 VDD108.t57 VDD108.n292 322.223
R14716 VDD108.t246 VDD108.n115 322.223
R14717 VDD108.n192 VDD108.t67 320.635
R14718 VDD108.n301 VDD108.t372 320.635
R14719 VDD108.n119 VDD108.t409 320.635
R14720 VDD108.t307 VDD108.t426 303.031
R14721 VDD108.t196 VDD108.t418 303.031
R14722 VDD108.t344 VDD108.t202 303.031
R14723 VDD108.t413 VDD108.t212 303.031
R14724 VDD108.t123 VDD108.t452 303.031
R14725 VDD108.t106 VDD108.t386 303.031
R14726 VDD108.t234 VDD108.t354 303.031
R14727 VDD108.t150 VDD108.t381 303.031
R14728 VDD108.t98 VDD108.t363 303.031
R14729 VDD108.t391 VDD108.t179 303.031
R14730 VDD108.t90 VDD108.t227 303.031
R14731 VDD108.t338 VDD108.t187 303.031
R14732 VDD108.t93 VDD108.t62 303.031
R14733 VDD108.t437 VDD108.t404 303.031
R14734 VDD108.t214 VDD108.t442 303.031
R14735 VDD108.t352 VDD108.t132 303.031
R14736 VDD108.t341 VDD108.t256 303.031
R14737 VDD108.t310 VDD108.t424 303.031
R14738 VDD108.n252 VDD108.t295 242.857
R14739 VDD108.n254 VDD108.t47 242.857
R14740 VDD108.t349 VDD108.n257 242.857
R14741 VDD108.n261 VDD108.t103 242.857
R14742 VDD108.n447 VDD108.t428 193.183
R14743 VDD108.n448 VDD108.t434 193.183
R14744 VDD108.n457 VDD108.t253 193.183
R14745 VDD108.n458 VDD108.t307 193.183
R14746 VDD108.n428 VDD108.t193 193.183
R14747 VDD108.n434 VDD108.t282 193.183
R14748 VDD108.n435 VDD108.t206 193.183
R14749 VDD108.n441 VDD108.t418 193.183
R14750 VDD108.n38 VDD108.t209 193.183
R14751 VDD108.n40 VDD108.t285 193.183
R14752 VDD108.n43 VDD108.t344 193.183
R14753 VDD108.n46 VDD108.t413 193.183
R14754 VDD108.n209 VDD108.t292 193.183
R14755 VDD108.n286 VDD108.t360 193.183
R14756 VDD108.n289 VDD108.t50 193.183
R14757 VDD108.n294 VDD108.t85 193.183
R14758 VDD108.n299 VDD108.t98 193.183
R14759 VDD108.n242 VDD108.t224 193.183
R14760 VDD108.n243 VDD108.t393 193.183
R14761 VDD108.n249 VDD108.t274 193.183
R14762 VDD108.n250 VDD108.t90 193.183
R14763 VDD108.n219 VDD108.t64 193.183
R14764 VDD108.n221 VDD108.t396 193.183
R14765 VDD108.n224 VDD108.t338 193.183
R14766 VDD108.n227 VDD108.t93 193.183
R14767 VDD108.n5 VDD108.t421 193.183
R14768 VDD108.n7 VDD108.t431 193.183
R14769 VDD108.n10 VDD108.t341 193.183
R14770 VDD108.n13 VDD108.t310 193.183
R14771 VDD108.t452 VDD108.n66 191.288
R14772 VDD108.t138 VDD108.n70 191.288
R14773 VDD108.t244 VDD108.n72 191.288
R14774 VDD108.n74 VDD108.t121 191.288
R14775 VDD108.t386 VDD108.n170 191.288
R14776 VDD108.t354 VDD108.n174 191.288
R14777 VDD108.t72 VDD108.n178 191.288
R14778 VDD108.n180 VDD108.t109 191.288
R14779 VDD108.t381 VDD108.n200 191.288
R14780 VDD108.n201 VDD108.t166 191.288
R14781 VDD108.t74 VDD108.n383 191.288
R14782 VDD108.n384 VDD108.t148 191.288
R14783 VDD108.t111 VDD108.n290 191.288
R14784 VDD108.n364 VDD108.t391 191.288
R14785 VDD108.n363 VDD108.t280 191.288
R14786 VDD108.t70 VDD108.n329 191.288
R14787 VDD108.n331 VDD108.t182 191.288
R14788 VDD108.n406 VDD108.t437 191.288
R14789 VDD108.n405 VDD108.t315 191.288
R14790 VDD108.n404 VDD108.t331 191.288
R14791 VDD108.n403 VDD108.t402 191.288
R14792 VDD108.t222 VDD108.n113 191.288
R14793 VDD108.t442 VDD108.n94 191.288
R14794 VDD108.n95 VDD108.t352 191.288
R14795 VDD108.t242 VDD108.n103 191.288
R14796 VDD108.n104 VDD108.t217 191.288
R14797 VDD108.n207 VDD108.t67 142.857
R14798 VDD108.t372 VDD108.n296 142.857
R14799 VDD108.t409 VDD108.n117 142.857
R14800 VDD108.t153 VDD108.n252 138.095
R14801 VDD108.t83 VDD108.n254 138.095
R14802 VDD108.t161 VDD108.n257 138.095
R14803 VDD108.n261 VDD108.t34 138.095
R14804 VDD108.n156 VDD108.t320 118.156
R14805 VDD108.n351 VDD108.t266 118.156
R14806 VDD108.n66 VDD108.t399 111.743
R14807 VDD108.n70 VDD108.t126 111.743
R14808 VDD108.n72 VDD108.t129 111.743
R14809 VDD108.n74 VDD108.t155 111.743
R14810 VDD108.n170 VDD108.t27 111.743
R14811 VDD108.n174 VDD108.t163 111.743
R14812 VDD108.n178 VDD108.t168 111.743
R14813 VDD108.n180 VDD108.t140 111.743
R14814 VDD108.n200 VDD108.t176 111.743
R14815 VDD108.n201 VDD108.t116 111.743
R14816 VDD108.n383 VDD108.t237 111.743
R14817 VDD108.n384 VDD108.t76 111.743
R14818 VDD108.n290 VDD108.t383 111.743
R14819 VDD108.n364 VDD108.t113 111.743
R14820 VDD108.t260 VDD108.n363 111.743
R14821 VDD108.n329 VDD108.t263 111.743
R14822 VDD108.n331 VDD108.t326 111.743
R14823 VDD108.n406 VDD108.t219 111.743
R14824 VDD108.t269 VDD108.n405 111.743
R14825 VDD108.t323 VDD108.n404 111.743
R14826 VDD108.t335 VDD108.n403 111.743
R14827 VDD108.n113 VDD108.t449 111.743
R14828 VDD108.n94 VDD108.t14 111.743
R14829 VDD108.n95 VDD108.t298 111.743
R14830 VDD108.n103 VDD108.t135 111.743
R14831 VDD108.n104 VDD108.t184 111.743
R14832 VDD108.t0 VDD108.n207 111.112
R14833 VDD108.n296 VDD108.t57 111.112
R14834 VDD108.n117 VDD108.t246 111.112
R14835 VDD108.t240 VDD108.n447 109.849
R14836 VDD108.n448 VDD108.t258 109.849
R14837 VDD108.t174 VDD108.n457 109.849
R14838 VDD108.n458 VDD108.t18 109.849
R14839 VDD108.n428 VDD108.t303 109.849
R14840 VDD108.t200 VDD108.n434 109.849
R14841 VDD108.n435 VDD108.t198 109.849
R14842 VDD108.t11 VDD108.n441 109.849
R14843 VDD108.t60 VDD108.n38 109.849
R14844 VDD108.t204 VDD108.n40 109.849
R14845 VDD108.t55 VDD108.n43 109.849
R14846 VDD108.n46 VDD108.t24 109.849
R14847 VDD108.n209 VDD108.t96 109.849
R14848 VDD108.t53 VDD108.n286 109.849
R14849 VDD108.t79 VDD108.n289 109.849
R14850 VDD108.t365 VDD108.n294 109.849
R14851 VDD108.t229 VDD108.n299 109.849
R14852 VDD108.t191 VDD108.n242 109.849
R14853 VDD108.n243 VDD108.t189 109.849
R14854 VDD108.t358 VDD108.n249 109.849
R14855 VDD108.t290 VDD108.n250 109.849
R14856 VDD108.t146 VDD108.n219 109.849
R14857 VDD108.t272 VDD108.n221 109.849
R14858 VDD108.t301 VDD108.n224 109.849
R14859 VDD108.n227 VDD108.t21 109.849
R14860 VDD108.t249 VDD108.n5 109.849
R14861 VDD108.t251 VDD108.n7 109.849
R14862 VDD108.t329 VDD108.n10 109.849
R14863 VDD108.n13 VDD108.t31 109.849
R14864 VDD108.n260 VDD108.t81 97.6195
R14865 VDD108.n303 VDD108.t101 62.1896
R14866 VDD108.n373 VDD108.t88 62.1896
R14867 VDD108.n192 VDD108.t305 61.8817
R14868 VDD108.n208 VDD108.t5 60.9761
R14869 VDD108.n462 VDD108.t313 59.702
R14870 VDD108.n442 VDD108.t416 59.702
R14871 VDD108.n64 VDD108.t446 59.702
R14872 VDD108.n196 VDD108.t378 59.702
R14873 VDD108.n325 VDD108.t388 59.702
R14874 VDD108.n108 VDD108.t439 59.702
R14875 VDD108.n301 VDD108.t2 59.4064
R14876 VDD108.n119 VDD108.t143 59.4064
R14877 VDD108.n292 VDD108.t373 58.5371
R14878 VDD108.n115 VDD108.t158 58.5371
R14879 VDD108.n49 VDD108.t23 30.9379
R14880 VDD108.n47 VDD108.t10 30.9379
R14881 VDD108.n264 VDD108.t20 30.9379
R14882 VDD108.n162 VDD108.t40 30.9379
R14883 VDD108.n82 VDD108.t36 30.9379
R14884 VDD108.n14 VDD108.t17 30.9379
R14885 VDD108.n15 VDD108.t30 30.9379
R14886 VDD108.n165 VDD108.t26 30.3459
R14887 VDD108.n85 VDD108.t13 30.3459
R14888 VDD108.n263 VDD108.t33 29.9642
R14889 VDD108.n49 VDD108.t458 24.5101
R14890 VDD108.n47 VDD108.t463 24.5101
R14891 VDD108.n269 VDD108.t457 24.5101
R14892 VDD108.n264 VDD108.t462 24.5101
R14893 VDD108.n162 VDD108.t464 24.5101
R14894 VDD108.n82 VDD108.t455 24.5101
R14895 VDD108.n14 VDD108.t461 24.5101
R14896 VDD108.n15 VDD108.t456 24.5101
R14897 VDD108.n166 VDD108.t467 24.4392
R14898 VDD108.n86 VDD108.t466 24.4392
R14899 VDD108.n164 VDD108.n163 8.14079
R14900 VDD108.n84 VDD108.n83 8.14079
R14901 VDD108.n270 VDD108.n269 8.0005
R14902 VDD108.n167 VDD108.n166 8.0005
R14903 VDD108.n87 VDD108.n86 8.0005
R14904 VDD108.n465 VDD108.n464 7.02949
R14905 VDD108.n266 VDD108.n265 6.99025
R14906 VDD108.n52 VDD108.n46 6.3005
R14907 VDD108.n55 VDD108.n43 6.3005
R14908 VDD108.n58 VDD108.n40 6.3005
R14909 VDD108.n61 VDD108.n38 6.3005
R14910 VDD108.n207 VDD108.n206 6.3005
R14911 VDD108.n210 VDD108.n209 6.3005
R14912 VDD108.n383 VDD108.n382 6.3005
R14913 VDD108.n203 VDD108.n201 6.3005
R14914 VDD108.n200 VDD108.n199 6.3005
R14915 VDD108.n308 VDD108.n296 6.3005
R14916 VDD108.n317 VDD108.n289 6.3005
R14917 VDD108.n311 VDD108.n294 6.3005
R14918 VDD108.n306 VDD108.n299 6.3005
R14919 VDD108.n316 VDD108.n290 6.3005
R14920 VDD108.n353 VDD108.n352 6.3005
R14921 VDD108.n346 VDD108.n332 6.3005
R14922 VDD108.n350 VDD108.n349 6.3005
R14923 VDD108.n363 VDD108.n362 6.3005
R14924 VDD108.n359 VDD108.n329 6.3005
R14925 VDD108.n356 VDD108.n331 6.3005
R14926 VDD108.n365 VDD108.n364 6.3005
R14927 VDD108.n369 VDD108.n286 6.3005
R14928 VDD108.n283 VDD108.n252 6.3005
R14929 VDD108.n280 VDD108.n254 6.3005
R14930 VDD108.n277 VDD108.n257 6.3005
R14931 VDD108.n274 VDD108.n261 6.3005
R14932 VDD108.n237 VDD108.n219 6.3005
R14933 VDD108.n234 VDD108.n221 6.3005
R14934 VDD108.n231 VDD108.n224 6.3005
R14935 VDD108.n228 VDD108.n227 6.3005
R14936 VDD108.n242 VDD108.n241 6.3005
R14937 VDD108.n244 VDD108.n243 6.3005
R14938 VDD108.n249 VDD108.n248 6.3005
R14939 VDD108.n375 VDD108.n250 6.3005
R14940 VDD108.n385 VDD108.n384 6.3005
R14941 VDD108.n398 VDD108.n170 6.3005
R14942 VDD108.n395 VDD108.n174 6.3005
R14943 VDD108.n392 VDD108.n178 6.3005
R14944 VDD108.n389 VDD108.n180 6.3005
R14945 VDD108.n158 VDD108.n157 6.3005
R14946 VDD108.n151 VDD108.n137 6.3005
R14947 VDD108.n155 VDD108.n154 6.3005
R14948 VDD108.n403 VDD108.n402 6.3005
R14949 VDD108.n404 VDD108.n133 6.3005
R14950 VDD108.n405 VDD108.n129 6.3005
R14951 VDD108.n121 VDD108.n117 6.3005
R14952 VDD108.n125 VDD108.n113 6.3005
R14953 VDD108.n407 VDD108.n406 6.3005
R14954 VDD108.n105 VDD108.n104 6.3005
R14955 VDD108.n103 VDD108.n102 6.3005
R14956 VDD108.n96 VDD108.n95 6.3005
R14957 VDD108.n94 VDD108.n93 6.3005
R14958 VDD108.n414 VDD108.n74 6.3005
R14959 VDD108.n417 VDD108.n72 6.3005
R14960 VDD108.n420 VDD108.n70 6.3005
R14961 VDD108.n423 VDD108.n66 6.3005
R14962 VDD108.n441 VDD108.n440 6.3005
R14963 VDD108.n436 VDD108.n435 6.3005
R14964 VDD108.n434 VDD108.n433 6.3005
R14965 VDD108.n429 VDD108.n428 6.3005
R14966 VDD108.n19 VDD108.n13 6.3005
R14967 VDD108.n22 VDD108.n10 6.3005
R14968 VDD108.n25 VDD108.n7 6.3005
R14969 VDD108.n28 VDD108.n5 6.3005
R14970 VDD108.n447 VDD108.n446 6.3005
R14971 VDD108.n449 VDD108.n448 6.3005
R14972 VDD108.n457 VDD108.n456 6.3005
R14973 VDD108.n459 VDD108.n458 6.3005
R14974 VDD108.n30 VDD108.t417 5.85907
R14975 VDD108.n202 VDD108.t6 5.85907
R14976 VDD108.n461 VDD108.t314 5.85907
R14977 VDD108.n312 VDD108.n293 5.85007
R14978 VDD108.n304 VDD108.t230 5.22601
R14979 VDD108.n410 VDD108.n409 5.21771
R14980 VDD108.n334 VDD108.n333 5.213
R14981 VDD108.n228 VDD108.t22 5.213
R14982 VDD108.n139 VDD108.n138 5.213
R14983 VDD108.n368 VDD108.t54 5.18919
R14984 VDD108 VDD108.n195 5.16369
R14985 VDD108.n197 VDD108.n194 5.13761
R14986 VDD108.n439 VDD108.t12 5.13287
R14987 VDD108.n437 VDD108.t199 5.13287
R14988 VDD108.n34 VDD108.n33 5.13287
R14989 VDD108.n432 VDD108.t201 5.13287
R14990 VDD108.n431 VDD108.n35 5.13287
R14991 VDD108.n430 VDD108.t304 5.13287
R14992 VDD108.n427 VDD108.n36 5.13287
R14993 VDD108.n51 VDD108.t25 5.13287
R14994 VDD108.n54 VDD108.t56 5.13287
R14995 VDD108.n57 VDD108.t205 5.13287
R14996 VDD108.n59 VDD108.n39 5.13287
R14997 VDD108.n60 VDD108.t61 5.13287
R14998 VDD108.n62 VDD108.n37 5.13287
R14999 VDD108.n386 VDD108.t149 5.13287
R15000 VDD108.n186 VDD108.n185 5.13287
R15001 VDD108.n381 VDD108.t97 5.13287
R15002 VDD108.n380 VDD108.t75 5.13287
R15003 VDD108.n184 VDD108.n183 5.13287
R15004 VDD108.n187 VDD108.t167 5.13287
R15005 VDD108.n204 VDD108.n191 5.13287
R15006 VDD108.n370 VDD108.n285 5.13287
R15007 VDD108.n319 VDD108.n287 5.13287
R15008 VDD108.n315 VDD108.t80 5.13287
R15009 VDD108.n313 VDD108.n291 5.13287
R15010 VDD108.n310 VDD108.t366 5.13287
R15011 VDD108.n314 VDD108.t112 5.13287
R15012 VDD108.n318 VDD108.n288 5.13287
R15013 VDD108.n324 VDD108.n323 5.13287
R15014 VDD108.n354 VDD108.t368 5.13287
R15015 VDD108.n344 VDD108.n343 5.13287
R15016 VDD108.n345 VDD108.t69 5.13287
R15017 VDD108.n347 VDD108.n342 5.13287
R15018 VDD108.n339 VDD108.n335 5.13287
R15019 VDD108.n355 VDD108.t183 5.13287
R15020 VDD108.n357 VDD108.n330 5.13287
R15021 VDD108.n358 VDD108.t71 5.13287
R15022 VDD108.n360 VDD108.n328 5.13287
R15023 VDD108.n361 VDD108.t281 5.13287
R15024 VDD108.n327 VDD108.n326 5.13287
R15025 VDD108.n284 VDD108.n251 5.13287
R15026 VDD108.n282 VDD108.t154 5.13287
R15027 VDD108.n281 VDD108.n253 5.13287
R15028 VDD108.n279 VDD108.t84 5.13287
R15029 VDD108.n276 VDD108.t162 5.13287
R15030 VDD108.n238 VDD108.n218 5.13287
R15031 VDD108.n236 VDD108.t147 5.13287
R15032 VDD108.n235 VDD108.n220 5.13287
R15033 VDD108.n233 VDD108.t273 5.13287
R15034 VDD108.n230 VDD108.t302 5.13287
R15035 VDD108.n239 VDD108.n217 5.13287
R15036 VDD108.n240 VDD108.t192 5.13287
R15037 VDD108.n216 VDD108.n215 5.13287
R15038 VDD108.n245 VDD108.t190 5.13287
R15039 VDD108.n246 VDD108.n214 5.13287
R15040 VDD108.n247 VDD108.t359 5.13287
R15041 VDD108.n374 VDD108.t291 5.13287
R15042 VDD108.n388 VDD108.t110 5.13287
R15043 VDD108.n390 VDD108.n179 5.13287
R15044 VDD108.n391 VDD108.t73 5.13287
R15045 VDD108.n393 VDD108.n177 5.13287
R15046 VDD108.n396 VDD108.n173 5.13287
R15047 VDD108.n159 VDD108.t408 5.13287
R15048 VDD108.n149 VDD108.n148 5.13287
R15049 VDD108.n150 VDD108.t334 5.13287
R15050 VDD108.n152 VDD108.n147 5.13287
R15051 VDD108.n144 VDD108.n140 5.13287
R15052 VDD108.n401 VDD108.t403 5.13287
R15053 VDD108.n136 VDD108.n134 5.13287
R15054 VDD108.n135 VDD108.t332 5.13287
R15055 VDD108.n132 VDD108.n130 5.13287
R15056 VDD108.n131 VDD108.t316 5.13287
R15057 VDD108.n128 VDD108.n127 5.13287
R15058 VDD108.n124 VDD108.t223 5.13287
R15059 VDD108.n126 VDD108.n112 5.13287
R15060 VDD108.n106 VDD108.t218 5.13287
R15061 VDD108.n100 VDD108.n99 5.13287
R15062 VDD108.n101 VDD108.t243 5.13287
R15063 VDD108.n98 VDD108.n75 5.13287
R15064 VDD108.n79 VDD108.n78 5.13287
R15065 VDD108.n460 VDD108.t19 5.13287
R15066 VDD108.n455 VDD108.t175 5.13287
R15067 VDD108.n451 VDD108.n0 5.13287
R15068 VDD108.n450 VDD108.t259 5.13287
R15069 VDD108.n2 VDD108.n1 5.13287
R15070 VDD108.n445 VDD108.t241 5.13287
R15071 VDD108.n444 VDD108.n3 5.13287
R15072 VDD108.n18 VDD108.t32 5.13287
R15073 VDD108.n21 VDD108.t330 5.13287
R15074 VDD108.n24 VDD108.t252 5.13287
R15075 VDD108.n26 VDD108.n6 5.13287
R15076 VDD108.n27 VDD108.t250 5.13287
R15077 VDD108.n29 VDD108.n4 5.13287
R15078 VDD108.n413 VDD108.t122 5.12655
R15079 VDD108.n415 VDD108.n73 5.12655
R15080 VDD108.n416 VDD108.t245 5.12655
R15081 VDD108.n418 VDD108.n71 5.12655
R15082 VDD108.n419 VDD108.t139 5.12655
R15083 VDD108.n421 VDD108.n69 5.12655
R15084 VDD108.n424 VDD108.n65 5.12655
R15085 VDD108 VDD108.n463 5.11937
R15086 VDD108 VDD108.t102 5.11529
R15087 VDD108.n193 VDD108.t306 5.09407
R15088 VDD108.n302 VDD108.n300 5.09407
R15089 VDD108.n182 VDD108.n181 5.09407
R15090 VDD108.n372 VDD108.t89 5.09407
R15091 VDD108.n120 VDD108.n118 5.09407
R15092 VDD108.n123 VDD108.n114 5.09407
R15093 VDD108.n411 VDD108.n107 5.09407
R15094 VDD108.n425 VDD108.n63 5.09407
R15095 VDD108.n400 VDD108.n399 5.08521
R15096 VDD108.n378 VDD108.n377 4.99361
R15097 VDD108.n273 VDD108.t35 4.8755
R15098 VDD108.n169 VDD108.n160 4.8755
R15099 VDD108.n89 VDD108.n80 4.8755
R15100 VDD108.n266 VDD108.n262 4.51272
R15101 VDD108.n269 VDD108.n268 4.5005
R15102 VDD108 VDD108.n14 4.35564
R15103 VDD108.n205 VDD108.t1 4.12326
R15104 VDD108.n309 VDD108.n295 4.12326
R15105 VDD108.n122 VDD108.n116 4.12326
R15106 VDD108 VDD108.n49 4.09565
R15107 VDD108.n48 VDD108.n47 4.08504
R15108 VDD108 VDD108.n15 4.00785
R15109 VDD108 VDD108.n465 3.85641
R15110 VDD108.n267 VDD108.n263 3.6022
R15111 VDD108.n17 VDD108 3.06902
R15112 VDD108.n50 VDD108.n48 2.93012
R15113 VDD108.n17 VDD108.n16 2.86671
R15114 VDD108.n438 VDD108.n32 2.85787
R15115 VDD108.n53 VDD108.n45 2.85787
R15116 VDD108.n56 VDD108.n42 2.85787
R15117 VDD108.n190 VDD108.n189 2.85787
R15118 VDD108.n307 VDD108.n298 2.85787
R15119 VDD108.n348 VDD108.n341 2.85787
R15120 VDD108.n338 VDD108.n337 2.85787
R15121 VDD108.n322 VDD108.n321 2.85787
R15122 VDD108.n278 VDD108.n256 2.85787
R15123 VDD108.n275 VDD108.n259 2.85787
R15124 VDD108.n232 VDD108.n223 2.85787
R15125 VDD108.n229 VDD108.n226 2.85787
R15126 VDD108.n213 VDD108.n212 2.85787
R15127 VDD108.n394 VDD108.n176 2.85787
R15128 VDD108.n397 VDD108.n172 2.85787
R15129 VDD108.n153 VDD108.n146 2.85787
R15130 VDD108.n143 VDD108.n142 2.85787
R15131 VDD108.n111 VDD108.n110 2.85787
R15132 VDD108.n97 VDD108.n77 2.85787
R15133 VDD108.n92 VDD108.n91 2.85787
R15134 VDD108.n454 VDD108.n453 2.85787
R15135 VDD108.n20 VDD108.n12 2.85787
R15136 VDD108.n23 VDD108.n9 2.85787
R15137 VDD108.n422 VDD108.n68 2.85155
R15138 VDD108.n50 VDD108 2.83528
R15139 VDD108.n18 VDD108.n17 2.28244
R15140 VDD108.n32 VDD108.t197 2.2755
R15141 VDD108.n32 VDD108.n31 2.2755
R15142 VDD108.n45 VDD108.t213 2.2755
R15143 VDD108.n45 VDD108.n44 2.2755
R15144 VDD108.n42 VDD108.t203 2.2755
R15145 VDD108.n42 VDD108.n41 2.2755
R15146 VDD108.n189 VDD108.t382 2.2755
R15147 VDD108.n189 VDD108.n188 2.2755
R15148 VDD108.n298 VDD108.t364 2.2755
R15149 VDD108.n298 VDD108.n297 2.2755
R15150 VDD108.n341 VDD108.t348 2.2755
R15151 VDD108.n341 VDD108.n340 2.2755
R15152 VDD108.n337 VDD108.t377 2.2755
R15153 VDD108.n337 VDD108.n336 2.2755
R15154 VDD108.n321 VDD108.t392 2.2755
R15155 VDD108.n321 VDD108.n320 2.2755
R15156 VDD108.n256 VDD108.t82 2.2755
R15157 VDD108.n256 VDD108.n255 2.2755
R15158 VDD108.n259 VDD108.t289 2.2755
R15159 VDD108.n259 VDD108.n258 2.2755
R15160 VDD108.n223 VDD108.t188 2.2755
R15161 VDD108.n223 VDD108.n222 2.2755
R15162 VDD108.n226 VDD108.t63 2.2755
R15163 VDD108.n226 VDD108.n225 2.2755
R15164 VDD108.n212 VDD108.t228 2.2755
R15165 VDD108.n212 VDD108.n211 2.2755
R15166 VDD108.n176 VDD108.t355 2.2755
R15167 VDD108.n176 VDD108.n175 2.2755
R15168 VDD108.n172 VDD108.t387 2.2755
R15169 VDD108.n172 VDD108.n171 2.2755
R15170 VDD108.n146 VDD108.t357 2.2755
R15171 VDD108.n146 VDD108.n145 2.2755
R15172 VDD108.n142 VDD108.t445 2.2755
R15173 VDD108.n142 VDD108.n141 2.2755
R15174 VDD108.n110 VDD108.t438 2.2755
R15175 VDD108.n110 VDD108.n109 2.2755
R15176 VDD108.n77 VDD108.t353 2.2755
R15177 VDD108.n77 VDD108.n76 2.2755
R15178 VDD108.n91 VDD108.t443 2.2755
R15179 VDD108.n91 VDD108.n90 2.2755
R15180 VDD108.n68 VDD108.t453 2.2755
R15181 VDD108.n68 VDD108.n67 2.2755
R15182 VDD108.n453 VDD108.t427 2.2755
R15183 VDD108.n453 VDD108.n452 2.2755
R15184 VDD108.n12 VDD108.t425 2.2755
R15185 VDD108.n12 VDD108.n11 2.2755
R15186 VDD108.n9 VDD108.t257 2.2755
R15187 VDD108.n9 VDD108.n8 2.2755
R15188 VDD108.n51 VDD108.n50 2.27489
R15189 VDD108.n163 VDD108.n162 2.11346
R15190 VDD108.n83 VDD108.n82 2.11346
R15191 VDD108.n265 VDD108.n264 2.11318
R15192 VDD108.n165 VDD108.n164 1.81921
R15193 VDD108.n85 VDD108.n84 1.81921
R15194 VDD108.n426 VDD108.n425 1.78842
R15195 VDD108.n197 VDD108 1.77385
R15196 VDD108 VDD108.n324 1.77343
R15197 VDD108.n268 VDD108.n266 1.54696
R15198 VDD108.n239 VDD108.n238 1.16167
R15199 VDD108.n355 VDD108.n354 1.16051
R15200 VDD108.n401 VDD108.n400 1.12915
R15201 VDD108.n388 VDD108.n387 1.0737
R15202 VDD108.n426 VDD108.n62 1.02928
R15203 VDD108.n443 VDD108.n29 1.02928
R15204 VDD108.n371 VDD108.n284 1.01882
R15205 VDD108.n412 VDD108.n106 1.01824
R15206 VDD108.n269 VDD108.n263 0.798596
R15207 VDD108.n378 VDD108 0.59265
R15208 VDD108 VDD108.n366 0.468962
R15209 VDD108.n408 VDD108 0.468962
R15210 VDD108.n166 VDD108.n165 0.423118
R15211 VDD108.n86 VDD108.n85 0.423118
R15212 VDD108.n121 VDD108.n120 0.389068
R15213 VDD108.n379 VDD108.n378 0.346452
R15214 VDD108.n274 VDD108.n273 0.337997
R15215 VDD108.n93 VDD108.n89 0.337997
R15216 VDD108.n273 VDD108.n272 0.328132
R15217 VDD108.n169 VDD108.n168 0.328132
R15218 VDD108.n89 VDD108.n88 0.328132
R15219 VDD108 VDD108.n376 0.316077
R15220 VDD108 VDD108.n126 0.274338
R15221 VDD108 VDD108.n122 0.269908
R15222 VDD108.n399 VDD108.n169 0.257868
R15223 VDD108.n57 VDD108.n56 0.233919
R15224 VDD108.n54 VDD108.n53 0.233919
R15225 VDD108.n339 VDD108.n338 0.233919
R15226 VDD108.n348 VDD108.n347 0.233919
R15227 VDD108.n279 VDD108.n278 0.233919
R15228 VDD108.n276 VDD108.n275 0.233919
R15229 VDD108.n233 VDD108.n232 0.233919
R15230 VDD108.n230 VDD108.n229 0.233919
R15231 VDD108.n397 VDD108.n396 0.233919
R15232 VDD108.n394 VDD108.n393 0.233919
R15233 VDD108.n144 VDD108.n143 0.233919
R15234 VDD108.n153 VDD108.n152 0.233919
R15235 VDD108.n92 VDD108.n79 0.233919
R15236 VDD108.n98 VDD108.n97 0.233919
R15237 VDD108.n24 VDD108.n23 0.233919
R15238 VDD108.n21 VDD108.n20 0.233919
R15239 VDD108.n367 VDD108 0.216814
R15240 VDD108.n379 VDD108 0.216814
R15241 VDD108.n124 VDD108.n123 0.170499
R15242 VDD108 VDD108.n424 0.166121
R15243 VDD108.n465 VDD108 0.156451
R15244 VDD108.n387 VDD108.n386 0.14292
R15245 VDD108.n60 VDD108.n59 0.141016
R15246 VDD108.n345 VDD108.n344 0.141016
R15247 VDD108.n361 VDD108.n360 0.141016
R15248 VDD108.n358 VDD108.n357 0.141016
R15249 VDD108.n282 VDD108.n281 0.141016
R15250 VDD108.n236 VDD108.n235 0.141016
R15251 VDD108.n240 VDD108.n216 0.141016
R15252 VDD108.n246 VDD108.n245 0.141016
R15253 VDD108.n391 VDD108.n390 0.141016
R15254 VDD108.n150 VDD108.n149 0.141016
R15255 VDD108.n132 VDD108.n131 0.141016
R15256 VDD108.n136 VDD108.n135 0.141016
R15257 VDD108.n101 VDD108.n100 0.141016
R15258 VDD108.n27 VDD108.n26 0.141016
R15259 VDD108 VDD108.n410 0.140259
R15260 VDD108.n387 VDD108.n182 0.139745
R15261 VDD108.n305 VDD108.n302 0.137219
R15262 VDD108.n198 VDD108.n193 0.13637
R15263 VDD108.n419 VDD108.n418 0.125672
R15264 VDD108.n416 VDD108.n415 0.125672
R15265 VDD108.n327 VDD108 0.123016
R15266 VDD108.n128 VDD108 0.123016
R15267 VDD108.n247 VDD108 0.122435
R15268 VDD108.n413 VDD108.n412 0.117172
R15269 VDD108 VDD108.n213 0.111984
R15270 VDD108 VDD108.n322 0.111403
R15271 VDD108 VDD108.n111 0.111403
R15272 VDD108 VDD108.n421 0.109638
R15273 VDD108.n122 VDD108 0.109408
R15274 VDD108.n163 VDD108 0.107393
R15275 VDD108.n83 VDD108 0.107393
R15276 VDD108.n62 VDD108.n61 0.107339
R15277 VDD108.n59 VDD108.n58 0.107339
R15278 VDD108.n346 VDD108.n345 0.107339
R15279 VDD108.n354 VDD108.n353 0.107339
R15280 VDD108.n362 VDD108.n361 0.107339
R15281 VDD108.n359 VDD108.n358 0.107339
R15282 VDD108.n356 VDD108.n355 0.107339
R15283 VDD108.n284 VDD108.n283 0.107339
R15284 VDD108.n281 VDD108.n280 0.107339
R15285 VDD108.n238 VDD108.n237 0.107339
R15286 VDD108.n235 VDD108.n234 0.107339
R15287 VDD108.n241 VDD108.n239 0.107339
R15288 VDD108.n244 VDD108.n216 0.107339
R15289 VDD108.n248 VDD108.n246 0.107339
R15290 VDD108.n386 VDD108.n385 0.107339
R15291 VDD108.n392 VDD108.n391 0.107339
R15292 VDD108.n389 VDD108.n388 0.107339
R15293 VDD108.n151 VDD108.n150 0.107339
R15294 VDD108.n159 VDD108.n158 0.107339
R15295 VDD108.n131 VDD108.n129 0.107339
R15296 VDD108.n135 VDD108.n133 0.107339
R15297 VDD108.n402 VDD108.n401 0.107339
R15298 VDD108.n125 VDD108.n124 0.107339
R15299 VDD108.n102 VDD108.n101 0.107339
R15300 VDD108.n106 VDD108.n105 0.107339
R15301 VDD108.n29 VDD108.n28 0.107339
R15302 VDD108.n26 VDD108.n25 0.107339
R15303 VDD108.n265 VDD108 0.106795
R15304 VDD108.n338 VDD108 0.106758
R15305 VDD108 VDD108.n348 0.106758
R15306 VDD108 VDD108.n397 0.106758
R15307 VDD108 VDD108.n394 0.106758
R15308 VDD108.n143 VDD108 0.106758
R15309 VDD108 VDD108.n153 0.106758
R15310 VDD108 VDD108.n92 0.106758
R15311 VDD108.n97 VDD108 0.106758
R15312 VDD108.n56 VDD108 0.106177
R15313 VDD108.n53 VDD108 0.106177
R15314 VDD108.n278 VDD108 0.106177
R15315 VDD108.n275 VDD108 0.106177
R15316 VDD108.n232 VDD108 0.106177
R15317 VDD108.n229 VDD108 0.106177
R15318 VDD108.n23 VDD108 0.106177
R15319 VDD108.n20 VDD108 0.106177
R15320 VDD108.n412 VDD108.n411 0.104
R15321 VDD108.n422 VDD108 0.0992931
R15322 VDD108.n420 VDD108.n419 0.0956724
R15323 VDD108.n417 VDD108.n416 0.0956724
R15324 VDD108.n414 VDD108.n413 0.0956724
R15325 VDD108 VDD108.n422 0.0951552
R15326 VDD108.n374 VDD108 0.0847644
R15327 VDD108.n55 VDD108.n54 0.080629
R15328 VDD108.n52 VDD108.n51 0.080629
R15329 VDD108.n349 VDD108.n339 0.080629
R15330 VDD108.n277 VDD108.n276 0.080629
R15331 VDD108.n231 VDD108.n230 0.080629
R15332 VDD108.n399 VDD108.n398 0.080629
R15333 VDD108.n396 VDD108.n395 0.080629
R15334 VDD108.n154 VDD108.n144 0.080629
R15335 VDD108.n96 VDD108.n79 0.080629
R15336 VDD108.n22 VDD108.n21 0.080629
R15337 VDD108.n19 VDD108.n18 0.080629
R15338 VDD108 VDD108.n60 0.0794677
R15339 VDD108 VDD108.n57 0.0794677
R15340 VDD108 VDD108.n282 0.0794677
R15341 VDD108 VDD108.n279 0.0794677
R15342 VDD108 VDD108.n236 0.0794677
R15343 VDD108 VDD108.n233 0.0794677
R15344 VDD108 VDD108.n240 0.0794677
R15345 VDD108.n245 VDD108 0.0794677
R15346 VDD108 VDD108.n247 0.0794677
R15347 VDD108 VDD108.n27 0.0794677
R15348 VDD108 VDD108.n24 0.0794677
R15349 VDD108.n347 VDD108 0.0788871
R15350 VDD108.n344 VDD108 0.0788871
R15351 VDD108 VDD108.n327 0.0788871
R15352 VDD108.n360 VDD108 0.0788871
R15353 VDD108.n357 VDD108 0.0788871
R15354 VDD108.n393 VDD108 0.0788871
R15355 VDD108.n390 VDD108 0.0788871
R15356 VDD108.n152 VDD108 0.0788871
R15357 VDD108.n149 VDD108 0.0788871
R15358 VDD108 VDD108.n128 0.0788871
R15359 VDD108 VDD108.n132 0.0788871
R15360 VDD108 VDD108.n136 0.0788871
R15361 VDD108 VDD108.n98 0.0788871
R15362 VDD108.n100 VDD108 0.0788871
R15363 VDD108.n126 VDD108 0.0754032
R15364 VDD108.n161 VDD108 0.0733571
R15365 VDD108.n81 VDD108 0.0733571
R15366 VDD108.n424 VDD108.n423 0.0718793
R15367 VDD108.n193 VDD108 0.0709717
R15368 VDD108.n421 VDD108 0.0703276
R15369 VDD108.n418 VDD108 0.0703276
R15370 VDD108.n415 VDD108 0.0703276
R15371 VDD108.n302 VDD108 0.0701226
R15372 VDD108 VDD108.n182 0.0701226
R15373 VDD108.n120 VDD108 0.0701226
R15374 VDD108.n123 VDD108 0.0701226
R15375 VDD108.n271 VDD108 0.0690714
R15376 VDD108.n376 VDD108.n213 0.0616715
R15377 VDD108.n371 VDD108.n370 0.0601785
R15378 VDD108.n366 VDD108.n324 0.0556613
R15379 VDD108.n304 VDD108 0.0531999
R15380 VDD108.n372 VDD108.n371 0.0531705
R15381 VDD108.n370 VDD108.n369 0.0489211
R15382 VDD108.n272 VDD108.n271 0.0471071
R15383 VDD108.n168 VDD108.n161 0.0471071
R15384 VDD108.n88 VDD108.n81 0.0471071
R15385 VDD108.n366 VDD108.n322 0.0417258
R15386 VDD108.n408 VDD108.n111 0.0417258
R15387 VDD108.n410 VDD108.n408 0.0417109
R15388 VDD108.n411 VDD108 0.0415
R15389 VDD108.n425 VDD108 0.0415
R15390 VDD108.n167 VDD108.n164 0.0387491
R15391 VDD108.n87 VDD108.n84 0.0387491
R15392 VDD108.n439 VDD108.n30 0.037789
R15393 VDD108.n461 VDD108.n460 0.0376465
R15394 VDD108.n375 VDD108.n374 0.0368158
R15395 VDD108 VDD108.n190 0.0366978
R15396 VDD108.n307 VDD108 0.0365
R15397 VDD108.n270 VDD108.n262 0.0358571
R15398 VDD108.n168 VDD108.n167 0.0358571
R15399 VDD108.n88 VDD108.n87 0.0358571
R15400 VDD108.n205 VDD108.n204 0.0349176
R15401 VDD108.n310 VDD108.n309 0.0349176
R15402 VDD108.n272 VDD108.n270 0.03425
R15403 VDD108 VDD108.n187 0.033533
R15404 VDD108.n313 VDD108 0.0333352
R15405 VDD108 VDD108.n368 0.033241
R15406 VDD108.n400 VDD108.n159 0.0318548
R15407 VDD108.n187 VDD108.n186 0.0307637
R15408 VDD108.n314 VDD108.n313 0.0307637
R15409 VDD108.n431 VDD108.n430 0.0283517
R15410 VDD108.n432 VDD108.n34 0.0283517
R15411 VDD108.n445 VDD108.n2 0.0282452
R15412 VDD108.n451 VDD108.n450 0.0282452
R15413 VDD108 VDD108.n310 0.0274011
R15414 VDD108.n204 VDD108 0.0272033
R15415 VDD108.n427 VDD108.n426 0.0267404
R15416 VDD108.n444 VDD108.n443 0.0266401
R15417 VDD108.n368 VDD108.n367 0.0252441
R15418 VDD108 VDD108.n437 0.0246688
R15419 VDD108.n455 VDD108 0.0245764
R15420 VDD108.n198 VDD108.n197 0.0230424
R15421 VDD108.n438 VDD108 0.0225972
R15422 VDD108 VDD108.n454 0.0225127
R15423 VDD108 VDD108.n372 0.0217216
R15424 VDD108.n429 VDD108.n427 0.0216765
R15425 VDD108.n433 VDD108.n431 0.0216765
R15426 VDD108.n436 VDD108.n34 0.0216765
R15427 VDD108.n446 VDD108.n444 0.0215955
R15428 VDD108.n449 VDD108.n2 0.0215955
R15429 VDD108.n456 VDD108.n451 0.0215955
R15430 VDD108 VDD108.n438 0.0214463
R15431 VDD108.n454 VDD108 0.0213662
R15432 VDD108.n366 VDD108.n365 0.0201154
R15433 VDD108.n408 VDD108.n407 0.0201154
R15434 VDD108.n210 VDD108.n184 0.0192912
R15435 VDD108.n382 VDD108.n381 0.0192912
R15436 VDD108.n318 VDD108.n317 0.0192912
R15437 VDD108.n316 VDD108.n315 0.0192912
R15438 VDD108.n186 VDD108.n184 0.0181044
R15439 VDD108.n381 VDD108.n380 0.0181044
R15440 VDD108.n319 VDD108.n318 0.0181044
R15441 VDD108.n315 VDD108.n314 0.0181044
R15442 VDD108.n440 VDD108.n439 0.0163824
R15443 VDD108.n460 VDD108.n459 0.0163217
R15444 VDD108.n430 VDD108 0.0161522
R15445 VDD108 VDD108.n432 0.0161522
R15446 VDD108.n437 VDD108 0.0161522
R15447 VDD108 VDD108.n445 0.0160924
R15448 VDD108.n450 VDD108 0.0160924
R15449 VDD108 VDD108.n455 0.0160924
R15450 VDD108.n308 VDD108.n307 0.0157308
R15451 VDD108.n206 VDD108.n190 0.015533
R15452 VDD108.n199 VDD108.n198 0.0149396
R15453 VDD108.n306 VDD108.n305 0.0147418
R15454 VDD108.n16 VDD108 0.0113333
R15455 VDD108.n376 VDD108 0.00944737
R15456 VDD108.n271 VDD108 0.00907143
R15457 VDD108.n305 VDD108.n304 0.00906907
R15458 VDD108 VDD108.n205 0.00781868
R15459 VDD108.n367 VDD108.n319 0.00762088
R15460 VDD108.n309 VDD108 0.00762088
R15461 VDD108.n380 VDD108.n379 0.00742308
R15462 VDD108 VDD108.n121 0.00579412
R15463 VDD108 VDD108.n125 0.00572581
R15464 VDD108.n48 VDD108 0.00564286
R15465 VDD108.n443 VDD108 0.00508599
R15466 VDD108.n161 VDD108 0.00478571
R15467 VDD108.n81 VDD108 0.00478571
R15468 VDD108.n16 VDD108 0.00466667
R15469 VDD108.n267 VDD108.n262 0.00371429
R15470 VDD108.n312 VDD108.n311 0.00366484
R15471 VDD108.n203 VDD108.n202 0.00346703
R15472 VDD108 VDD108.n316 0.00228022
R15473 VDD108 VDD108.n346 0.00224194
R15474 VDD108.n353 VDD108 0.00224194
R15475 VDD108.n362 VDD108 0.00224194
R15476 VDD108 VDD108.n359 0.00224194
R15477 VDD108 VDD108.n356 0.00224194
R15478 VDD108.n385 VDD108 0.00224194
R15479 VDD108 VDD108.n392 0.00224194
R15480 VDD108 VDD108.n389 0.00224194
R15481 VDD108 VDD108.n151 0.00224194
R15482 VDD108.n158 VDD108 0.00224194
R15483 VDD108.n129 VDD108 0.00224194
R15484 VDD108.n133 VDD108 0.00224194
R15485 VDD108.n402 VDD108 0.00224194
R15486 VDD108.n102 VDD108 0.00224194
R15487 VDD108.n105 VDD108 0.00224194
R15488 VDD108.n268 VDD108.n267 0.00210714
R15489 VDD108 VDD108.n210 0.00208242
R15490 VDD108 VDD108.n420 0.00205172
R15491 VDD108 VDD108.n417 0.00205172
R15492 VDD108 VDD108.n414 0.00205172
R15493 VDD108.n206 VDD108 0.00188462
R15494 VDD108 VDD108.n308 0.00188462
R15495 VDD108.n61 VDD108 0.00166129
R15496 VDD108.n58 VDD108 0.00166129
R15497 VDD108 VDD108.n55 0.00166129
R15498 VDD108 VDD108.n52 0.00166129
R15499 VDD108.n283 VDD108 0.00166129
R15500 VDD108.n280 VDD108 0.00166129
R15501 VDD108 VDD108.n277 0.00166129
R15502 VDD108 VDD108.n274 0.00166129
R15503 VDD108.n237 VDD108 0.00166129
R15504 VDD108.n234 VDD108 0.00166129
R15505 VDD108 VDD108.n231 0.00166129
R15506 VDD108 VDD108.n228 0.00166129
R15507 VDD108.n241 VDD108 0.00166129
R15508 VDD108 VDD108.n244 0.00166129
R15509 VDD108.n248 VDD108 0.00166129
R15510 VDD108.n28 VDD108 0.00166129
R15511 VDD108.n25 VDD108 0.00166129
R15512 VDD108 VDD108.n22 0.00166129
R15513 VDD108 VDD108.n19 0.00166129
R15514 VDD108 VDD108.n203 0.00109341
R15515 VDD108.n382 VDD108 0.00109341
R15516 VDD108 VDD108.n334 0.00108064
R15517 VDD108.n349 VDD108 0.00108064
R15518 VDD108.n398 VDD108 0.00108064
R15519 VDD108.n395 VDD108 0.00108064
R15520 VDD108 VDD108.n139 0.00108064
R15521 VDD108.n154 VDD108 0.00108064
R15522 VDD108.n93 VDD108 0.00108064
R15523 VDD108 VDD108.n96 0.00108064
R15524 VDD108.n365 VDD108 0.00107692
R15525 VDD108.n407 VDD108 0.00107692
R15526 VDD108.n369 VDD108 0.00102632
R15527 VDD108 VDD108.n375 0.00102632
R15528 VDD108.n423 VDD108 0.00101724
R15529 VDD108.n202 VDD108 0.000895604
R15530 VDD108.n317 VDD108 0.000895604
R15531 VDD108 VDD108.n312 0.000895604
R15532 VDD108.n311 VDD108 0.000895604
R15533 VDD108 VDD108.n306 0.000895604
R15534 VDD108 VDD108.n429 0.000730179
R15535 VDD108.n433 VDD108 0.000730179
R15536 VDD108 VDD108.n436 0.000730179
R15537 VDD108.n440 VDD108 0.000730179
R15538 VDD108 VDD108.n30 0.000730179
R15539 VDD108.n446 VDD108 0.000729299
R15540 VDD108 VDD108.n449 0.000729299
R15541 VDD108.n456 VDD108 0.000729299
R15542 VDD108.n459 VDD108 0.000729299
R15543 VDD108 VDD108.n461 0.000729299
R15544 VDD108.n199 VDD108 0.000697802
R15545 VDD105.n388 VDD105.n49 190685
R15546 VDD105.n388 VDD105.t473 83097.6
R15547 VDD105.n285 VDD105.t302 29077.7
R15548 VDD105.n353 VDD105.n352 11185.2
R15549 VDD105.n312 VDD105.n311 11185.2
R15550 VDD105.t111 VDD105.n43 1105.93
R15551 VDD105.n289 VDD105.t195 1105.93
R15552 VDD105.t167 VDD105.t173 961.905
R15553 VDD105.t435 VDD105.t333 961.905
R15554 VDD105.t335 VDD105.t9 961.905
R15555 VDD105.t184 VDD105.t221 961.905
R15556 VDD105.t356 VDD105.t15 961.905
R15557 VDD105.t407 VDD105.t83 961.905
R15558 VDD105.t159 VDD105.t215 765.152
R15559 VDD105.t464 VDD105.t25 765.152
R15560 VDD105.t77 VDD105.t33 765.152
R15561 VDD105.t320 VDD105.t200 765.152
R15562 VDD105.t328 VDD105.t351 765.152
R15563 VDD105.t300 VDD105.t188 765.152
R15564 VDD105.t203 VDD105.t206 765.152
R15565 VDD105.t349 VDD105.t331 765.152
R15566 VDD105.t368 VDD105.t277 765.152
R15567 VDD105.t353 VDD105.t106 765.152
R15568 VDD105.t120 VDD105.t23 765.152
R15569 VDD105.t377 VDD105.t13 765.152
R15570 VDD105.t177 VDD105.t359 765.152
R15571 VDD105.t268 VDD105.t128 765.152
R15572 VDD105.t271 VDD105.t372 765.152
R15573 VDD105.t279 VDD105.t249 765.152
R15574 VDD105.t312 VDD105.t260 765.152
R15575 VDD105.t315 VDD105.t116 765.152
R15576 VDD105.t153 VDD105.t101 765.152
R15577 VDD105.t298 VDD105.t292 765.152
R15578 VDD105.t17 VDD105.t223 765.152
R15579 VDD105.t325 VDD105.t237 765.152
R15580 VDD105.t309 VDD105.t257 765.152
R15581 VDD105.t254 VDD105.t114 765.152
R15582 VDD105.t274 VDD105.t452 765.152
R15583 VDD105.t265 VDD105.t125 765.152
R15584 VDD105.t122 VDD105.t370 765.152
R15585 VDD105.t338 VDD105.t341 765.152
R15586 VDD105.t182 VDD105.t7 765.152
R15587 VDD105.t141 VDD105.t208 765.152
R15588 VDD105.t170 VDD105.t230 765.152
R15589 VDD105.t284 VDD105.t162 765.152
R15590 VDD105.t426 VDD105.t186 765.152
R15591 VDD105.t262 VDD105.t89 765.152
R15592 VDD105.t289 VDD105.t295 765.152
R15593 VDD105.t227 VDD105.t225 765.152
R15594 VDD105.t197 VDD105.t343 765.152
R15595 VDD105.t28 VDD105.t466 765.152
R15596 VDD105.t409 VDD105.t31 765.152
R15597 VDD105.n352 VDD105.t180 676.191
R15598 VDD105.n311 VDD105.t118 676.191
R15599 VDD105.t164 VDD105.n49 669.048
R15600 VDD105.t85 VDD105.t318 645.307
R15601 VDD105.t108 VDD105.t150 642.843
R15602 VDD105.n388 VDD105.n45 525.424
R15603 VDD105.n286 VDD105.n285 525.424
R15604 VDD105.n353 VDD105.t193 485.714
R15605 VDD105.n312 VDD105.t57 485.714
R15606 VDD105 VDD105.n140 429.187
R15607 VDD105 VDD105.n295 427.092
R15608 VDD105.n301 VDD105 427.092
R15609 VDD105 VDD105.n201 426.699
R15610 VDD105 VDD105.n213 426.699
R15611 VDD105 VDD105.n433 426.699
R15612 VDD105.t428 VDD105.n353 426.44
R15613 VDD105.t148 VDD105.n312 426.44
R15614 VDD105 VDD105.n290 425.019
R15615 VDD105 VDD105.n34 424.618
R15616 VDD105 VDD105.n38 424.618
R15617 VDD105 VDD105.n42 422.557
R15618 VDD105.n433 VDD105.t156 386.365
R15619 VDD105.t92 VDD105.n34 386.365
R15620 VDD105.t460 VDD105.n38 386.365
R15621 VDD105.n140 VDD105.t2 386.365
R15622 VDD105.n301 VDD105.t379 386.365
R15623 VDD105.n295 VDD105.t433 386.365
R15624 VDD105.t210 VDD105.n201 386.365
R15625 VDD105.n213 VDD105.t60 386.365
R15626 VDD105.t473 VDD105.t435 380.952
R15627 VDD105.t221 VDD105.t420 380.952
R15628 VDD105.t83 VDD105.t143 380.952
R15629 VDD105.n34 VDD105.t95 378.788
R15630 VDD105.n38 VDD105.t232 378.788
R15631 VDD105.n42 VDD105.t99 378.788
R15632 VDD105.t381 VDD105.n301 378.788
R15633 VDD105.n295 VDD105.t135 378.788
R15634 VDD105.n290 VDD105.t384 378.788
R15635 VDD105.t215 VDD105.t458 303.031
R15636 VDD105.t188 VDD105.t430 303.031
R15637 VDD105.t392 VDD105.t349 303.031
R15638 VDD105.t414 VDD105.t368 303.031
R15639 VDD105.t387 VDD105.t120 303.031
R15640 VDD105.t132 VDD105.t377 303.031
R15641 VDD105.t302 VDD105.t177 303.031
R15642 VDD105.t249 VDD105.t448 303.031
R15643 VDD105.t101 VDD105.t242 303.031
R15644 VDD105.t237 VDD105.t450 303.031
R15645 VDD105.t395 VDD105.t309 303.031
R15646 VDD105.t452 VDD105.t307 303.031
R15647 VDD105.t397 VDD105.t265 303.031
R15648 VDD105.t402 VDD105.t182 303.031
R15649 VDD105.t423 VDD105.t141 303.031
R15650 VDD105.t399 VDD105.t284 303.031
R15651 VDD105.t470 VDD105.t426 303.031
R15652 VDD105.t89 VDD105.t247 303.031
R15653 VDD105.t390 VDD105.t289 303.031
R15654 VDD105.t343 VDD105.t444 303.031
R15655 VDD105.t405 VDD105.t28 303.031
R15656 VDD105.t282 VDD105.n49 292.858
R15657 VDD105.n352 VDD105.t4 285.714
R15658 VDD105.n311 VDD105.t20 285.714
R15659 VDD105.n380 VDD105.t437 242.857
R15660 VDD105.n381 VDD105.t167 242.857
R15661 VDD105.n387 VDD105.t164 242.857
R15662 VDD105.n339 VDD105.t218 242.857
R15663 VDD105.n340 VDD105.t335 242.857
R15664 VDD105.t4 VDD105.n351 242.857
R15665 VDD105.t420 VDD105.n350 242.857
R15666 VDD105.n167 VDD105.t80 242.857
R15667 VDD105.n168 VDD105.t356 242.857
R15668 VDD105.t20 VDD105.n310 242.857
R15669 VDD105.t143 VDD105.n309 242.857
R15670 VDD105.n127 VDD105.t190 193.183
R15671 VDD105.n133 VDD105.t200 193.183
R15672 VDD105.n134 VDD105.t328 193.183
R15673 VDD105.n139 VDD105.t430 193.183
R15674 VDD105.n72 VDD105.t365 193.183
R15675 VDD105.n74 VDD105.t203 193.183
R15676 VDD105.n77 VDD105.t392 193.183
R15677 VDD105.n80 VDD105.t414 193.183
R15678 VDD105.n143 VDD105.t374 193.183
R15679 VDD105.n145 VDD105.t353 193.183
R15680 VDD105.n148 VDD105.t387 193.183
R15681 VDD105.n151 VDD105.t132 193.183
R15682 VDD105.n302 VDD105.t381 193.183
R15683 VDD105.n300 VDD105.t135 193.183
R15684 VDD105.n294 VDD105.t384 193.183
R15685 VDD105.n315 VDD105.t138 193.183
R15686 VDD105.n317 VDD105.t338 193.183
R15687 VDD105.n320 VDD105.t402 193.183
R15688 VDD105.n323 VDD105.t423 193.183
R15689 VDD105.n356 VDD105.t417 193.183
R15690 VDD105.n358 VDD105.t170 193.183
R15691 VDD105.n361 VDD105.t399 193.183
R15692 VDD105.n364 VDD105.t470 193.183
R15693 VDD105.t458 VDD105.n441 191.288
R15694 VDD105.n442 VDD105.t464 191.288
R15695 VDD105.t33 VDD105.n450 191.288
R15696 VDD105.n451 VDD105.t213 191.288
R15697 VDD105.t95 VDD105.n32 191.288
R15698 VDD105.t232 VDD105.n36 191.288
R15699 VDD105.t99 VDD105.n40 191.288
R15700 VDD105.n284 VDD105.t128 191.288
R15701 VDD105.t372 VDD105.n197 191.288
R15702 VDD105.n199 VDD105.t175 191.288
R15703 VDD105.t448 VDD105.n203 191.288
R15704 VDD105.t260 VDD105.n207 191.288
R15705 VDD105.t116 VDD105.n209 191.288
R15706 VDD105.n211 VDD105.t252 191.288
R15707 VDD105.t242 VDD105.n418 191.288
R15708 VDD105.n419 VDD105.t298 191.288
R15709 VDD105.t223 VDD105.n427 191.288
R15710 VDD105.n428 VDD105.t104 191.288
R15711 VDD105.t450 VDD105.n225 191.288
R15712 VDD105.n226 VDD105.t395 191.288
R15713 VDD105.t114 VDD105.n234 191.288
R15714 VDD105.n235 VDD105.t240 191.288
R15715 VDD105.t307 VDD105.n262 191.288
R15716 VDD105.n263 VDD105.t397 191.288
R15717 VDD105.t370 VDD105.n271 191.288
R15718 VDD105.n272 VDD105.t446 191.288
R15719 VDD105.t247 VDD105.n13 191.288
R15720 VDD105.n14 VDD105.t390 191.288
R15721 VDD105.t225 VDD105.n22 191.288
R15722 VDD105.n23 VDD105.t97 191.288
R15723 VDD105.t444 VDD105.n496 191.288
R15724 VDD105.n497 VDD105.t405 191.288
R15725 VDD105.t31 VDD105.n505 191.288
R15726 VDD105.n506 VDD105.t346 191.288
R15727 VDD105.t173 VDD105.n380 138.095
R15728 VDD105.n381 VDD105.t282 138.095
R15729 VDD105.t333 VDD105.n387 138.095
R15730 VDD105.t9 VDD105.n339 138.095
R15731 VDD105.n340 VDD105.t180 138.095
R15732 VDD105.n351 VDD105.t184 138.095
R15733 VDD105.n350 VDD105.t193 138.095
R15734 VDD105.t15 VDD105.n167 138.095
R15735 VDD105.n168 VDD105.t118 138.095
R15736 VDD105.n310 VDD105.t407 138.095
R15737 VDD105.n309 VDD105.t57 138.095
R15738 VDD105.t348 VDD105.t440 120.755
R15739 VDD105.t463 VDD105.t304 120.755
R15740 VDD105.n441 VDD105.t156 111.743
R15741 VDD105.n442 VDD105.t159 111.743
R15742 VDD105.n450 VDD105.t25 111.743
R15743 VDD105.n451 VDD105.t77 111.743
R15744 VDD105.n32 VDD105.t234 111.743
R15745 VDD105.n36 VDD105.t92 111.743
R15746 VDD105.n40 VDD105.t460 111.743
R15747 VDD105.t359 VDD105.n284 111.743
R15748 VDD105.n197 VDD105.t268 111.743
R15749 VDD105.n199 VDD105.t271 111.743
R15750 VDD105.n203 VDD105.t210 111.743
R15751 VDD105.n207 VDD105.t279 111.743
R15752 VDD105.n209 VDD105.t312 111.743
R15753 VDD105.n211 VDD105.t315 111.743
R15754 VDD105.n418 VDD105.t60 111.743
R15755 VDD105.n419 VDD105.t153 111.743
R15756 VDD105.n427 VDD105.t292 111.743
R15757 VDD105.n428 VDD105.t17 111.743
R15758 VDD105.n225 VDD105.t67 111.743
R15759 VDD105.n226 VDD105.t325 111.743
R15760 VDD105.n234 VDD105.t257 111.743
R15761 VDD105.n235 VDD105.t254 111.743
R15762 VDD105.n262 VDD105.t74 111.743
R15763 VDD105.n263 VDD105.t274 111.743
R15764 VDD105.n271 VDD105.t125 111.743
R15765 VDD105.n272 VDD105.t122 111.743
R15766 VDD105.n13 VDD105.t53 111.743
R15767 VDD105.n14 VDD105.t262 111.743
R15768 VDD105.n22 VDD105.t295 111.743
R15769 VDD105.n23 VDD105.t227 111.743
R15770 VDD105.n496 VDD105.t42 111.743
R15771 VDD105.n497 VDD105.t197 111.743
R15772 VDD105.n505 VDD105.t466 111.743
R15773 VDD105.n506 VDD105.t409 111.743
R15774 VDD105.n127 VDD105.t320 109.849
R15775 VDD105.t351 VDD105.n133 109.849
R15776 VDD105.n134 VDD105.t300 109.849
R15777 VDD105.t2 VDD105.n139 109.849
R15778 VDD105.t206 VDD105.n72 109.849
R15779 VDD105.t331 VDD105.n74 109.849
R15780 VDD105.t277 VDD105.n77 109.849
R15781 VDD105.n80 VDD105.t71 109.849
R15782 VDD105.t106 VDD105.n143 109.849
R15783 VDD105.t23 VDD105.n145 109.849
R15784 VDD105.t13 VDD105.n148 109.849
R15785 VDD105.n151 VDD105.t64 109.849
R15786 VDD105.n302 VDD105.t146 109.849
R15787 VDD105.t379 VDD105.n300 109.849
R15788 VDD105.t433 VDD105.n294 109.849
R15789 VDD105.t341 VDD105.n315 109.849
R15790 VDD105.t7 VDD105.n317 109.849
R15791 VDD105.t208 VDD105.n320 109.849
R15792 VDD105.n323 VDD105.t50 109.849
R15793 VDD105.t230 VDD105.n356 109.849
R15794 VDD105.t162 VDD105.n358 109.849
R15795 VDD105.t186 VDD105.n361 109.849
R15796 VDD105.n364 VDD105.t39 109.849
R15797 VDD105.n391 VDD105.t286 105.66
R15798 VDD105.n185 VDD105.t87 105.66
R15799 VDD105.t286 VDD105.t36 63.3967
R15800 VDD105.t87 VDD105.t46 63.3967
R15801 VDD105.n433 VDD105.t441 62.1896
R15802 VDD105.n201 VDD105.t455 62.1896
R15803 VDD105.n213 VDD105.t244 62.1896
R15804 VDD105.n34 VDD105.t322 61.8817
R15805 VDD105.n38 VDD105.t362 61.8817
R15806 VDD105.t150 VDD105.n42 61.5769
R15807 VDD105.n140 VDD105.t412 59.702
R15808 VDD105.n301 VDD105.t11 59.4064
R15809 VDD105.n295 VDD105.t0 59.4064
R15810 VDD105.n290 VDD105.t85 59.1138
R15811 VDD105.n43 VDD105.t108 55.0852
R15812 VDD105.n45 VDD105.t111 55.0852
R15813 VDD105.n286 VDD105.t195 55.0852
R15814 VDD105.t318 VDD105.n289 55.0852
R15815 VDD105.n389 VDD105.n388 45.2835
R15816 VDD105.n190 VDD105.t46 44.5288
R15817 VDD105.n285 VDD105.n190 44.5288
R15818 VDD105.t36 VDD105.n389 43.7741
R15819 VDD105.n81 VDD105.t70 30.9379
R15820 VDD105.n83 VDD105.t49 30.9379
R15821 VDD105.n487 VDD105.t41 30.9379
R15822 VDD105.n461 VDD105.t66 30.9379
R15823 VDD105.n104 VDD105.t56 30.721
R15824 VDD105.n479 VDD105.t59 30.7204
R15825 VDD105.n467 VDD105.t45 30.7203
R15826 VDD105.n94 VDD105.t35 30.7203
R15827 VDD105.n101 VDD105.t63 30.3459
R15828 VDD105.n473 VDD105.t73 30.2877
R15829 VDD105.n483 VDD105.t52 30.2877
R15830 VDD105.n89 VDD105.t38 30.0062
R15831 VDD105.n483 VDD105.t487 24.9141
R15832 VDD105.n101 VDD105.t481 24.8618
R15833 VDD105.n81 VDD105.t479 24.5101
R15834 VDD105.n83 VDD105.t490 24.5101
R15835 VDD105.n487 VDD105.t483 24.5101
R15836 VDD105.n472 VDD105.t477 24.5101
R15837 VDD105.n461 VDD105.t488 24.5101
R15838 VDD105.n104 VDD105.t485 24.4816
R15839 VDD105.n94 VDD105.t476 24.4814
R15840 VDD105.n467 VDD105.t492 24.4814
R15841 VDD105.n479 VDD105.t484 24.4813
R15842 VDD105.n91 VDD105.t493 24.4392
R15843 VDD105.t440 VDD105.n391 15.0948
R15844 VDD105.n185 VDD105.t463 15.0948
R15845 VDD105 VDD105.t428 10.5649
R15846 VDD105 VDD105.t148 10.5649
R15847 VDD105.n91 VDD105.n90 8.0005
R15848 VDD105.n472 VDD105.n471 8.0005
R15849 VDD105 VDD105.t348 7.80993
R15850 VDD105.t304 VDD105 7.80993
R15851 VDD105.n512 VDD105.n510 6.74465
R15852 VDD105.n111 VDD105.n110 6.39748
R15853 VDD105.n488 VDD105.n486 6.39705
R15854 VDD105.n391 VDD105 6.30126
R15855 VDD105 VDD105.n185 6.30126
R15856 VDD105.n115 VDD105.n80 6.3005
R15857 VDD105.n118 VDD105.n77 6.3005
R15858 VDD105.n121 VDD105.n74 6.3005
R15859 VDD105.n124 VDD105.n72 6.3005
R15860 VDD105.n139 VDD105.n138 6.3005
R15861 VDD105.n135 VDD105.n134 6.3005
R15862 VDD105.n133 VDD105.n132 6.3005
R15863 VDD105.n128 VDD105.n127 6.3005
R15864 VDD105.n152 VDD105.n151 6.3005
R15865 VDD105.n155 VDD105.n148 6.3005
R15866 VDD105.n158 VDD105.n145 6.3005
R15867 VDD105.n161 VDD105.n143 6.3005
R15868 VDD105.n225 VDD105.n224 6.3005
R15869 VDD105.n227 VDD105.n226 6.3005
R15870 VDD105.n234 VDD105.n233 6.3005
R15871 VDD105.n236 VDD105.n235 6.3005
R15872 VDD105.n249 VDD105.n203 6.3005
R15873 VDD105.n246 VDD105.n207 6.3005
R15874 VDD105.n243 VDD105.n209 6.3005
R15875 VDD105.n240 VDD105.n211 6.3005
R15876 VDD105.n262 VDD105.n261 6.3005
R15877 VDD105.n264 VDD105.n263 6.3005
R15878 VDD105.n271 VDD105.n270 6.3005
R15879 VDD105.n273 VDD105.n272 6.3005
R15880 VDD105.n284 VDD105.n283 6.3005
R15881 VDD105.n280 VDD105.n197 6.3005
R15882 VDD105.n277 VDD105.n199 6.3005
R15883 VDD105.n190 VDD105.n189 6.3005
R15884 VDD105 VDD105.n286 6.3005
R15885 VDD105.n289 VDD105.n288 6.3005
R15886 VDD105.n294 VDD105.n293 6.3005
R15887 VDD105.n300 VDD105.n299 6.3005
R15888 VDD105.n303 VDD105.n302 6.3005
R15889 VDD105.n309 VDD105.n308 6.3005
R15890 VDD105.n310 VDD105.n172 6.3005
R15891 VDD105.n169 VDD105.n168 6.3005
R15892 VDD105.n167 VDD105.n166 6.3005
R15893 VDD105.n324 VDD105.n323 6.3005
R15894 VDD105.n327 VDD105.n320 6.3005
R15895 VDD105.n330 VDD105.n317 6.3005
R15896 VDD105.n333 VDD105.n315 6.3005
R15897 VDD105.n350 VDD105.n349 6.3005
R15898 VDD105.n351 VDD105.n344 6.3005
R15899 VDD105.n341 VDD105.n340 6.3005
R15900 VDD105.n339 VDD105.n338 6.3005
R15901 VDD105.n365 VDD105.n364 6.3005
R15902 VDD105.n368 VDD105.n361 6.3005
R15903 VDD105.n371 VDD105.n358 6.3005
R15904 VDD105.n374 VDD105.n356 6.3005
R15905 VDD105.n387 VDD105.n386 6.3005
R15906 VDD105.n382 VDD105.n381 6.3005
R15907 VDD105.n380 VDD105.n379 6.3005
R15908 VDD105.n395 VDD105.n389 6.3005
R15909 VDD105 VDD105.n45 6.3005
R15910 VDD105.n398 VDD105.n43 6.3005
R15911 VDD105.n403 VDD105.n40 6.3005
R15912 VDD105.n407 VDD105.n36 6.3005
R15913 VDD105.n411 VDD105.n32 6.3005
R15914 VDD105.n418 VDD105.n417 6.3005
R15915 VDD105.n420 VDD105.n419 6.3005
R15916 VDD105.n427 VDD105.n426 6.3005
R15917 VDD105.n429 VDD105.n428 6.3005
R15918 VDD105.n13 VDD105.n12 6.3005
R15919 VDD105.n15 VDD105.n14 6.3005
R15920 VDD105.n22 VDD105.n21 6.3005
R15921 VDD105.n24 VDD105.n23 6.3005
R15922 VDD105.n507 VDD105.n506 6.3005
R15923 VDD105.n505 VDD105.n504 6.3005
R15924 VDD105.n498 VDD105.n497 6.3005
R15925 VDD105.n496 VDD105.n495 6.3005
R15926 VDD105.n441 VDD105.n440 6.3005
R15927 VDD105.n443 VDD105.n442 6.3005
R15928 VDD105.n450 VDD105.n449 6.3005
R15929 VDD105.n452 VDD105.n451 6.3005
R15930 VDD105.n476 VDD105.n475 5.30733
R15931 VDD105.n100 VDD105.n99 5.30657
R15932 VDD105 VDD105.n509 5.22726
R15933 VDD105.n152 VDD105.t65 5.213
R15934 VDD105.n224 VDD105.n220 5.213
R15935 VDD105.n261 VDD105.n257 5.213
R15936 VDD105.n324 VDD105.t51 5.213
R15937 VDD105.n365 VDD105.t40 5.213
R15938 VDD105.n12 VDD105.n8 5.213
R15939 VDD105 VDD105.t469 5.16454
R15940 VDD105 VDD105.n184 5.16369
R15941 VDD105.n181 VDD105.t319 5.14212
R15942 VDD105.n400 VDD105.n399 5.14212
R15943 VDD105.n28 VDD105.n27 5.13287
R15944 VDD105.n414 VDD105.n413 5.13287
R15945 VDD105.n421 VDD105.t299 5.13287
R15946 VDD105.n422 VDD105.n26 5.13287
R15947 VDD105.n425 VDD105.t224 5.13287
R15948 VDD105.n424 VDD105.n423 5.13287
R15949 VDD105.n430 VDD105.t105 5.13287
R15950 VDD105.n393 VDD105.t37 5.13287
R15951 VDD105.n64 VDD105.t3 5.13287
R15952 VDD105.n136 VDD105.t301 5.13287
R15953 VDD105.n68 VDD105.n67 5.13287
R15954 VDD105.n131 VDD105.t352 5.13287
R15955 VDD105.n130 VDD105.n69 5.13287
R15956 VDD105.n129 VDD105.t321 5.13287
R15957 VDD105.n126 VDD105.n70 5.13287
R15958 VDD105.n117 VDD105.t278 5.13287
R15959 VDD105.n120 VDD105.t332 5.13287
R15960 VDD105.n122 VDD105.n73 5.13287
R15961 VDD105.n123 VDD105.t207 5.13287
R15962 VDD105.n125 VDD105.n71 5.13287
R15963 VDD105.n154 VDD105.t14 5.13287
R15964 VDD105.n157 VDD105.t24 5.13287
R15965 VDD105.n159 VDD105.n144 5.13287
R15966 VDD105.n160 VDD105.t107 5.13287
R15967 VDD105.n162 VDD105.n142 5.13287
R15968 VDD105.n187 VDD105.n183 5.13287
R15969 VDD105.n219 VDD105.n218 5.13287
R15970 VDD105.n229 VDD105.n215 5.13287
R15971 VDD105.n232 VDD105.t115 5.13287
R15972 VDD105.n231 VDD105.n230 5.13287
R15973 VDD105.n237 VDD105.t241 5.13287
R15974 VDD105.n250 VDD105.n202 5.13287
R15975 VDD105.n247 VDD105.n206 5.13287
R15976 VDD105.n245 VDD105.t261 5.13287
R15977 VDD105.n244 VDD105.n208 5.13287
R15978 VDD105.n242 VDD105.t117 5.13287
R15979 VDD105.n241 VDD105.n210 5.13287
R15980 VDD105.n239 VDD105.t253 5.13287
R15981 VDD105.n256 VDD105.n255 5.13287
R15982 VDD105.n266 VDD105.n252 5.13287
R15983 VDD105.n269 VDD105.t371 5.13287
R15984 VDD105.n268 VDD105.n267 5.13287
R15985 VDD105.n274 VDD105.t447 5.13287
R15986 VDD105.n195 VDD105.n191 5.13287
R15987 VDD105.n282 VDD105.t129 5.13287
R15988 VDD105.n281 VDD105.n196 5.13287
R15989 VDD105.n279 VDD105.t373 5.13287
R15990 VDD105.n278 VDD105.n198 5.13287
R15991 VDD105.n276 VDD105.t176 5.13287
R15992 VDD105.n179 VDD105.t434 5.13287
R15993 VDD105.n292 VDD105.n180 5.13287
R15994 VDD105.n298 VDD105.t380 5.13287
R15995 VDD105.n297 VDD105.n178 5.13287
R15996 VDD105.n304 VDD105.t147 5.13287
R15997 VDD105.n176 VDD105.n175 5.13287
R15998 VDD105.n59 VDD105.t58 5.13287
R15999 VDD105.n305 VDD105.t408 5.13287
R16000 VDD105.n171 VDD105.n60 5.13287
R16001 VDD105.n170 VDD105.t119 5.13287
R16002 VDD105.n62 VDD105.n61 5.13287
R16003 VDD105.n165 VDD105.t16 5.13287
R16004 VDD105.n164 VDD105.n63 5.13287
R16005 VDD105.n326 VDD105.t209 5.13287
R16006 VDD105.n329 VDD105.t8 5.13287
R16007 VDD105.n331 VDD105.n316 5.13287
R16008 VDD105.n332 VDD105.t342 5.13287
R16009 VDD105.n334 VDD105.n314 5.13287
R16010 VDD105.n54 VDD105.t194 5.13287
R16011 VDD105.n347 VDD105.t185 5.13287
R16012 VDD105.n343 VDD105.n55 5.13287
R16013 VDD105.n342 VDD105.t181 5.13287
R16014 VDD105.n57 VDD105.n56 5.13287
R16015 VDD105.n337 VDD105.t10 5.13287
R16016 VDD105.n336 VDD105.n58 5.13287
R16017 VDD105.n367 VDD105.t187 5.13287
R16018 VDD105.n370 VDD105.t163 5.13287
R16019 VDD105.n372 VDD105.n357 5.13287
R16020 VDD105.n373 VDD105.t231 5.13287
R16021 VDD105.n375 VDD105.n355 5.13287
R16022 VDD105.n385 VDD105.t334 5.13287
R16023 VDD105.n384 VDD105.n50 5.13287
R16024 VDD105.n383 VDD105.t283 5.13287
R16025 VDD105.n52 VDD105.n51 5.13287
R16026 VDD105.n378 VDD105.t174 5.13287
R16027 VDD105.n377 VDD105.n53 5.13287
R16028 VDD105.n404 VDD105.n39 5.13287
R16029 VDD105.n402 VDD105.t100 5.13287
R16030 VDD105.n408 VDD105.n35 5.13287
R16031 VDD105.n406 VDD105.t233 5.13287
R16032 VDD105.n412 VDD105.n31 5.13287
R16033 VDD105.n410 VDD105.t96 5.13287
R16034 VDD105.n7 VDD105.n6 5.13287
R16035 VDD105.n17 VDD105.n3 5.13287
R16036 VDD105.n20 VDD105.t226 5.13287
R16037 VDD105.n19 VDD105.n18 5.13287
R16038 VDD105.n25 VDD105.t98 5.13287
R16039 VDD105.n434 VDD105.n1 5.13287
R16040 VDD105.n438 VDD105.n437 5.13287
R16041 VDD105.n444 VDD105.t465 5.13287
R16042 VDD105.n445 VDD105.n0 5.13287
R16043 VDD105.n448 VDD105.t34 5.13287
R16044 VDD105.n447 VDD105.n446 5.13287
R16045 VDD105.n453 VDD105.t214 5.13287
R16046 VDD105.n458 VDD105.n457 5.13287
R16047 VDD105.n500 VDD105.n454 5.13287
R16048 VDD105.n503 VDD105.t32 5.13287
R16049 VDD105.n502 VDD105.n501 5.13287
R16050 VDD105.n508 VDD105.t347 5.13287
R16051 VDD105 VDD105.n511 5.13104
R16052 VDD105.n287 VDD105.t196 5.09693
R16053 VDD105.n397 VDD105.n44 5.09693
R16054 VDD105.n141 VDD105.t413 5.09407
R16055 VDD105.n214 VDD105.n212 5.09407
R16056 VDD105.n251 VDD105.n200 5.09407
R16057 VDD105.n291 VDD105.t86 5.09407
R16058 VDD105.n296 VDD105.t1 5.09407
R16059 VDD105.n177 VDD105.t12 5.09407
R16060 VDD105.n313 VDD105.t149 5.09407
R16061 VDD105.n354 VDD105.t429 5.09407
R16062 VDD105.n401 VDD105.n41 5.09407
R16063 VDD105.n405 VDD105.n37 5.09407
R16064 VDD105.n409 VDD105.n33 5.09407
R16065 VDD105.n432 VDD105.n2 5.09407
R16066 VDD105.n114 VDD105.t72 4.8755
R16067 VDD105.n491 VDD105.n490 4.8755
R16068 VDD105.n110 VDD105.n100 4.84121
R16069 VDD105.n486 VDD105.n476 4.84121
R16070 VDD105 VDD105.n512 4.65302
R16071 VDD105.n92 VDD105.n91 4.5005
R16072 VDD105.n95 VDD105.n93 4.5005
R16073 VDD105.n96 VDD105.n93 4.5005
R16074 VDD105.n84 VDD105.n82 4.5005
R16075 VDD105.n85 VDD105.n82 4.5005
R16076 VDD105.n105 VDD105.n103 4.5005
R16077 VDD105.n106 VDD105.n103 4.5005
R16078 VDD105.n466 VDD105.n465 4.5005
R16079 VDD105.n468 VDD105.n465 4.5005
R16080 VDD105.n460 VDD105.n459 4.5005
R16081 VDD105.n462 VDD105.n459 4.5005
R16082 VDD105.n478 VDD105.n477 4.5005
R16083 VDD105.n480 VDD105.n477 4.5005
R16084 VDD105.n392 VDD105 4.40201
R16085 VDD105.n186 VDD105 4.40201
R16086 VDD105.n394 VDD105.n390 3.94862
R16087 VDD105.n188 VDD105.t88 3.94862
R16088 VDD105.n89 VDD105.n88 3.61662
R16089 VDD105.n186 VDD105 3.52487
R16090 VDD105.n392 VDD105 3.47987
R16091 VDD105.n488 VDD105.n487 2.88198
R16092 VDD105.n111 VDD105.n81 2.88182
R16093 VDD105.n194 VDD105.n193 2.88011
R16094 VDD105.n48 VDD105.n47 2.87966
R16095 VDD105.n416 VDD105.n30 2.85787
R16096 VDD105.n137 VDD105.n66 2.85787
R16097 VDD105.n116 VDD105.n79 2.85787
R16098 VDD105.n119 VDD105.n76 2.85787
R16099 VDD105.n153 VDD105.n150 2.85787
R16100 VDD105.n156 VDD105.n147 2.85787
R16101 VDD105.n223 VDD105.n222 2.85787
R16102 VDD105.n228 VDD105.n217 2.85787
R16103 VDD105.n248 VDD105.n205 2.85787
R16104 VDD105.n260 VDD105.n259 2.85787
R16105 VDD105.n265 VDD105.n254 2.85787
R16106 VDD105.n307 VDD105.n174 2.85787
R16107 VDD105.n325 VDD105.n322 2.85787
R16108 VDD105.n328 VDD105.n319 2.85787
R16109 VDD105.n348 VDD105.n346 2.85787
R16110 VDD105.n366 VDD105.n363 2.85787
R16111 VDD105.n369 VDD105.n360 2.85787
R16112 VDD105.n11 VDD105.n10 2.85787
R16113 VDD105.n16 VDD105.n5 2.85787
R16114 VDD105.n439 VDD105.n436 2.85787
R16115 VDD105.n494 VDD105.n493 2.85787
R16116 VDD105.n499 VDD105.n456 2.85787
R16117 VDD105.n30 VDD105.t243 2.2755
R16118 VDD105.n30 VDD105.n29 2.2755
R16119 VDD105.n47 VDD105.t436 2.2755
R16120 VDD105.n47 VDD105.n46 2.2755
R16121 VDD105.n66 VDD105.t189 2.2755
R16122 VDD105.n66 VDD105.n65 2.2755
R16123 VDD105.n79 VDD105.t369 2.2755
R16124 VDD105.n79 VDD105.n78 2.2755
R16125 VDD105.n76 VDD105.t350 2.2755
R16126 VDD105.n76 VDD105.n75 2.2755
R16127 VDD105.n150 VDD105.t378 2.2755
R16128 VDD105.n150 VDD105.n149 2.2755
R16129 VDD105.n147 VDD105.t121 2.2755
R16130 VDD105.n147 VDD105.n146 2.2755
R16131 VDD105.n193 VDD105.t303 2.2755
R16132 VDD105.n193 VDD105.n192 2.2755
R16133 VDD105.n222 VDD105.t451 2.2755
R16134 VDD105.n222 VDD105.n221 2.2755
R16135 VDD105.n217 VDD105.t396 2.2755
R16136 VDD105.n217 VDD105.n216 2.2755
R16137 VDD105.n205 VDD105.t449 2.2755
R16138 VDD105.n205 VDD105.n204 2.2755
R16139 VDD105.n259 VDD105.t308 2.2755
R16140 VDD105.n259 VDD105.n258 2.2755
R16141 VDD105.n254 VDD105.t398 2.2755
R16142 VDD105.n254 VDD105.n253 2.2755
R16143 VDD105.n174 VDD105.t84 2.2755
R16144 VDD105.n174 VDD105.n173 2.2755
R16145 VDD105.n322 VDD105.t142 2.2755
R16146 VDD105.n322 VDD105.n321 2.2755
R16147 VDD105.n319 VDD105.t183 2.2755
R16148 VDD105.n319 VDD105.n318 2.2755
R16149 VDD105.n346 VDD105.t222 2.2755
R16150 VDD105.n346 VDD105.n345 2.2755
R16151 VDD105.n363 VDD105.t427 2.2755
R16152 VDD105.n363 VDD105.n362 2.2755
R16153 VDD105.n360 VDD105.t285 2.2755
R16154 VDD105.n360 VDD105.n359 2.2755
R16155 VDD105.n10 VDD105.t248 2.2755
R16156 VDD105.n10 VDD105.n9 2.2755
R16157 VDD105.n5 VDD105.t391 2.2755
R16158 VDD105.n5 VDD105.n4 2.2755
R16159 VDD105.n436 VDD105.t459 2.2755
R16160 VDD105.n436 VDD105.n435 2.2755
R16161 VDD105.n493 VDD105.t445 2.2755
R16162 VDD105.n493 VDD105.n492 2.2755
R16163 VDD105.n456 VDD105.t406 2.2755
R16164 VDD105.n456 VDD105.n455 2.2755
R16165 VDD105.n98 VDD105.n97 2.2439
R16166 VDD105.n108 VDD105.n107 2.2439
R16167 VDD105.n470 VDD105.n469 2.2439
R16168 VDD105.n482 VDD105.n481 2.2439
R16169 VDD105.n87 VDD105.n86 2.24362
R16170 VDD105.n464 VDD105.n463 2.24362
R16171 VDD105.n462 VDD105.n461 2.12269
R16172 VDD105.n84 VDD105.n83 2.12257
R16173 VDD105.n474 VDD105.n473 1.82213
R16174 VDD105.n484 VDD105.n483 1.82213
R16175 VDD105 VDD105.n28 1.81843
R16176 VDD105 VDD105.n250 1.81843
R16177 VDD105 VDD105.n404 1.81843
R16178 VDD105 VDD105.n408 1.81843
R16179 VDD105.n434 VDD105 1.81843
R16180 VDD105.n102 VDD105.n101 1.81789
R16181 VDD105 VDD105.n64 1.77285
R16182 VDD105 VDD105.n179 1.77285
R16183 VDD105.n298 VDD105 1.77285
R16184 VDD105 VDD105.n59 1.77285
R16185 VDD105 VDD105.n54 1.77285
R16186 VDD105.n99 VDD105.n98 1.62565
R16187 VDD105.n109 VDD105.n108 1.62565
R16188 VDD105.n485 VDD105.n482 1.6239
R16189 VDD105.n475 VDD105.n470 1.6239
R16190 VDD105.n480 VDD105.n479 1.39892
R16191 VDD105.n468 VDD105.n467 1.3985
R16192 VDD105.n105 VDD105.n104 1.39782
R16193 VDD105.n95 VDD105.n94 1.39728
R16194 VDD105.n126 VDD105.n125 1.16167
R16195 VDD105.n475 VDD105.n474 1.12224
R16196 VDD105.n99 VDD105.n92 1.12171
R16197 VDD105.n109 VDD105.n102 1.12171
R16198 VDD105.n485 VDD105.n484 1.12167
R16199 VDD105.n163 VDD105.n162 1.07428
R16200 VDD105.n335 VDD105.n334 1.07428
R16201 VDD105.n376 VDD105.n375 1.07428
R16202 VDD105.n238 VDD105.n237 1.0737
R16203 VDD105.n275 VDD105.n274 1.0737
R16204 VDD105.n431 VDD105.n25 1.0737
R16205 VDD105.n509 VDD105.n508 1.03044
R16206 VDD105.n91 VDD105.n89 0.840632
R16207 VDD105.n415 VDD105.n412 0.715235
R16208 VDD105.n491 VDD105.n489 0.603658
R16209 VDD105.n486 VDD105.n485 0.523557
R16210 VDD105.n110 VDD105.n109 0.5228
R16211 VDD105.n100 VDD105.n87 0.497812
R16212 VDD105.n476 VDD105.n464 0.497812
R16213 VDD105 VDD105.n304 0.434967
R16214 VDD105.n473 VDD105.n472 0.404541
R16215 VDD105 VDD105.n396 0.339236
R16216 VDD105 VDD105.n182 0.338387
R16217 VDD105.n115 VDD105.n114 0.337997
R16218 VDD105.n495 VDD105.n491 0.337997
R16219 VDD105 VDD105.n181 0.334577
R16220 VDD105 VDD105.n400 0.334577
R16221 VDD105.n114 VDD105.n113 0.333658
R16222 VDD105.n398 VDD105.n397 0.318198
R16223 VDD105.n288 VDD105.n287 0.317357
R16224 VDD105.n306 VDD105 0.280768
R16225 VDD105.n120 VDD105.n119 0.233919
R16226 VDD105.n117 VDD105.n116 0.233919
R16227 VDD105.n157 VDD105.n156 0.233919
R16228 VDD105.n154 VDD105.n153 0.233919
R16229 VDD105.n223 VDD105.n219 0.233919
R16230 VDD105.n229 VDD105.n228 0.233919
R16231 VDD105.n260 VDD105.n256 0.233919
R16232 VDD105.n266 VDD105.n265 0.233919
R16233 VDD105.n329 VDD105.n328 0.233919
R16234 VDD105.n326 VDD105.n325 0.233919
R16235 VDD105.n370 VDD105.n369 0.233919
R16236 VDD105.n367 VDD105.n366 0.233919
R16237 VDD105.n11 VDD105.n7 0.233919
R16238 VDD105.n17 VDD105.n16 0.233919
R16239 VDD105.n494 VDD105.n458 0.233919
R16240 VDD105.n500 VDD105.n499 0.233919
R16241 VDD105.n402 VDD105.n401 0.170499
R16242 VDD105.n406 VDD105.n405 0.170499
R16243 VDD105.n410 VDD105.n409 0.170499
R16244 VDD105.n292 VDD105.n291 0.170231
R16245 VDD105.n297 VDD105.n296 0.170231
R16246 VDD105.n177 VDD105.n176 0.170231
R16247 VDD105.n287 VDD105 0.147133
R16248 VDD105.n397 VDD105 0.146292
R16249 VDD105.n239 VDD105.n238 0.143967
R16250 VDD105.n276 VDD105.n275 0.143967
R16251 VDD105.n431 VDD105.n430 0.143967
R16252 VDD105.n164 VDD105.n163 0.143501
R16253 VDD105.n336 VDD105.n335 0.143501
R16254 VDD105.n377 VDD105.n376 0.143501
R16255 VDD105.n512 VDD105 0.142752
R16256 VDD105.n123 VDD105.n122 0.141016
R16257 VDD105.n130 VDD105.n129 0.141016
R16258 VDD105.n131 VDD105.n68 0.141016
R16259 VDD105.n160 VDD105.n159 0.141016
R16260 VDD105.n232 VDD105.n231 0.141016
R16261 VDD105.n245 VDD105.n244 0.141016
R16262 VDD105.n242 VDD105.n241 0.141016
R16263 VDD105.n269 VDD105.n268 0.141016
R16264 VDD105.n282 VDD105.n281 0.141016
R16265 VDD105.n279 VDD105.n278 0.141016
R16266 VDD105.n165 VDD105.n62 0.141016
R16267 VDD105.n171 VDD105.n170 0.141016
R16268 VDD105.n332 VDD105.n331 0.141016
R16269 VDD105.n337 VDD105.n57 0.141016
R16270 VDD105.n343 VDD105.n342 0.141016
R16271 VDD105.n373 VDD105.n372 0.141016
R16272 VDD105.n378 VDD105.n52 0.141016
R16273 VDD105.n384 VDD105.n383 0.141016
R16274 VDD105.n422 VDD105.n421 0.141016
R16275 VDD105.n425 VDD105.n424 0.141016
R16276 VDD105.n20 VDD105.n19 0.141016
R16277 VDD105.n503 VDD105.n502 0.141016
R16278 VDD105.n445 VDD105.n444 0.141016
R16279 VDD105.n448 VDD105.n447 0.141016
R16280 VDD105.n238 VDD105.n214 0.139745
R16281 VDD105.n432 VDD105.n431 0.139745
R16282 VDD105.n163 VDD105.n141 0.138896
R16283 VDD105.n335 VDD105.n313 0.138896
R16284 VDD105.n509 VDD105.n453 0.130565
R16285 VDD105 VDD105.n251 0.128708
R16286 VDD105 VDD105.n354 0.127858
R16287 VDD105 VDD105.n247 0.123016
R16288 VDD105.n195 VDD105 0.123016
R16289 VDD105 VDD105.n438 0.123016
R16290 VDD105 VDD105.n136 0.122435
R16291 VDD105 VDD105.n347 0.122435
R16292 VDD105.n385 VDD105 0.122435
R16293 VDD105.n484 VDD105 0.112066
R16294 VDD105.n137 VDD105 0.111984
R16295 VDD105.n307 VDD105 0.111984
R16296 VDD105.n348 VDD105 0.111984
R16297 VDD105.n489 VDD105 0.111564
R16298 VDD105.n248 VDD105 0.111403
R16299 VDD105.n416 VDD105 0.111403
R16300 VDD105.n439 VDD105 0.111403
R16301 VDD105.n102 VDD105 0.110941
R16302 VDD105 VDD105.n48 0.108832
R16303 VDD105 VDD105.n194 0.108613
R16304 VDD105.n125 VDD105.n124 0.107339
R16305 VDD105.n122 VDD105.n121 0.107339
R16306 VDD105.n128 VDD105.n126 0.107339
R16307 VDD105.n132 VDD105.n130 0.107339
R16308 VDD105.n135 VDD105.n68 0.107339
R16309 VDD105.n162 VDD105.n161 0.107339
R16310 VDD105.n159 VDD105.n158 0.107339
R16311 VDD105.n233 VDD105.n232 0.107339
R16312 VDD105.n237 VDD105.n236 0.107339
R16313 VDD105.n246 VDD105.n245 0.107339
R16314 VDD105.n243 VDD105.n242 0.107339
R16315 VDD105.n240 VDD105.n239 0.107339
R16316 VDD105.n270 VDD105.n269 0.107339
R16317 VDD105.n274 VDD105.n273 0.107339
R16318 VDD105.n283 VDD105.n282 0.107339
R16319 VDD105.n280 VDD105.n279 0.107339
R16320 VDD105.n277 VDD105.n276 0.107339
R16321 VDD105.n293 VDD105.n292 0.107339
R16322 VDD105.n299 VDD105.n297 0.107339
R16323 VDD105.n303 VDD105.n176 0.107339
R16324 VDD105.n166 VDD105.n164 0.107339
R16325 VDD105.n169 VDD105.n62 0.107339
R16326 VDD105.n172 VDD105.n171 0.107339
R16327 VDD105.n334 VDD105.n333 0.107339
R16328 VDD105.n331 VDD105.n330 0.107339
R16329 VDD105.n338 VDD105.n336 0.107339
R16330 VDD105.n341 VDD105.n57 0.107339
R16331 VDD105.n344 VDD105.n343 0.107339
R16332 VDD105.n375 VDD105.n374 0.107339
R16333 VDD105.n372 VDD105.n371 0.107339
R16334 VDD105.n379 VDD105.n377 0.107339
R16335 VDD105.n382 VDD105.n52 0.107339
R16336 VDD105.n386 VDD105.n384 0.107339
R16337 VDD105.n403 VDD105.n402 0.107339
R16338 VDD105.n407 VDD105.n406 0.107339
R16339 VDD105.n411 VDD105.n410 0.107339
R16340 VDD105.n421 VDD105.n420 0.107339
R16341 VDD105.n426 VDD105.n425 0.107339
R16342 VDD105.n430 VDD105.n429 0.107339
R16343 VDD105.n21 VDD105.n20 0.107339
R16344 VDD105.n25 VDD105.n24 0.107339
R16345 VDD105.n504 VDD105.n503 0.107339
R16346 VDD105.n508 VDD105.n507 0.107339
R16347 VDD105.n444 VDD105.n443 0.107339
R16348 VDD105.n449 VDD105.n448 0.107339
R16349 VDD105.n453 VDD105.n452 0.107339
R16350 VDD105 VDD105.n223 0.106758
R16351 VDD105.n228 VDD105 0.106758
R16352 VDD105 VDD105.n248 0.106758
R16353 VDD105 VDD105.n260 0.106758
R16354 VDD105.n265 VDD105 0.106758
R16355 VDD105 VDD105.n416 0.106758
R16356 VDD105 VDD105.n11 0.106758
R16357 VDD105.n16 VDD105 0.106758
R16358 VDD105 VDD105.n494 0.106758
R16359 VDD105.n499 VDD105 0.106758
R16360 VDD105 VDD105.n439 0.106758
R16361 VDD105.n119 VDD105 0.106177
R16362 VDD105.n116 VDD105 0.106177
R16363 VDD105 VDD105.n137 0.106177
R16364 VDD105.n156 VDD105 0.106177
R16365 VDD105.n153 VDD105 0.106177
R16366 VDD105 VDD105.n307 0.106177
R16367 VDD105.n328 VDD105 0.106177
R16368 VDD105.n325 VDD105 0.106177
R16369 VDD105 VDD105.n348 0.106177
R16370 VDD105.n369 VDD105 0.106177
R16371 VDD105.n366 VDD105 0.106177
R16372 VDD105.n471 VDD105 0.0850665
R16373 VDD105.n90 VDD105 0.0839415
R16374 VDD105 VDD105.n415 0.0829516
R16375 VDD105 VDD105.n306 0.082371
R16376 VDD105.n96 VDD105 0.0816915
R16377 VDD105.n466 VDD105 0.0816915
R16378 VDD105.n118 VDD105.n117 0.080629
R16379 VDD105.n138 VDD105.n64 0.080629
R16380 VDD105.n155 VDD105.n154 0.080629
R16381 VDD105.n227 VDD105.n219 0.080629
R16382 VDD105.n250 VDD105.n249 0.080629
R16383 VDD105.n264 VDD105.n256 0.080629
R16384 VDD105.n308 VDD105.n59 0.080629
R16385 VDD105.n327 VDD105.n326 0.080629
R16386 VDD105.n349 VDD105.n54 0.080629
R16387 VDD105.n368 VDD105.n367 0.080629
R16388 VDD105.n417 VDD105.n28 0.080629
R16389 VDD105.n15 VDD105.n7 0.080629
R16390 VDD105.n498 VDD105.n458 0.080629
R16391 VDD105.n440 VDD105.n434 0.080629
R16392 VDD105.n106 VDD105 0.0805665
R16393 VDD105.n478 VDD105 0.0805665
R16394 VDD105 VDD105.n123 0.0794677
R16395 VDD105 VDD105.n120 0.0794677
R16396 VDD105.n129 VDD105 0.0794677
R16397 VDD105 VDD105.n131 0.0794677
R16398 VDD105.n136 VDD105 0.0794677
R16399 VDD105 VDD105.n160 0.0794677
R16400 VDD105 VDD105.n157 0.0794677
R16401 VDD105 VDD105.n165 0.0794677
R16402 VDD105.n170 VDD105 0.0794677
R16403 VDD105.n305 VDD105 0.0794677
R16404 VDD105 VDD105.n332 0.0794677
R16405 VDD105 VDD105.n329 0.0794677
R16406 VDD105 VDD105.n337 0.0794677
R16407 VDD105.n342 VDD105 0.0794677
R16408 VDD105.n347 VDD105 0.0794677
R16409 VDD105 VDD105.n373 0.0794677
R16410 VDD105 VDD105.n370 0.0794677
R16411 VDD105 VDD105.n378 0.0794677
R16412 VDD105.n383 VDD105 0.0794677
R16413 VDD105 VDD105.n385 0.0794677
R16414 VDD105 VDD105.n181 0.0794623
R16415 VDD105.n400 VDD105 0.0794623
R16416 VDD105 VDD105.n229 0.0788871
R16417 VDD105.n231 VDD105 0.0788871
R16418 VDD105.n247 VDD105 0.0788871
R16419 VDD105.n244 VDD105 0.0788871
R16420 VDD105.n241 VDD105 0.0788871
R16421 VDD105 VDD105.n266 0.0788871
R16422 VDD105.n268 VDD105 0.0788871
R16423 VDD105 VDD105.n195 0.0788871
R16424 VDD105.n281 VDD105 0.0788871
R16425 VDD105.n278 VDD105 0.0788871
R16426 VDD105.n414 VDD105 0.0788871
R16427 VDD105 VDD105.n422 0.0788871
R16428 VDD105.n424 VDD105 0.0788871
R16429 VDD105 VDD105.n17 0.0788871
R16430 VDD105.n19 VDD105 0.0788871
R16431 VDD105 VDD105.n500 0.0788871
R16432 VDD105.n502 VDD105 0.0788871
R16433 VDD105.n438 VDD105 0.0788871
R16434 VDD105 VDD105.n445 0.0788871
R16435 VDD105.n447 VDD105 0.0788871
R16436 VDD105 VDD105.n179 0.0759839
R16437 VDD105 VDD105.n298 0.0759839
R16438 VDD105.n304 VDD105 0.0759839
R16439 VDD105.n404 VDD105 0.0754032
R16440 VDD105.n408 VDD105 0.0754032
R16441 VDD105.n412 VDD105 0.0754032
R16442 VDD105.n460 VDD105 0.0749415
R16443 VDD105.n85 VDD105 0.0738165
R16444 VDD105.n113 VDD105.n111 0.0725
R16445 VDD105.n141 VDD105 0.0709717
R16446 VDD105.n291 VDD105 0.0709717
R16447 VDD105.n296 VDD105 0.0709717
R16448 VDD105 VDD105.n177 0.0709717
R16449 VDD105.n313 VDD105 0.0709717
R16450 VDD105.n354 VDD105 0.0709717
R16451 VDD105.n214 VDD105 0.0701226
R16452 VDD105.n251 VDD105 0.0701226
R16453 VDD105.n401 VDD105 0.0701226
R16454 VDD105.n405 VDD105 0.0701226
R16455 VDD105.n409 VDD105 0.0701226
R16456 VDD105 VDD105.n432 0.0701226
R16457 VDD105.n112 VDD105 0.0700455
R16458 VDD105 VDD105.n182 0.0491131
R16459 VDD105.n396 VDD105 0.0487847
R16460 VDD105.n113 VDD105.n112 0.0455
R16461 VDD105.n187 VDD105.n186 0.0409015
R16462 VDD105.n393 VDD105.n392 0.040573
R16463 VDD105.n306 VDD105.n305 0.0405645
R16464 VDD105.n415 VDD105.n414 0.0405645
R16465 VDD105.n489 VDD105.n488 0.0344894
R16466 VDD105.n97 VDD105.n96 0.0275
R16467 VDD105.n90 VDD105.n88 0.0275
R16468 VDD105.n469 VDD105.n466 0.0275
R16469 VDD105.n474 VDD105.n471 0.0275
R16470 VDD105.n107 VDD105.n106 0.026375
R16471 VDD105.n481 VDD105.n478 0.026375
R16472 VDD105.n98 VDD105.n93 0.025705
R16473 VDD105.n108 VDD105.n103 0.025705
R16474 VDD105.n470 VDD105.n465 0.025705
R16475 VDD105.n482 VDD105.n477 0.025705
R16476 VDD105.n188 VDD105.n187 0.025135
R16477 VDD105.n394 VDD105.n393 0.025135
R16478 VDD105.n189 VDD105.n188 0.0211934
R16479 VDD105.n395 VDD105.n394 0.0211934
R16480 VDD105.n86 VDD105.n85 0.02075
R16481 VDD105.n463 VDD105.n460 0.019625
R16482 VDD105.n87 VDD105.n82 0.0169383
R16483 VDD105.n464 VDD105.n459 0.0169383
R16484 VDD105.n396 VDD105.n48 0.0132147
R16485 VDD105.n194 VDD105.n182 0.0131133
R16486 VDD105.n275 VDD105 0.0115377
R16487 VDD105.n376 VDD105 0.0115377
R16488 VDD105.n463 VDD105.n462 0.010625
R16489 VDD105.n86 VDD105.n84 0.0095
R16490 VDD105 VDD105.n403 0.00572581
R16491 VDD105 VDD105.n407 0.00572581
R16492 VDD105 VDD105.n411 0.00572581
R16493 VDD105.n293 VDD105 0.00514516
R16494 VDD105.n299 VDD105 0.00514516
R16495 VDD105 VDD105.n303 0.00514516
R16496 VDD105.n112 VDD105 0.00459091
R16497 VDD105.n107 VDD105.n105 0.003875
R16498 VDD105.n481 VDD105.n480 0.003875
R16499 VDD105.n97 VDD105.n95 0.00275
R16500 VDD105.n469 VDD105.n468 0.00275
R16501 VDD105.n233 VDD105 0.00224194
R16502 VDD105.n236 VDD105 0.00224194
R16503 VDD105 VDD105.n246 0.00224194
R16504 VDD105 VDD105.n243 0.00224194
R16505 VDD105 VDD105.n240 0.00224194
R16506 VDD105.n270 VDD105 0.00224194
R16507 VDD105.n273 VDD105 0.00224194
R16508 VDD105.n283 VDD105 0.00224194
R16509 VDD105 VDD105.n280 0.00224194
R16510 VDD105 VDD105.n277 0.00224194
R16511 VDD105.n420 VDD105 0.00224194
R16512 VDD105.n426 VDD105 0.00224194
R16513 VDD105.n429 VDD105 0.00224194
R16514 VDD105.n21 VDD105 0.00224194
R16515 VDD105.n24 VDD105 0.00224194
R16516 VDD105.n504 VDD105 0.00224194
R16517 VDD105.n507 VDD105 0.00224194
R16518 VDD105.n443 VDD105 0.00224194
R16519 VDD105.n449 VDD105 0.00224194
R16520 VDD105.n452 VDD105 0.00224194
R16521 VDD105.n288 VDD105 0.00219811
R16522 VDD105 VDD105.n398 0.00219811
R16523 VDD105.n124 VDD105 0.00166129
R16524 VDD105.n121 VDD105 0.00166129
R16525 VDD105 VDD105.n118 0.00166129
R16526 VDD105 VDD105.n115 0.00166129
R16527 VDD105 VDD105.n128 0.00166129
R16528 VDD105.n132 VDD105 0.00166129
R16529 VDD105 VDD105.n135 0.00166129
R16530 VDD105.n138 VDD105 0.00166129
R16531 VDD105.n161 VDD105 0.00166129
R16532 VDD105.n158 VDD105 0.00166129
R16533 VDD105 VDD105.n155 0.00166129
R16534 VDD105 VDD105.n152 0.00166129
R16535 VDD105.n166 VDD105 0.00166129
R16536 VDD105 VDD105.n169 0.00166129
R16537 VDD105 VDD105.n172 0.00166129
R16538 VDD105.n308 VDD105 0.00166129
R16539 VDD105.n333 VDD105 0.00166129
R16540 VDD105.n330 VDD105 0.00166129
R16541 VDD105 VDD105.n327 0.00166129
R16542 VDD105 VDD105.n324 0.00166129
R16543 VDD105.n338 VDD105 0.00166129
R16544 VDD105 VDD105.n341 0.00166129
R16545 VDD105 VDD105.n344 0.00166129
R16546 VDD105.n349 VDD105 0.00166129
R16547 VDD105.n374 VDD105 0.00166129
R16548 VDD105.n371 VDD105 0.00166129
R16549 VDD105 VDD105.n368 0.00166129
R16550 VDD105 VDD105.n365 0.00166129
R16551 VDD105.n379 VDD105 0.00166129
R16552 VDD105 VDD105.n382 0.00166129
R16553 VDD105.n386 VDD105 0.00166129
R16554 VDD105.n92 VDD105.n88 0.001625
R16555 VDD105 VDD105.n395 0.00115693
R16556 VDD105.n224 VDD105 0.00108064
R16557 VDD105 VDD105.n227 0.00108064
R16558 VDD105.n249 VDD105 0.00108064
R16559 VDD105.n261 VDD105 0.00108064
R16560 VDD105 VDD105.n264 0.00108064
R16561 VDD105.n417 VDD105 0.00108064
R16562 VDD105.n12 VDD105 0.00108064
R16563 VDD105 VDD105.n15 0.00108064
R16564 VDD105.n495 VDD105 0.00108064
R16565 VDD105 VDD105.n498 0.00108064
R16566 VDD105.n440 VDD105 0.00108064
R16567 VDD105.n189 VDD105 0.000828467
R16568 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t7 37.1981
R16569 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n4 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t3 31.528
R16570 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t6 30.5752
R16571 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t5 24.6493
R16572 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t8 17.6611
R16573 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 17.0533
R16574 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n4 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t4 15.3826
R16575 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n4 7.62758
R16576 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n5 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n3 3.28711
R16577 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n7 2.99416
R16578 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 2.81128
R16579 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n5 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 2.66613
R16580 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n7 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t1 2.2755
R16581 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n7 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n6 2.2755
R16582 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n5 2.2505
R16583 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n1 1.80834
R16584 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n2 1.43706
R16585 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n0 0.281955
R16586 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n8 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t2 36.935
R16587 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n7 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t9 36.935
R16588 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n12 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t8 36.935
R16589 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n9 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t5 36.935
R16590 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n10 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t10 30.5752
R16591 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n13 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t3 25.4744
R16592 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n6 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t13 25.4742
R16593 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n10 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t12 21.7814
R16594 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n8 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t14 18.1962
R16595 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n7 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t7 18.1962
R16596 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n12 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t6 18.1962
R16597 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n9 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t15 18.1962
R16598 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n6 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t4 14.142
R16599 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n13 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t11 14.1417
R16600 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n5 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t1 9.33985
R16601 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n0 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n11 7.41483
R16602 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n15 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n14 5.37091
R16603 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n5 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t0 5.17836
R16604 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n2 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n12 2.13265
R16605 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n2 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK 0.077103
R16606 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n13 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n3 1.42996
R16607 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n0 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n2 1.11863
R16608 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n14 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n3 1.19586
R16609 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n8 2.13265
R16610 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n11 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n10 1.80883
R16611 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n1 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK 2.63776
R16612 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n0 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK 2.51943
R16613 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n9 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK 2.13281
R16614 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n7 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK 2.13261
R16615 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n4 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n6 1.43004
R16616 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n3 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK 0.196041
R16617 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n4 0.196041
R16618 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n5 0.115328
R16619 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n11 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK 0.108371
R16620 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n4 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n15 1.19586
R16621 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n1 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK 1.11863
R16622 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n14 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n0 1.01264
R16623 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n15 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n1 0.894314
R16624 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n5 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.t6 36.935
R16625 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n2 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.t9 31.4332
R16626 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n6 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.t7 31.4332
R16627 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n3 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.t3 30.4613
R16628 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n3 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.t5 24.7562
R16629 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n5 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.t10 18.1962
R16630 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n2 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.t8 15.3826
R16631 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n6 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.t4 15.3826
R16632 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n4 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1 8.5575
R16633 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.t1 7.09905
R16634 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n6 6.86029
R16635 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n2 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1 5.69501
R16636 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n7 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1 5.01077
R16637 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n1 3.25053
R16638 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n8 2.43532
R16639 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n1 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.t2 2.2755
R16640 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n1 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n0 2.2755
R16641 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n5 2.13459
R16642 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n3 1.81638
R16643 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n8 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n7 1.45395
R16644 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n8 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n4 1.23718
R16645 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n7 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1 1.12067
R16646 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n4 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1 0.976433
R16647 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t8 37.1986
R16648 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t6 31.528
R16649 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n3 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t3 30.6315
R16650 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n3 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t4 24.5953
R16651 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t5 17.6614
R16652 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n4 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 17.0516
R16653 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t7 15.3826
R16654 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n1 7.62751
R16655 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n5 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n4 3.28711
R16656 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n7 2.99416
R16657 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n4 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 2.81128
R16658 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n5 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 2.67866
R16659 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n7 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t1 2.2755
R16660 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n7 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n6 2.2755
R16661 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n5 2.2505
R16662 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n3 1.80496
R16663 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n2 1.43709
R16664 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n0 0.281955
R16665 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n5 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.t4 36.935
R16666 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n2 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.t7 31.4332
R16667 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n6 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.t3 31.4332
R16668 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n3 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.t10 30.4613
R16669 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n3 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.t6 24.7562
R16670 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n5 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.t9 18.1962
R16671 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n2 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.t5 15.3826
R16672 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n6 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.t8 15.3826
R16673 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n4 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1 8.5575
R16674 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.t1 7.09905
R16675 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n6 6.86029
R16676 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n2 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1 5.69501
R16677 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n7 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1 5.01077
R16678 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n1 3.25053
R16679 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n8 2.43532
R16680 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n1 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.t0 2.2755
R16681 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n1 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n0 2.2755
R16682 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n5 2.13459
R16683 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n3 1.81638
R16684 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n8 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n7 1.45395
R16685 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n8 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n4 1.23718
R16686 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n7 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1 1.12067
R16687 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n4 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1 0.976433
R16688 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.n2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.t5 37.1981
R16689 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.n1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.t3 31.528
R16690 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.n2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.t6 17.6611
R16691 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.n1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.t4 15.3826
R16692 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.n1 7.62751
R16693 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.n3 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB 6.09789
R16694 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.n0 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.n5 2.99416
R16695 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.n3 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB 2.67866
R16696 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.n5 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.t0 2.2755
R16697 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.n5 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.n4 2.2755
R16698 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.n0 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.n3 2.2505
R16699 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.n2 1.43706
R16700 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.n0 0.281955
R16701 Vdiv96.n3 Vdiv96.t2 31.528
R16702 Vdiv96.n3 Vdiv96.t3 15.3826
R16703 Vdiv96 Vdiv96.n8 10.9696
R16704 Vdiv96.n11 Vdiv96.n10 9.33985
R16705 Vdiv96.n4 Vdiv96.n3 5.60588
R16706 Vdiv96.n11 Vdiv96.n9 5.17836
R16707 Vdiv96.n6 Vdiv96.n0 4.52731
R16708 Vdiv96.n6 Vdiv96.n5 4.5005
R16709 Vdiv96.n8 Vdiv96.n7 4.5005
R16710 Vdiv96.n1 Vdiv96.n0 1.50562
R16711 Vdiv96.n2 Vdiv96.n1 0.899631
R16712 Vdiv96.n2 Vdiv96 0.0781829
R16713 Vdiv96 Vdiv96.n11 0.0749828
R16714 Vdiv96 Vdiv96.n2 0.0376545
R16715 Vdiv96.n8 Vdiv96.n0 0.0266
R16716 Vdiv96.n7 Vdiv96.n6 0.00624468
R16717 Vdiv96.n7 Vdiv96.n1 0.00260066
R16718 Vdiv96.n5 Vdiv96 0.00197541
R16719 Vdiv96.n4 Vdiv96 0.00189862
R16720 Vdiv96.n5 Vdiv96.n4 0.00157662
R16721 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n3 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t7 37.1981
R16722 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n5 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t4 31.4332
R16723 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n2 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t6 30.5752
R16724 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n2 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t2 24.6493
R16725 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n3 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t5 17.6611
R16726 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n4 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 17.0516
R16727 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n5 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t3 15.3826
R16728 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n5 7.62776
R16729 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n6 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n4 3.28711
R16730 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n7 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n1 2.99416
R16731 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n4 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 2.81128
R16732 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n6 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 2.67895
R16733 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t0 2.2755
R16734 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n0 2.2755
R16735 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n7 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n6 2.2505
R16736 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n2 1.80883
R16737 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n3 1.43706
R16738 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n7 0.4325
R16739 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n5 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.t5 36.935
R16740 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n4 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.t3 31.4332
R16741 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n6 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.t9 31.4332
R16742 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n3 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.t10 30.5184
R16743 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n3 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.t8 24.7029
R16744 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n5 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.t4 18.1962
R16745 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n4 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.t7 15.3826
R16746 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n6 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.t6 15.3826
R16747 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.t2 7.09905
R16748 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n6 6.86134
R16749 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n7 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1 5.0096
R16750 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n0 8.55639
R16751 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n4 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1 5.69501
R16752 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n2 3.25226
R16753 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n8 2.43532
R16754 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.t0 2.2755
R16755 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n1 2.2755
R16756 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n5 2.13479
R16757 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n3 1.81225
R16758 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n8 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n7 1.45511
R16759 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n8 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n0 1.23718
R16760 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n7 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1 1.12056
R16761 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n0 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1 0.976034
R16762 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n10 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t9 36.935
R16763 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n9 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t13 36.935
R16764 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n14 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t3 36.935
R16765 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n11 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t6 36.935
R16766 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n12 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t11 30.5752
R16767 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n18 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t14 25.4742
R16768 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n15 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t2 25.4742
R16769 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n12 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t8 21.7814
R16770 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n10 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t12 18.1962
R16771 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n9 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t15 18.1962
R16772 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n14 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t4 18.1962
R16773 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n11 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t7 18.1962
R16774 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n18 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t5 14.142
R16775 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n15 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t10 14.142
R16776 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n8 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t1 9.33985
R16777 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n0 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n13 7.41653
R16778 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n17 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n16 5.37091
R16779 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n8 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t0 5.17836
R16780 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n9 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n4 2.13175
R16781 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n3 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n2 1.11873
R16782 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n11 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n5 2.13275
R16783 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n1 0.0786548
R16784 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n14 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n1 2.13252
R16785 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n15 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n6 1.42979
R16786 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n7 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n18 1.42979
R16787 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n7 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n17 1.19668
R16788 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n0 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n1 1.11863
R16789 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n3 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n10 2.13252
R16790 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n13 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n12 1.80834
R16791 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n2 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n4 2.63066
R16792 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n0 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n5 2.51833
R16793 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n5 0.0794261
R16794 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n8 0.115328
R16795 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n13 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK 0.105738
R16796 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n4 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK 0.0794261
R16797 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n3 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK 0.0786538
R16798 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n7 0.19529
R16799 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n6 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK 0.19529
R16800 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n16 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n6 1.19668
R16801 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n16 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n0 1.01264
R16802 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n17 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n2 0.890034
R16803 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n2 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t9 36.935
R16804 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n6 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t8 31.4332
R16805 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n8 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t12 31.4332
R16806 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n3 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t4 31.4332
R16807 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n5 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t5 30.5752
R16808 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n5 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t6 21.7814
R16809 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n2 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t3 18.1962
R16810 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n6 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t7 15.3826
R16811 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n8 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t11 15.3826
R16812 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n3 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t10 15.3826
R16813 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t2 7.09905
R16814 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n8 6.86658
R16815 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n6 6.86658
R16816 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n3 6.86029
R16817 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n9 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2 5.61266
R16818 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n4 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2 5.01077
R16819 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n1 3.25053
R16820 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n7 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2 3.01024
R16821 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n9 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n7 2.84996
R16822 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n10 2.34645
R16823 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n1 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t0 2.2755
R16824 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n1 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n0 2.2755
R16825 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n2 2.13459
R16826 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n5 1.80883
R16827 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n7 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2 1.67882
R16828 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n10 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n4 1.5246
R16829 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n10 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n9 1.44585
R16830 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n4 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2 1.12067
R16831 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n3 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t2 37.1981
R16832 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n5 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t4 31.4332
R16833 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n4 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t6 30.4613
R16834 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n4 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t3 24.7562
R16835 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n3 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t5 17.6611
R16836 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n5 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t7 15.3826
R16837 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n0 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 12.0716
R16838 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n5 7.62076
R16839 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n6 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 6.09789
R16840 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n7 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n2 2.99416
R16841 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n2 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t0 2.2755
R16842 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n2 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n1 2.2755
R16843 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n7 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n6 2.2505
R16844 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n0 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 2.24788
R16845 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n6 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n0 1.94903
R16846 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n4 1.81638
R16847 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n3 1.43706
R16848 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n7 0.4325
R16849 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.n2 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.t3 36.935
R16850 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.n3 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.t5 31.4332
R16851 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.n5 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.t7 29.8135
R16852 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.n5 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.t4 27.8352
R16853 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.n2 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.t6 18.1962
R16854 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.n3 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.t8 15.3826
R16855 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.t2 7.09905
R16856 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.n3 6.86029
R16857 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.n4 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 5.01077
R16858 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.n6 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 3.41843
R16859 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.n1 3.25053
R16860 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.n1 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.t0 2.2755
R16861 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.n1 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.n0 2.2755
R16862 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.n6 2.2505
R16863 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.n2 2.13459
R16864 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.n5 1.74998
R16865 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.n6 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.n4 1.50381
R16866 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.n4 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 1.12067
R16867 CLK.n59 CLK.t91 36.935
R16868 CLK.n54 CLK.t41 36.935
R16869 CLK.n74 CLK.t27 36.935
R16870 CLK.n66 CLK.t14 36.935
R16871 CLK.n99 CLK.t87 36.935
R16872 CLK.n94 CLK.t25 36.935
R16873 CLK.n9 CLK.t92 36.935
R16874 CLK.n2 CLK.t76 36.935
R16875 CLK.n32 CLK.t70 36.935
R16876 CLK.n40 CLK.t29 36.935
R16877 CLK.n278 CLK.t90 36.935
R16878 CLK.n273 CLK.t75 36.935
R16879 CLK.n293 CLK.t69 36.935
R16880 CLK.n285 CLK.t57 36.935
R16881 CLK.n194 CLK.t16 36.935
R16882 CLK.n188 CLK.t53 36.935
R16883 CLK.n208 CLK.t24 36.935
R16884 CLK.n202 CLK.t5 36.935
R16885 CLK.n226 CLK.t48 36.935
R16886 CLK.n220 CLK.t4 36.935
R16887 CLK.n250 CLK.t68 36.935
R16888 CLK.n244 CLK.t40 36.935
R16889 CLK.n237 CLK.t22 36.935
R16890 CLK.n151 CLK.t60 36.935
R16891 CLK.n145 CLK.t32 36.935
R16892 CLK.n166 CLK.t0 36.935
R16893 CLK.n159 CLK.t62 36.935
R16894 CLK.n118 CLK.t50 36.935
R16895 CLK.n124 CLK.t88 36.935
R16896 CLK.n110 CLK.t79 31.528
R16897 CLK.n156 CLK.t63 30.6315
R16898 CLK.n71 CLK.t47 30.5752
R16899 CLK.n290 CLK.t36 30.5752
R16900 CLK.n26 CLK.t6 25.5364
R16901 CLK.n213 CLK.t59 25.5364
R16902 CLK.n231 CLK.t56 25.5364
R16903 CLK.n255 CLK.t80 25.5361
R16904 CLK.n262 CLK.t85 25.5361
R16905 CLK.n173 CLK.t19 25.5361
R16906 CLK.n180 CLK.t46 25.5361
R16907 CLK.n81 CLK.t77 25.4744
R16908 CLK.n105 CLK.t67 25.4744
R16909 CLK.n300 CLK.t38 25.4744
R16910 CLK.n307 CLK.t55 25.4744
R16911 CLK.n115 CLK.t81 25.4744
R16912 CLK.n50 CLK.t64 25.4742
R16913 CLK.n18 CLK.t42 25.2177
R16914 CLK.n71 CLK.t54 21.7814
R16915 CLK.n290 CLK.t44 21.7814
R16916 CLK.n156 CLK.t35 21.7275
R16917 CLK.n59 CLK.t33 18.1962
R16918 CLK.n54 CLK.t18 18.1962
R16919 CLK.n74 CLK.t71 18.1962
R16920 CLK.n66 CLK.t82 18.1962
R16921 CLK.n99 CLK.t15 18.1962
R16922 CLK.n94 CLK.t20 18.1962
R16923 CLK.n9 CLK.t78 18.1962
R16924 CLK.n2 CLK.t65 18.1962
R16925 CLK.n32 CLK.t83 18.1962
R16926 CLK.n40 CLK.t30 18.1962
R16927 CLK.n278 CLK.t21 18.1962
R16928 CLK.n273 CLK.t13 18.1962
R16929 CLK.n293 CLK.t8 18.1962
R16930 CLK.n285 CLK.t2 18.1962
R16931 CLK.n194 CLK.t49 18.1962
R16932 CLK.n188 CLK.t3 18.1962
R16933 CLK.n208 CLK.t61 18.1962
R16934 CLK.n202 CLK.t37 18.1962
R16935 CLK.n226 CLK.t58 18.1962
R16936 CLK.n220 CLK.t34 18.1962
R16937 CLK.n250 CLK.t10 18.1962
R16938 CLK.n244 CLK.t86 18.1962
R16939 CLK.n237 CLK.t52 18.1962
R16940 CLK.n151 CLK.t72 18.1962
R16941 CLK.n145 CLK.t28 18.1962
R16942 CLK.n166 CLK.t9 18.1962
R16943 CLK.n159 CLK.t31 18.1962
R16944 CLK.n118 CLK.t84 18.1962
R16945 CLK.n124 CLK.t17 18.1962
R16946 CLK.n110 CLK.t7 15.3826
R16947 CLK.n50 CLK.t89 14.142
R16948 CLK.n81 CLK.t45 14.1417
R16949 CLK.n105 CLK.t74 14.1417
R16950 CLK.n300 CLK.t1 14.1417
R16951 CLK.n307 CLK.t12 14.1417
R16952 CLK.n115 CLK.t66 14.1417
R16953 CLK.n26 CLK.t93 14.0749
R16954 CLK.n213 CLK.t26 14.0749
R16955 CLK.n231 CLK.t23 14.0749
R16956 CLK.n255 CLK.t39 14.0734
R16957 CLK.n262 CLK.t43 14.0734
R16958 CLK.n173 CLK.t73 14.0734
R16959 CLK.n180 CLK.t11 14.0734
R16960 CLK.n19 CLK.t51 13.6765
R16961 CLK.n47 CLK.n46 8.843
R16962 CLK.n111 CLK.n110 7.62171
R16963 CLK.n73 CLK.n72 7.41483
R16964 CLK.n292 CLK.n291 7.41483
R16965 CLK.n164 CLK.n157 7.41437
R16966 CLK.n90 CLK 6.87797
R16967 CLK.n269 CLK.n268 6.74647
R16968 CLK.n142 CLK.n141 6.61208
R16969 CLK.n312 CLK.n311 6.5934
R16970 CLK.n113 CLK.n112 6.33303
R16971 CLK.n184 CLK 6.14196
R16972 CLK.n269 CLK.n184 6.04302
R16973 CLK.n260 CLK 5.77906
R16974 CLK.n109 CLK 5.51417
R16975 CLK.n178 CLK.n177 5.37352
R16976 CLK.n86 CLK.n85 5.37091
R16977 CLK.n305 CLK.n304 5.37091
R16978 CLK.n311 CLK 5.24048
R16979 CLK.n264 CLK.n261 5.11659
R16980 CLK.n112 CLK.n111 5.0581
R16981 CLK.n47 CLK.n24 4.73335
R16982 CLK.n268 CLK.n266 4.56336
R16983 CLK.n56 CLK.n53 4.5005
R16984 CLK.n58 CLK.n57 4.5005
R16985 CLK.n62 CLK.n60 4.5005
R16986 CLK.n62 CLK.n61 4.5005
R16987 CLK.n68 CLK.n65 4.5005
R16988 CLK.n70 CLK.n69 4.5005
R16989 CLK.n77 CLK.n75 4.5005
R16990 CLK.n77 CLK.n76 4.5005
R16991 CLK.n80 CLK.n79 4.5005
R16992 CLK.n82 CLK.n79 4.5005
R16993 CLK.n89 CLK.n88 4.5005
R16994 CLK.n88 CLK.n51 4.5005
R16995 CLK.n96 CLK.n93 4.5005
R16996 CLK.n98 CLK.n97 4.5005
R16997 CLK.n102 CLK.n100 4.5005
R16998 CLK.n102 CLK.n101 4.5005
R16999 CLK.n108 CLK.n107 4.5005
R17000 CLK.n107 CLK.n106 4.5005
R17001 CLK.n23 CLK.n17 4.5005
R17002 CLK.n23 CLK.n22 4.5005
R17003 CLK.n16 CLK.n14 4.5005
R17004 CLK.n16 CLK.n15 4.5005
R17005 CLK.n275 CLK.n272 4.5005
R17006 CLK.n277 CLK.n276 4.5005
R17007 CLK.n281 CLK.n279 4.5005
R17008 CLK.n281 CLK.n280 4.5005
R17009 CLK.n287 CLK.n284 4.5005
R17010 CLK.n289 CLK.n288 4.5005
R17011 CLK.n296 CLK.n294 4.5005
R17012 CLK.n296 CLK.n295 4.5005
R17013 CLK.n299 CLK.n298 4.5005
R17014 CLK.n301 CLK.n298 4.5005
R17015 CLK.n310 CLK.n309 4.5005
R17016 CLK.n309 CLK.n308 4.5005
R17017 CLK.n190 CLK.n187 4.5005
R17018 CLK.n190 CLK.n189 4.5005
R17019 CLK.n193 CLK.n192 4.5005
R17020 CLK.n195 CLK.n192 4.5005
R17021 CLK.n204 CLK.n201 4.5005
R17022 CLK.n204 CLK.n203 4.5005
R17023 CLK.n207 CLK.n206 4.5005
R17024 CLK.n209 CLK.n206 4.5005
R17025 CLK.n216 CLK.n215 4.5005
R17026 CLK.n215 CLK.n214 4.5005
R17027 CLK.n222 CLK.n219 4.5005
R17028 CLK.n222 CLK.n221 4.5005
R17029 CLK.n225 CLK.n224 4.5005
R17030 CLK.n227 CLK.n224 4.5005
R17031 CLK.n234 CLK.n233 4.5005
R17032 CLK.n233 CLK.n232 4.5005
R17033 CLK.n246 CLK.n243 4.5005
R17034 CLK.n246 CLK.n245 4.5005
R17035 CLK.n249 CLK.n248 4.5005
R17036 CLK.n251 CLK.n248 4.5005
R17037 CLK.n258 CLK.n257 4.5005
R17038 CLK.n257 CLK.n256 4.5005
R17039 CLK.n238 CLK.n235 4.5005
R17040 CLK.n265 CLK.n264 4.5005
R17041 CLK.n264 CLK.n263 4.5005
R17042 CLK.n148 CLK.n146 4.5005
R17043 CLK.n148 CLK.n147 4.5005
R17044 CLK.n152 CLK.n150 4.5005
R17045 CLK.n153 CLK.n150 4.5005
R17046 CLK.n162 CLK.n160 4.5005
R17047 CLK.n162 CLK.n161 4.5005
R17048 CLK.n167 CLK.n165 4.5005
R17049 CLK.n168 CLK.n165 4.5005
R17050 CLK.n172 CLK.n171 4.5005
R17051 CLK.n174 CLK.n171 4.5005
R17052 CLK.n182 CLK.n181 4.5005
R17053 CLK.n183 CLK.n182 4.5005
R17054 CLK.n313 CLK.n109 4.44251
R17055 CLK.n261 CLK 4.43149
R17056 CLK.n312 CLK.n142 4.25721
R17057 CLK.n266 CLK 4.10231
R17058 CLK.n259 CLK.n240 4.05348
R17059 CLK.n20 CLK.n19 3.5993
R17060 CLK.n260 CLK.n259 3.5258
R17061 CLK.n259 CLK 2.3355
R17062 CLK CLK.n0 2.27847
R17063 CLK.n267 CLK 2.27103
R17064 CLK.n136 CLK.n135 2.2567
R17065 CLK.n63 CLK.n52 2.25107
R17066 CLK.n78 CLK.n64 2.25107
R17067 CLK.n103 CLK.n92 2.25107
R17068 CLK.n12 CLK.n11 2.25107
R17069 CLK.n282 CLK.n271 2.25107
R17070 CLK.n297 CLK.n283 2.25107
R17071 CLK.n197 CLK.n196 2.25107
R17072 CLK.n211 CLK.n210 2.25107
R17073 CLK.n229 CLK.n228 2.25107
R17074 CLK.n253 CLK.n252 2.25107
R17075 CLK.n155 CLK.n154 2.25107
R17076 CLK.n170 CLK.n169 2.25107
R17077 CLK.n129 CLK.n121 2.25107
R17078 CLK.n43 CLK.n42 2.2505
R17079 CLK.n48 CLK.n47 2.2505
R17080 CLK.n236 CLK.n235 2.24763
R17081 CLK.n240 CLK.n239 2.2455
R17082 CLK.n176 CLK.n175 2.24385
R17083 CLK.n179 CLK.n143 2.24385
R17084 CLK.n84 CLK.n83 2.24352
R17085 CLK.n87 CLK.n49 2.24352
R17086 CLK.n303 CLK.n302 2.24352
R17087 CLK.n306 CLK.n270 2.24352
R17088 CLK.n130 CLK.n117 2.24319
R17089 CLK.n212 CLK.n199 2.24235
R17090 CLK.n230 CLK.n217 2.24235
R17091 CLK.n254 CLK.n241 2.24235
R17092 CLK.n198 CLK.n185 2.24235
R17093 CLK.n30 CLK.n29 2.24235
R17094 CLK.n104 CLK.n91 2.24196
R17095 CLK.n67 CLK.n66 2.12464
R17096 CLK.n55 CLK.n54 2.12444
R17097 CLK.n95 CLK.n94 2.12444
R17098 CLK.n274 CLK.n273 2.12444
R17099 CLK.n286 CLK.n285 2.12444
R17100 CLK.n125 CLK.n124 2.12444
R17101 CLK.n238 CLK.n237 2.12226
R17102 CLK.n152 CLK.n151 2.12207
R17103 CLK.n167 CLK.n166 2.12207
R17104 CLK.n60 CLK.n59 2.12188
R17105 CLK.n75 CLK.n74 2.12188
R17106 CLK.n100 CLK.n99 2.12188
R17107 CLK.n279 CLK.n278 2.12188
R17108 CLK.n294 CLK.n293 2.12188
R17109 CLK.n146 CLK.n145 2.12188
R17110 CLK.n160 CLK.n159 2.12188
R17111 CLK.n119 CLK.n118 2.12188
R17112 CLK.n3 CLK.n2 2.12175
R17113 CLK.n33 CLK.n32 2.12175
R17114 CLK.n189 CLK.n188 2.12175
R17115 CLK.n203 CLK.n202 2.12175
R17116 CLK.n221 CLK.n220 2.12175
R17117 CLK.n245 CLK.n244 2.12175
R17118 CLK.n10 CLK.n9 2.12075
R17119 CLK.n41 CLK.n40 2.12075
R17120 CLK.n195 CLK.n194 2.12075
R17121 CLK.n209 CLK.n208 2.12075
R17122 CLK.n227 CLK.n226 2.12075
R17123 CLK.n251 CLK.n250 2.12075
R17124 CLK.n90 CLK.n48 1.8876
R17125 CLK.n72 CLK.n71 1.80883
R17126 CLK.n291 CLK.n290 1.80883
R17127 CLK.n157 CLK.n156 1.80496
R17128 CLK.n7 CLK.n6 1.74297
R17129 CLK.n192 CLK.n191 1.74297
R17130 CLK.n206 CLK.n205 1.74297
R17131 CLK.n224 CLK.n223 1.74297
R17132 CLK.n248 CLK.n247 1.74297
R17133 CLK.n150 CLK.n149 1.74297
R17134 CLK.n62 CLK.n58 1.71671
R17135 CLK.n102 CLK.n98 1.71671
R17136 CLK.n281 CLK.n277 1.71671
R17137 CLK.n128 CLK.n127 1.71671
R17138 CLK.n261 CLK.n260 1.62556
R17139 CLK.n164 CLK.n163 1.62464
R17140 CLK.n73 CLK.n70 1.59838
R17141 CLK.n292 CLK.n289 1.59838
R17142 CLK.n55 CLK.n53 1.50503
R17143 CLK.n67 CLK.n65 1.50503
R17144 CLK.n95 CLK.n93 1.50503
R17145 CLK.n274 CLK.n272 1.50503
R17146 CLK.n286 CLK.n284 1.50503
R17147 CLK.n126 CLK.n125 1.50503
R17148 CLK.n138 CLK.n136 1.50161
R17149 CLK.n6 CLK.n4 1.49778
R17150 CLK.n191 CLK.n186 1.49778
R17151 CLK.n205 CLK.n200 1.49778
R17152 CLK.n223 CLK.n218 1.49778
R17153 CLK.n247 CLK.n242 1.49778
R17154 CLK.n149 CLK.n144 1.49778
R17155 CLK.n163 CLK.n158 1.49778
R17156 CLK.n36 CLK.n34 1.49774
R17157 CLK.n256 CLK.n255 1.42775
R17158 CLK.n263 CLK.n262 1.42775
R17159 CLK.n174 CLK.n173 1.42775
R17160 CLK.n181 CLK.n180 1.42775
R17161 CLK.n27 CLK.n26 1.42706
R17162 CLK.n214 CLK.n213 1.42706
R17163 CLK.n232 CLK.n231 1.42706
R17164 CLK.n51 CLK.n50 1.42126
R17165 CLK.n82 CLK.n81 1.42118
R17166 CLK.n106 CLK.n105 1.42118
R17167 CLK.n301 CLK.n300 1.42118
R17168 CLK.n308 CLK.n307 1.42118
R17169 CLK.n116 CLK.n115 1.42118
R17170 CLK.n109 CLK.n90 1.40597
R17171 CLK.n141 CLK.n140 1.32117
R17172 CLK.n313 CLK.n312 1.23194
R17173 CLK.n198 CLK.n197 0.97145
R17174 CLK.n212 CLK.n211 0.97145
R17175 CLK.n230 CLK.n229 0.97145
R17176 CLK.n254 CLK.n253 0.97145
R17177 CLK.n104 CLK.n103 0.969075
R17178 CLK.n130 CLK.n129 0.964895
R17179 CLK.n46 CLK.n45 0.953968
R17180 CLK.n13 CLK.n12 0.930887
R17181 CLK.n268 CLK.n267 0.899626
R17182 CLK.n86 CLK.n63 0.882596
R17183 CLK.n85 CLK.n78 0.882596
R17184 CLK.n305 CLK.n282 0.882596
R17185 CLK.n304 CLK.n297 0.882596
R17186 CLK.n178 CLK.n155 0.882596
R17187 CLK.n177 CLK.n170 0.882596
R17188 CLK.n37 CLK.n36 0.879852
R17189 CLK.n45 CLK.n37 0.843227
R17190 CLK.n311 CLK.n269 0.823767
R17191 CLK.n19 CLK.n18 0.804397
R17192 CLK CLK.n313 0.7853
R17193 CLK.n80 CLK 0.1605
R17194 CLK CLK.n108 0.1605
R17195 CLK.n299 CLK 0.1605
R17196 CLK CLK.n216 0.1605
R17197 CLK CLK.n234 0.1605
R17198 CLK CLK.n258 0.1605
R17199 CLK CLK.n265 0.1605
R17200 CLK.n172 CLK 0.1605
R17201 CLK.n141 CLK.n113 0.158593
R17202 CLK.n28 CLK 0.1355
R17203 CLK.n77 CLK.n73 0.118826
R17204 CLK.n296 CLK.n292 0.118826
R17205 CLK.n165 CLK.n164 0.118826
R17206 CLK.n72 CLK 0.108371
R17207 CLK.n291 CLK 0.108371
R17208 CLK.n157 CLK 0.107668
R17209 CLK.n135 CLK.n134 0.09875
R17210 CLK.n17 CLK 0.0950833
R17211 CLK.n43 CLK.n38 0.0901918
R17212 CLK.n85 CLK.n84 0.0733415
R17213 CLK.n87 CLK.n86 0.0733415
R17214 CLK.n304 CLK.n303 0.0733415
R17215 CLK.n306 CLK.n305 0.0733415
R17216 CLK.n177 CLK.n176 0.0726935
R17217 CLK.n179 CLK.n178 0.0726935
R17218 CLK CLK.n89 0.05925
R17219 CLK CLK.n310 0.05925
R17220 CLK CLK.n183 0.05925
R17221 CLK.n236 CLK 0.052998
R17222 CLK.n135 CLK 0.04775
R17223 CLK.n8 CLK 0.0473512
R17224 CLK.n1 CLK 0.0473512
R17225 CLK.n31 CLK 0.0473512
R17226 CLK.n39 CLK 0.0473512
R17227 CLK.n193 CLK 0.0473512
R17228 CLK.n187 CLK 0.0473512
R17229 CLK.n207 CLK 0.0473512
R17230 CLK.n201 CLK 0.0473512
R17231 CLK.n225 CLK 0.0473512
R17232 CLK.n219 CLK 0.0473512
R17233 CLK.n249 CLK 0.0473512
R17234 CLK.n243 CLK 0.0473512
R17235 CLK.n61 CLK 0.0457995
R17236 CLK.n56 CLK 0.0457995
R17237 CLK.n76 CLK 0.0457995
R17238 CLK.n68 CLK 0.0457995
R17239 CLK.n101 CLK 0.0457995
R17240 CLK.n96 CLK 0.0457995
R17241 CLK.n280 CLK 0.0457995
R17242 CLK.n275 CLK 0.0457995
R17243 CLK.n295 CLK 0.0457995
R17244 CLK.n287 CLK 0.0457995
R17245 CLK.n153 CLK 0.0457995
R17246 CLK.n147 CLK 0.0457995
R17247 CLK.n168 CLK 0.0457995
R17248 CLK.n161 CLK 0.0457995
R17249 CLK.n120 CLK 0.0457995
R17250 CLK.n122 CLK 0.0457995
R17251 CLK.n46 CLK.n30 0.0435648
R17252 CLK.n133 CLK.n132 0.0403734
R17253 CLK.n58 CLK.n53 0.0386356
R17254 CLK.n70 CLK.n65 0.0386356
R17255 CLK.n98 CLK.n93 0.0386356
R17256 CLK.n277 CLK.n272 0.0386356
R17257 CLK.n289 CLK.n284 0.0386356
R17258 CLK.n127 CLK.n126 0.0386356
R17259 CLK.n61 CLK.n52 0.0377414
R17260 CLK.n57 CLK.n56 0.0377414
R17261 CLK.n76 CLK.n64 0.0377414
R17262 CLK.n69 CLK.n68 0.0377414
R17263 CLK.n101 CLK.n92 0.0377414
R17264 CLK.n97 CLK.n96 0.0377414
R17265 CLK.n280 CLK.n271 0.0377414
R17266 CLK.n276 CLK.n275 0.0377414
R17267 CLK.n295 CLK.n283 0.0377414
R17268 CLK.n288 CLK.n287 0.0377414
R17269 CLK.n154 CLK.n153 0.0377414
R17270 CLK.n147 CLK.n144 0.0377414
R17271 CLK.n169 CLK.n168 0.0377414
R17272 CLK.n161 CLK.n158 0.0377414
R17273 CLK.n121 CLK.n120 0.0377414
R17274 CLK.n123 CLK.n122 0.0377414
R17275 CLK.n11 CLK.n8 0.0361897
R17276 CLK.n4 CLK.n1 0.0361897
R17277 CLK.n34 CLK.n31 0.0361897
R17278 CLK.n42 CLK.n39 0.0361897
R17279 CLK.n196 CLK.n193 0.0361897
R17280 CLK.n187 CLK.n186 0.0361897
R17281 CLK.n210 CLK.n207 0.0361897
R17282 CLK.n201 CLK.n200 0.0361897
R17283 CLK.n228 CLK.n225 0.0361897
R17284 CLK.n219 CLK.n218 0.0361897
R17285 CLK.n252 CLK.n249 0.0361897
R17286 CLK.n243 CLK.n242 0.0361897
R17287 CLK.n138 CLK.n137 0.034882
R17288 CLK.n132 CLK.n131 0.03466
R17289 CLK.n140 CLK.n139 0.0328596
R17290 CLK.n83 CLK.n80 0.03175
R17291 CLK.n89 CLK.n49 0.03175
R17292 CLK.n108 CLK.n91 0.03175
R17293 CLK.n29 CLK.n28 0.03175
R17294 CLK.n302 CLK.n299 0.03175
R17295 CLK.n310 CLK.n270 0.03175
R17296 CLK.n216 CLK.n199 0.03175
R17297 CLK.n234 CLK.n217 0.03175
R17298 CLK.n258 CLK.n241 0.03175
R17299 CLK.n265 CLK.n185 0.03175
R17300 CLK.n175 CLK.n172 0.03175
R17301 CLK.n183 CLK.n143 0.03175
R17302 CLK.n111 CLK 0.0316785
R17303 CLK.n16 CLK.n13 0.0309615
R17304 CLK.n215 CLK.n212 0.0246174
R17305 CLK.n233 CLK.n230 0.0246174
R17306 CLK.n257 CLK.n254 0.0246174
R17307 CLK.n264 CLK.n198 0.0246174
R17308 CLK.n30 CLK.n25 0.0246174
R17309 CLK.n107 CLK.n104 0.0238218
R17310 CLK.n239 CLK.n238 0.0210263
R17311 CLK.n131 CLK.n130 0.0207183
R17312 CLK.n176 CLK.n171 0.0205196
R17313 CLK.n182 CLK.n179 0.0205196
R17314 CLK.n84 CLK.n79 0.0198632
R17315 CLK.n88 CLK.n87 0.0198632
R17316 CLK.n303 CLK.n298 0.0198632
R17317 CLK.n309 CLK.n306 0.0198632
R17318 CLK.n239 CLK.n236 0.0183424
R17319 CLK.n36 CLK.n35 0.0139789
R17320 CLK.n6 CLK.n5 0.0131772
R17321 CLK.n191 CLK.n190 0.0131772
R17322 CLK.n205 CLK.n204 0.0131772
R17323 CLK.n223 CLK.n222 0.0131772
R17324 CLK.n247 CLK.n246 0.0131772
R17325 CLK.n149 CLK.n148 0.0131772
R17326 CLK.n163 CLK.n162 0.0131772
R17327 CLK.n240 CLK.n235 0.0128848
R17328 CLK.n136 CLK.n133 0.012347
R17329 CLK.n63 CLK.n62 0.0122182
R17330 CLK.n78 CLK.n77 0.0122182
R17331 CLK.n103 CLK.n102 0.0122182
R17332 CLK.n12 CLK.n7 0.0122182
R17333 CLK.n282 CLK.n281 0.0122182
R17334 CLK.n297 CLK.n296 0.0122182
R17335 CLK.n197 CLK.n192 0.0122182
R17336 CLK.n211 CLK.n206 0.0122182
R17337 CLK.n229 CLK.n224 0.0122182
R17338 CLK.n253 CLK.n248 0.0122182
R17339 CLK.n155 CLK.n150 0.0122182
R17340 CLK.n170 CLK.n165 0.0122182
R17341 CLK.n129 CLK.n128 0.0122182
R17342 CLK.n112 CLK 0.0095
R17343 CLK.n45 CLK.n44 0.00913014
R17344 CLK.n24 CLK.n16 0.00542459
R17345 CLK.n11 CLK.n10 0.00515517
R17346 CLK.n4 CLK.n3 0.00515517
R17347 CLK.n34 CLK.n33 0.00515517
R17348 CLK.n42 CLK.n41 0.00515517
R17349 CLK.n196 CLK.n195 0.00515517
R17350 CLK.n189 CLK.n186 0.00515517
R17351 CLK.n210 CLK.n209 0.00515517
R17352 CLK.n203 CLK.n200 0.00515517
R17353 CLK.n228 CLK.n227 0.00515517
R17354 CLK.n221 CLK.n218 0.00515517
R17355 CLK.n252 CLK.n251 0.00515517
R17356 CLK.n245 CLK.n242 0.00515517
R17357 CLK.n113 CLK 0.00469786
R17358 CLK.n44 CLK.n43 0.00419863
R17359 CLK.n60 CLK.n52 0.00360345
R17360 CLK.n75 CLK.n64 0.00360345
R17361 CLK.n100 CLK.n92 0.00360345
R17362 CLK.n279 CLK.n271 0.00360345
R17363 CLK.n294 CLK.n283 0.00360345
R17364 CLK.n154 CLK.n152 0.00360345
R17365 CLK.n146 CLK.n144 0.00360345
R17366 CLK.n169 CLK.n167 0.00360345
R17367 CLK.n160 CLK.n158 0.00360345
R17368 CLK.n121 CLK.n119 0.00360345
R17369 CLK.n22 CLK.n20 0.003
R17370 CLK.n139 CLK.n114 0.00286842
R17371 CLK.n24 CLK.n23 0.00210846
R17372 CLK.n57 CLK.n55 0.00203726
R17373 CLK.n69 CLK.n67 0.00203726
R17374 CLK.n97 CLK.n95 0.00203726
R17375 CLK.n276 CLK.n274 0.00203726
R17376 CLK.n288 CLK.n286 0.00203726
R17377 CLK.n125 CLK.n123 0.00203726
R17378 CLK.n83 CLK.n82 0.00175
R17379 CLK.n51 CLK.n49 0.00175
R17380 CLK.n106 CLK.n91 0.00175
R17381 CLK.n29 CLK.n27 0.00175
R17382 CLK.n302 CLK.n301 0.00175
R17383 CLK.n308 CLK.n270 0.00175
R17384 CLK.n214 CLK.n199 0.00175
R17385 CLK.n232 CLK.n217 0.00175
R17386 CLK.n256 CLK.n241 0.00175
R17387 CLK.n263 CLK.n185 0.00175
R17388 CLK.n175 CLK.n174 0.00175
R17389 CLK.n181 CLK.n143 0.00175
R17390 CLK.n117 CLK.n116 0.00175
R17391 CLK.n139 CLK.n138 0.00151124
R17392 CLK.n22 CLK.n21 0.00133333
R17393 CLK.n142 CLK 0.00110798
R17394 CLK CLK.n266 0.000959184
R17395 CLK.n267 CLK 0.000959184
R17396 Vdiv100.n2 Vdiv100.t4 31.528
R17397 Vdiv100.n2 Vdiv100.t5 15.3826
R17398 Vdiv100.n9 Vdiv100 9.77396
R17399 Vdiv100.n7 Vdiv100.t2 9.28805
R17400 Vdiv100 Vdiv100.n2 7.62076
R17401 Vdiv100.n6 Vdiv100.n5 6.01414
R17402 Vdiv100.n6 Vdiv100.t0 6.01414
R17403 Vdiv100 Vdiv100.n8 5.89054
R17404 Vdiv100 Vdiv100.n14 4.53253
R17405 Vdiv100.n8 Vdiv100.t3 3.87536
R17406 Vdiv100.n7 Vdiv100.n6 3.74829
R17407 Vdiv100.n4 Vdiv100.n1 1.5005
R17408 Vdiv100.n12 Vdiv100.n11 1.5005
R17409 Vdiv100.n0 Vdiv100 0.0664402
R17410 Vdiv100.n8 Vdiv100.n7 0.0409348
R17411 Vdiv100.n1 Vdiv100.n0 0.0386356
R17412 Vdiv100.n10 Vdiv100.n9 0.0341364
R17413 Vdiv100.n4 Vdiv100.n3 0.0232273
R17414 Vdiv100.n14 Vdiv100.n13 0.0232273
R17415 Vdiv100 Vdiv100.n1 0.0127034
R17416 Vdiv100.n13 Vdiv100.n12 0.00504545
R17417 Vdiv100.n12 Vdiv100.n4 0.00322727
R17418 Vdiv100.n11 Vdiv100.n10 0.00322727
R17419 Vdiv100.n8 Vdiv100 0.0031087
R17420 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n17 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t14 36.935
R17421 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n18 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t15 36.935
R17422 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n12 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t9 36.935
R17423 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n19 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t5 31.4332
R17424 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n14 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t8 31.4332
R17425 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n20 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t6 30.9379
R17426 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n22 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t13 25.4744
R17427 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n20 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t7 21.6422
R17428 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n17 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t12 18.1962
R17429 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n18 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t16 18.1962
R17430 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n12 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t10 18.1962
R17431 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n19 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t4 15.3826
R17432 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n14 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t11 15.3826
R17433 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n22 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t3 14.1417
R17434 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n11 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t1 7.09905
R17435 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n15 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n14 6.86029
R17436 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n16 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n13 5.01077
R17437 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n2 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n4 0.0219501
R17438 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n1 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n0 0.0360559
R17439 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n19 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 5.69501
R17440 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n4 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n1 2.23369
R17441 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n2 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n0 1.11499
R17442 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n23 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n8 2.2429
R17443 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n8 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n7 0.0171915
R17444 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n11 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n10 3.25053
R17445 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n10 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t2 2.2755
R17446 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n10 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n9 2.2755
R17447 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n25 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n24 2.2505
R17448 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n7 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n6 2.24196
R17449 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n13 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n12 2.13459
R17450 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n3 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n20 2.13074
R17451 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n4 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n17 2.12093
R17452 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n1 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n5 2.64237
R17453 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n0 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n21 4.95192
R17454 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n21 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 4.19069
R17455 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n24 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n16 1.52773
R17456 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n18 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n5 2.13281
R17457 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n7 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n22 1.42118
R17458 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n16 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n15 1.12067
R17459 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n6 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n0 0.960138
R17460 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n23 0.646487
R17461 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n8 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 0.187192
R17462 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n25 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n11 0.0905
R17463 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n15 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 0.0857632
R17464 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n25 0.0834687
R17465 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n13 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 0.0800273
R17466 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n3 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 0.0980715
R17467 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n2 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 0.0672526
R17468 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n5 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 0.0771461
R17469 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n24 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 0.0322045
R17470 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n23 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n6 0.0238218
R17471 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n21 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n3 2.08419
R17472 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.n3 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.t3 36.935
R17473 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.n4 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.t6 31.4332
R17474 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.n2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.t8 29.8635
R17475 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.n2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.t5 27.7543
R17476 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.n3 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.t7 18.1962
R17477 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.n4 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.t4 15.3826
R17478 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.t0 7.09905
R17479 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.n4 6.86134
R17480 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.n5 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 5.0096
R17481 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.n6 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 3.41823
R17482 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.n1 3.25226
R17483 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.n1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.t2 2.2755
R17484 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.n1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.n0 2.2755
R17485 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.n6 2.2505
R17486 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.n3 2.13479
R17487 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.n2 1.7371
R17488 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.n6 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.n5 1.50498
R17489 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.n5 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 1.12056
R17490 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n19 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t7 36.935
R17491 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n18 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t9 36.935
R17492 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n22 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t16 36.935
R17493 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n21 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t14 36.935
R17494 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n13 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t18 36.935
R17495 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n15 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t13 31.4332
R17496 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n24 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t19 30.6613
R17497 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n20 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t3 25.4744
R17498 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n26 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t12 25.4744
R17499 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n24 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t20 21.6718
R17500 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n19 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t6 18.1962
R17501 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n18 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t8 18.1962
R17502 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n22 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t15 18.1962
R17503 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n21 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t4 18.1962
R17504 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n13 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t11 18.1962
R17505 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n15 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t5 15.3826
R17506 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n26 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t17 14.1417
R17507 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n20 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t10 14.1417
R17508 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n0 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n25 9.9005
R17509 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n12 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t1 7.09905
R17510 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n16 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n15 6.86029
R17511 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n17 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n14 5.01077
R17512 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n2 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n3 1.11863
R17513 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n4 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n5 1.11863
R17514 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n20 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n9 1.42995
R17515 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n0 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n1 1.11781
R17516 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n12 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n11 3.25053
R17517 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n11 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t2 2.2755
R17518 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n11 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n10 2.2755
R17519 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n28 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n27 2.2505
R17520 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n23 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n9 1.16587
R17521 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n14 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n13 2.13459
R17522 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n3 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n19 2.13265
R17523 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n5 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n22 2.13265
R17524 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n2 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n7 2.63776
R17525 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n4 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n8 2.63776
R17526 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n27 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n17 1.52773
R17527 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n18 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n7 2.13261
R17528 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n21 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n8 2.13281
R17529 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n1 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n26 1.42999
R17530 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n6 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n24 1.41101
R17531 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n17 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n16 1.12067
R17532 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n25 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n23 0.286289
R17533 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n1 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 0.196008
R17534 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n9 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 0.196051
R17535 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n28 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n12 0.0905
R17536 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n16 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 0.0857632
R17537 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n28 0.0834687
R17538 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n6 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 0.104828
R17539 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n14 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 0.0800273
R17540 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n8 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 0.0771461
R17541 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n7 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 0.0771461
R17542 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n5 0.077103
R17543 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n3 0.077103
R17544 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n27 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 0.0289903
R17545 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n25 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n6 7.13895
R17546 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n0 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n2 1.18681
R17547 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n23 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n4 0.938524
R17548 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n0 0.680217
R17549 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n4 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t5 37.1986
R17550 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n3 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t3 31.528
R17551 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n2 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t6 30.5184
R17552 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n2 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t7 24.7029
R17553 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n4 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t4 17.6614
R17554 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n3 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t8 15.3826
R17555 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n0 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 12.0843
R17556 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n0 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n3 9.86691
R17557 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n5 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 6.09789
R17558 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n7 2.99416
R17559 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n7 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t2 2.2755
R17560 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n7 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n6 2.2755
R17561 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n5 2.2505
R17562 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n0 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 2.24173
R17563 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n5 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n0 1.93723
R17564 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n2 1.81225
R17565 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n4 1.43709
R17566 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n1 0.281955
R17567 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n14 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t15 36.935
R17568 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n9 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t5 36.935
R17569 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n20 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t10 36.935
R17570 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n26 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t16 31.4332
R17571 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n23 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t7 30.9379
R17572 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n22 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t11 30.9379
R17573 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n6 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t13 25.4744
R17574 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n23 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t3 21.6422
R17575 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n22 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t8 21.6422
R17576 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n14 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t4 18.1962
R17577 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n9 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t9 18.1962
R17578 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n20 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t14 18.1962
R17579 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n26 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t6 15.3826
R17580 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n6 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t12 14.1417
R17581 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n4 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t0 7.09905
R17582 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n27 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n26 6.86029
R17583 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n24 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 6.54296
R17584 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n25 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n24 4.54543
R17585 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n0 1.50092
R17586 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n11 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n8 4.5005
R17587 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n13 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n12 4.5005
R17588 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n17 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n15 4.5005
R17589 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n17 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n16 4.5005
R17590 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n19 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n5 4.5005
R17591 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n23 4.11094
R17592 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n22 4.11094
R17593 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n28 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n25 3.5302
R17594 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n4 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n3 3.25053
R17595 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n3 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t2 2.2755
R17596 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n3 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n2 2.2755
R17597 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n29 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 2.25167
R17598 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n18 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n7 2.25107
R17599 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n21 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n20 2.13459
R17600 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n10 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n9 2.12444
R17601 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n15 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n14 2.12188
R17602 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n17 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n13 1.71671
R17603 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n28 1.52539
R17604 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n10 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n8 1.50503
R17605 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n25 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n21 1.37844
R17606 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n28 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n27 1.12067
R17607 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n0 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n18 0.932217
R17608 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n24 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 0.485557
R17609 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n5 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 0.1705
R17610 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n29 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n4 0.0905
R17611 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n27 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 0.0857632
R17612 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n29 0.0834687
R17613 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n21 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 0.0800273
R17614 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n16 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 0.0457995
R17615 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n11 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 0.0457995
R17616 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n13 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n8 0.0386356
R17617 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n16 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n7 0.0377414
R17618 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n12 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n11 0.0377414
R17619 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n19 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n0 0.0322517
R17620 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n5 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n1 0.0326665
R17621 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n18 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n17 0.0122182
R17622 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n15 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n7 0.00360345
R17623 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n12 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n10 0.00203726
R17624 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n6 1.42251
R17625 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n19 0.338856
R17626 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n5 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t4 37.1984
R17627 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n4 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t3 31.4332
R17628 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n3 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t2 30.5184
R17629 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n3 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t7 24.7029
R17630 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n5 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t5 17.6618
R17631 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n4 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t6 15.3826
R17632 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n0 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 12.0839
R17633 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n0 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n4 9.86691
R17634 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n6 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 6.09789
R17635 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n7 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n2 2.99416
R17636 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t0 2.2755
R17637 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n1 2.2755
R17638 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n7 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n6 2.2505
R17639 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n0 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 2.24134
R17640 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n6 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n0 1.93723
R17641 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n3 1.81224
R17642 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n5 1.43718
R17643 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n7 0.4325
R17644 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n2 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t10 36.935
R17645 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n6 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t5 31.4332
R17646 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n8 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t4 31.4332
R17647 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n3 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t8 31.4332
R17648 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n5 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t6 30.5752
R17649 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n5 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t11 21.7814
R17650 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n2 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t9 18.1962
R17651 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n6 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t3 15.3826
R17652 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n8 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t12 15.3826
R17653 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n3 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t7 15.3826
R17654 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t2 7.09905
R17655 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n8 6.86658
R17656 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n6 6.86658
R17657 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n3 6.86029
R17658 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n9 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2 5.61266
R17659 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n4 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2 5.01077
R17660 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n1 3.25053
R17661 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n7 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2 3.01024
R17662 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n9 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n7 2.84996
R17663 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n10 2.34645
R17664 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n1 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t0 2.2755
R17665 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n1 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n0 2.2755
R17666 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n2 2.13459
R17667 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n5 1.80883
R17668 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n7 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2 1.67882
R17669 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n10 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n4 1.5246
R17670 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n10 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n9 1.44585
R17671 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n4 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2 1.12067
R17672 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.n2 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.t6 36.935
R17673 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.n3 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.t7 31.4332
R17674 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.n5 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.t3 29.8135
R17675 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.n5 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.t8 27.8352
R17676 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.n2 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.t4 18.1962
R17677 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.n3 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.t5 15.3826
R17678 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.t0 7.09905
R17679 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.n3 6.86029
R17680 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.n4 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 5.01077
R17681 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.n6 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 3.41843
R17682 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.n1 3.25053
R17683 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.n1 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.t2 2.2755
R17684 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.n1 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.n0 2.2755
R17685 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.n6 2.2505
R17686 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.n2 2.13459
R17687 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.n5 1.74998
R17688 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.n6 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.n4 1.50381
R17689 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.n4 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 1.12067
R17690 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.n2 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.t8 36.935
R17691 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.n3 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.t7 31.4332
R17692 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.n5 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.t6 29.8135
R17693 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.n5 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.t5 27.8352
R17694 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.n2 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.t4 18.1962
R17695 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.n3 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.t3 15.3826
R17696 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.t2 7.09905
R17697 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.n3 6.86029
R17698 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.n4 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 5.01077
R17699 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.n6 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 3.41843
R17700 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.n1 3.25053
R17701 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.n1 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.t0 2.2755
R17702 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.n1 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.n0 2.2755
R17703 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.n6 2.2505
R17704 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.n2 2.13459
R17705 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.n5 1.74998
R17706 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.n6 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.n4 1.50381
R17707 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.n4 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 1.12067
R17708 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t4 37.1986
R17709 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t6 31.528
R17710 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n3 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t7 30.6315
R17711 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n3 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t8 24.5953
R17712 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t3 17.6614
R17713 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n4 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 17.0516
R17714 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t5 15.3826
R17715 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n1 7.62751
R17716 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n5 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n4 3.28711
R17717 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n7 2.99416
R17718 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n4 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 2.81128
R17719 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n5 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 2.67866
R17720 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n7 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t1 2.2755
R17721 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n7 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n6 2.2755
R17722 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n5 2.2505
R17723 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n3 1.80496
R17724 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n2 1.43709
R17725 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n0 0.281955
R17726 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n3 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t6 37.1981
R17727 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n5 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t5 31.4332
R17728 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n4 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t7 30.4613
R17729 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n4 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t4 24.7562
R17730 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n3 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t3 17.6611
R17731 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n5 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t2 15.3826
R17732 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n0 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 12.0716
R17733 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n5 7.62076
R17734 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n6 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 6.09789
R17735 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n7 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n2 2.99416
R17736 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n2 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t0 2.2755
R17737 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n2 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n1 2.2755
R17738 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n7 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n6 2.2505
R17739 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n0 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 2.24788
R17740 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n6 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n0 1.94903
R17741 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n4 1.81638
R17742 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n3 1.43706
R17743 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n7 0.4325
R17744 Vdiv105.n0 Vdiv105.t4 30.9379
R17745 Vdiv105.n0 Vdiv105.t5 21.6422
R17746 Vdiv105.n3 Vdiv105.t1 9.28805
R17747 Vdiv105 Vdiv105.n5 7.04952
R17748 Vdiv105.n2 Vdiv105.n1 6.01414
R17749 Vdiv105.n2 Vdiv105.t0 6.01414
R17750 Vdiv105 Vdiv105.n0 4.005
R17751 Vdiv105.n3 Vdiv105.n2 3.74829
R17752 Vdiv105.n5 Vdiv105.t2 3.74101
R17753 Vdiv105.n5 Vdiv105.n4 0.134848
R17754 Vdiv105.n4 Vdiv105.n3 0.0409348
R17755 Vdiv105.n4 Vdiv105 0.0031087
R17756 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n3 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t7 37.1981
R17757 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n5 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t5 31.4332
R17758 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n2 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t2 30.5752
R17759 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n2 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t3 24.6493
R17760 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n3 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t6 17.6611
R17761 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n4 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 17.0516
R17762 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n5 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t4 15.3826
R17763 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n5 7.62776
R17764 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n6 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n4 3.28711
R17765 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n7 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n1 2.99416
R17766 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n4 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 2.81128
R17767 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n6 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 2.67895
R17768 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t1 2.2755
R17769 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n0 2.2755
R17770 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n7 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n6 2.2505
R17771 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n2 1.80883
R17772 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n3 1.43706
R17773 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n7 0.4325
R17774 CLK_div_96_mag_0.JK_FF_mag_5.Q.n4 CLK_div_96_mag_0.JK_FF_mag_5.Q.t10 36.935
R17775 CLK_div_96_mag_0.JK_FF_mag_5.Q.n3 CLK_div_96_mag_0.JK_FF_mag_5.Q.t11 36.935
R17776 CLK_div_96_mag_0.JK_FF_mag_5.Q.n6 CLK_div_96_mag_0.JK_FF_mag_5.Q.t9 36.935
R17777 CLK_div_96_mag_0.JK_FF_mag_5.Q.n7 CLK_div_96_mag_0.JK_FF_mag_5.Q.t6 31.4332
R17778 CLK_div_96_mag_0.JK_FF_mag_5.Q.n5 CLK_div_96_mag_0.JK_FF_mag_5.Q.t4 25.5361
R17779 CLK_div_96_mag_0.JK_FF_mag_5.Q.n4 CLK_div_96_mag_0.JK_FF_mag_5.Q.t12 18.1962
R17780 CLK_div_96_mag_0.JK_FF_mag_5.Q.n3 CLK_div_96_mag_0.JK_FF_mag_5.Q.t3 18.1962
R17781 CLK_div_96_mag_0.JK_FF_mag_5.Q.n6 CLK_div_96_mag_0.JK_FF_mag_5.Q.t8 18.1962
R17782 CLK_div_96_mag_0.JK_FF_mag_5.Q.n7 CLK_div_96_mag_0.JK_FF_mag_5.Q.t5 15.3826
R17783 CLK_div_96_mag_0.JK_FF_mag_5.Q.n5 CLK_div_96_mag_0.JK_FF_mag_5.Q.t7 14.0734
R17784 CLK_div_96_mag_0.JK_FF_mag_5.Q CLK_div_96_mag_0.JK_FF_mag_5.Q.t0 7.09905
R17785 CLK_div_96_mag_0.JK_FF_mag_5.Q CLK_div_96_mag_0.JK_FF_mag_5.Q.n7 6.86029
R17786 CLK_div_96_mag_0.JK_FF_mag_5.Q.n8 CLK_div_96_mag_0.JK_FF_mag_5.Q 5.01077
R17787 CLK_div_96_mag_0.JK_FF_mag_5.Q.n9 CLK_div_96_mag_0.JK_FF_mag_5.Q 4.16836
R17788 CLK_div_96_mag_0.JK_FF_mag_5.Q CLK_div_96_mag_0.JK_FF_mag_5.Q.n2 3.25053
R17789 CLK_div_96_mag_0.JK_FF_mag_5.Q.n2 CLK_div_96_mag_0.JK_FF_mag_5.Q.t2 2.2755
R17790 CLK_div_96_mag_0.JK_FF_mag_5.Q.n2 CLK_div_96_mag_0.JK_FF_mag_5.Q.n1 2.2755
R17791 CLK_div_96_mag_0.JK_FF_mag_5.Q CLK_div_96_mag_0.JK_FF_mag_5.Q.n4 2.13151
R17792 CLK_div_96_mag_0.JK_FF_mag_5.Q.n0 CLK_div_96_mag_0.JK_FF_mag_5.Q 2.63808
R17793 CLK_div_96_mag_0.JK_FF_mag_5.Q CLK_div_96_mag_0.JK_FF_mag_5.Q.n9 2.34284
R17794 CLK_div_96_mag_0.JK_FF_mag_5.Q CLK_div_96_mag_0.JK_FF_mag_5.Q.n6 2.13459
R17795 CLK_div_96_mag_0.JK_FF_mag_5.Q CLK_div_96_mag_0.JK_FF_mag_5.Q.n3 2.13042
R17796 CLK_div_96_mag_0.JK_FF_mag_5.Q CLK_div_96_mag_0.JK_FF_mag_5.Q.n0 2.10738
R17797 CLK_div_96_mag_0.JK_FF_mag_5.Q.n9 CLK_div_96_mag_0.JK_FF_mag_5.Q.n8 1.52539
R17798 CLK_div_96_mag_0.JK_FF_mag_5.Q CLK_div_96_mag_0.JK_FF_mag_5.Q.n5 1.43628
R17799 CLK_div_96_mag_0.JK_FF_mag_5.Q.n8 CLK_div_96_mag_0.JK_FF_mag_5.Q 1.12067
R17800 CLK_div_96_mag_0.JK_FF_mag_5.Q CLK_div_96_mag_0.JK_FF_mag_5.Q.n0 1.11863
R17801 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t5 30.9379
R17802 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t4 30.664
R17803 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t2 24.5385
R17804 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t3 24.5101
R17805 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n2 7.46763
R17806 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n3 5.28703
R17807 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n1 4.09208
R17808 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 3.12156
R17809 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 1.86016
R17810 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n0 1.4252
R17811 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t4 37.1986
R17812 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t5 31.528
R17813 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t3 30.6344
R17814 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t6 27.3855
R17815 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t7 17.6614
R17816 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t8 15.3826
R17817 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n1 7.62751
R17818 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 6.09789
R17819 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n0 2.8877
R17820 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 2.67866
R17821 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n3 2.2505
R17822 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n2 1.43709
R17823 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.4325
R17824 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n5 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.t7 36.935
R17825 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n2 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.t10 31.4332
R17826 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n6 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.t4 31.4332
R17827 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n3 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.t8 30.4613
R17828 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n3 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.t5 24.7562
R17829 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n5 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.t3 18.1962
R17830 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n2 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.t9 15.3826
R17831 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n6 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.t6 15.3826
R17832 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n4 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1 8.5575
R17833 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.t2 7.09905
R17834 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n6 6.86029
R17835 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n2 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1 5.69501
R17836 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n7 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1 5.01077
R17837 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n1 3.25053
R17838 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n8 2.43532
R17839 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n1 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.t0 2.2755
R17840 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n1 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n0 2.2755
R17841 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n5 2.13459
R17842 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n3 1.81638
R17843 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n8 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n7 1.45395
R17844 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n8 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n4 1.23718
R17845 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n7 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1 1.12067
R17846 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n4 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1 0.976433
R17847 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n5 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.t3 36.935
R17848 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n2 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.t9 31.4332
R17849 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n6 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.t6 31.4332
R17850 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n3 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.t7 30.4613
R17851 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n3 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.t5 24.7562
R17852 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n5 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.t10 18.1962
R17853 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n2 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.t8 15.3826
R17854 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n6 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.t4 15.3826
R17855 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n4 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1 8.5575
R17856 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.t1 7.09905
R17857 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n6 6.86029
R17858 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n2 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1 5.69501
R17859 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n7 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1 5.01077
R17860 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n1 3.25053
R17861 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n8 2.43532
R17862 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n1 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.t0 2.2755
R17863 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n1 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n0 2.2755
R17864 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n5 2.13459
R17865 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n3 1.81638
R17866 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n8 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n7 1.45395
R17867 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n8 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n4 1.23718
R17868 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n7 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1 1.12067
R17869 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n4 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1 0.976433
R17870 Vdiv110 Vdiv110.n7 31.6239
R17871 Vdiv110.n3 Vdiv110.t4 30.9379
R17872 Vdiv110.n3 Vdiv110.t5 21.6422
R17873 Vdiv110.n11 Vdiv110.n10 9.28805
R17874 Vdiv110.n9 Vdiv110.n8 6.01414
R17875 Vdiv110.n9 Vdiv110.t0 6.01414
R17876 Vdiv110.n1 Vdiv110.n0 4.51956
R17877 Vdiv110.n4 Vdiv110.n2 4.51503
R17878 Vdiv110.n13 Vdiv110.n12 3.87405
R17879 Vdiv110.n11 Vdiv110.n9 3.74829
R17880 Vdiv110 Vdiv110.n3 2.8805
R17881 Vdiv110 Vdiv110.n1 2.251
R17882 Vdiv110.n2 Vdiv110.n0 2.24568
R17883 Vdiv110.n7 Vdiv110.n6 2.24307
R17884 Vdiv110.n5 Vdiv110 1.5005
R17885 Vdiv110.n13 Vdiv110.n11 0.0422391
R17886 Vdiv110 Vdiv110.n4 0.028625
R17887 Vdiv110.n7 Vdiv110.n0 0.0201512
R17888 Vdiv110.n6 Vdiv110.n1 0.0172252
R17889 Vdiv110.n5 Vdiv110.n2 0.0150082
R17890 Vdiv110.n4 Vdiv110 0.01175
R17891 Vdiv110 Vdiv110.n13 0.003
R17892 Vdiv110.n6 Vdiv110.n5 0.00275
R17893 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n4 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t4 37.1986
R17894 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n3 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t7 31.528
R17895 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n2 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t8 30.5184
R17896 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n2 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t6 24.7029
R17897 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n4 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t5 17.6614
R17898 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n3 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t3 15.3826
R17899 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n0 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 12.0843
R17900 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n0 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n3 9.86691
R17901 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n5 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 6.09789
R17902 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n7 2.99416
R17903 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n7 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t0 2.2755
R17904 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n7 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n6 2.2755
R17905 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n5 2.2505
R17906 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n0 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 2.24173
R17907 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n5 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n0 1.93723
R17908 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n2 1.81225
R17909 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n4 1.43709
R17910 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n1 0.281955
R17911 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n3 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t5 37.1981
R17912 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n5 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t4 31.4332
R17913 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n4 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t3 30.4613
R17914 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n4 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t7 24.7562
R17915 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n3 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t2 17.6611
R17916 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n5 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t6 15.3826
R17917 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n0 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 12.0716
R17918 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n5 7.62076
R17919 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n6 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 6.09789
R17920 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n7 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n2 2.99416
R17921 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n2 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t1 2.2755
R17922 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n2 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n1 2.2755
R17923 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n7 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n6 2.2505
R17924 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n0 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 2.24788
R17925 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n6 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n0 1.94903
R17926 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n4 1.81638
R17927 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n3 1.43706
R17928 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n7 0.4325
R17929 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n8 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t6 36.935
R17930 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n7 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t4 36.935
R17931 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n12 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t2 36.935
R17932 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n9 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t9 36.935
R17933 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n10 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t5 30.5752
R17934 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n13 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t3 25.4744
R17935 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n6 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t7 25.4742
R17936 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n10 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t8 21.7814
R17937 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n8 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t12 18.1962
R17938 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n7 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t11 18.1962
R17939 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n12 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t10 18.1962
R17940 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n9 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t14 18.1962
R17941 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n6 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t15 14.142
R17942 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n13 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t13 14.1417
R17943 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n5 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t0 9.33985
R17944 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n0 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n11 7.41483
R17945 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n15 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n14 5.37091
R17946 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n5 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t1 5.17836
R17947 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n2 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n12 2.13265
R17948 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n2 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK 0.077103
R17949 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n13 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n3 1.42996
R17950 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n0 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n2 1.11863
R17951 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n14 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n3 1.19586
R17952 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n8 2.13265
R17953 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n11 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n10 1.80883
R17954 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n1 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK 2.63776
R17955 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n0 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK 2.51943
R17956 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n9 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK 2.13281
R17957 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n7 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK 2.13261
R17958 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n4 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n6 1.43004
R17959 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n3 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK 0.196041
R17960 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n4 0.196041
R17961 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n5 0.115328
R17962 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n11 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK 0.108371
R17963 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n4 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n15 1.19586
R17964 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n1 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK 1.11863
R17965 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n14 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n0 1.01264
R17966 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n15 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n1 0.894314
R17967 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t6 37.1986
R17968 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t8 31.528
R17969 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t5 30.6344
R17970 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t7 27.3855
R17971 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t3 17.6614
R17972 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t4 15.3826
R17973 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n1 7.62751
R17974 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 6.09789
R17975 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n5 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t1 2.99416
R17976 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n0 2.8877
R17977 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 2.67866
R17978 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n4 2.2755
R17979 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n5 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n3 2.2505
R17980 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n2 1.43709
R17981 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n5 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.4325
R17982 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n5 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.t3 36.935
R17983 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n4 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.t6 31.4332
R17984 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n6 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.t4 31.4332
R17985 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n3 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.t9 30.5184
R17986 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n3 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.t7 24.7029
R17987 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n5 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.t5 18.1962
R17988 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n4 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.t10 15.3826
R17989 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n6 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.t8 15.3826
R17990 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.t1 7.09905
R17991 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n6 6.86134
R17992 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n7 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1 5.0096
R17993 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n0 8.55639
R17994 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n4 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1 5.69501
R17995 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n2 3.25226
R17996 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n8 2.43532
R17997 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n2 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.t2 2.2755
R17998 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n2 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n1 2.2755
R17999 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n5 2.13479
R18000 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n3 1.81225
R18001 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n8 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n7 1.45511
R18002 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n8 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n0 1.23718
R18003 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n7 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1 1.12056
R18004 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n0 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1 0.976034
R18005 Vdiv108.n9 Vdiv108.t4 36.935
R18006 Vdiv108.n0 Vdiv108.t8 31.528
R18007 Vdiv108.n7 Vdiv108.t7 31.528
R18008 Vdiv108.n9 Vdiv108.t6 18.1962
R18009 Vdiv108.n0 Vdiv108.t5 15.3826
R18010 Vdiv108.n7 Vdiv108.t3 15.3826
R18011 Vdiv108.n1 Vdiv108.n0 8.74076
R18012 Vdiv108.n5 Vdiv108.n2 7.09905
R18013 Vdiv108.n8 Vdiv108.n7 6.86134
R18014 Vdiv108.n11 Vdiv108.n10 5.01109
R18015 Vdiv108.n5 Vdiv108.n4 3.25085
R18016 Vdiv108.n12 Vdiv108.n6 2.36461
R18017 Vdiv108.n4 Vdiv108.t0 2.2755
R18018 Vdiv108.n4 Vdiv108.n3 2.2755
R18019 Vdiv108.n10 Vdiv108.n9 2.13398
R18020 Vdiv108.n12 Vdiv108.n11 1.47724
R18021 Vdiv108.n11 Vdiv108.n8 1.12725
R18022 Vdiv108 Vdiv108.n12 0.914492
R18023 Vdiv108 Vdiv108.n1 0.116616
R18024 Vdiv108.n6 Vdiv108.n5 0.0919062
R18025 Vdiv108.n8 Vdiv108 0.0857632
R18026 Vdiv108.n10 Vdiv108 0.0810725
R18027 Vdiv108.n6 Vdiv108 0.073625
R18028 Vdiv108.n1 Vdiv108 0.00202542
R18029 CLK_div_96_mag_0.JK_FF_mag_4.Q.n7 CLK_div_96_mag_0.JK_FF_mag_4.Q.t3 36.935
R18030 CLK_div_96_mag_0.JK_FF_mag_4.Q.n6 CLK_div_96_mag_0.JK_FF_mag_4.Q.t12 36.935
R18031 CLK_div_96_mag_0.JK_FF_mag_4.Q.n3 CLK_div_96_mag_0.JK_FF_mag_4.Q.t8 36.935
R18032 CLK_div_96_mag_0.JK_FF_mag_4.Q.n4 CLK_div_96_mag_0.JK_FF_mag_4.Q.t6 31.4332
R18033 CLK_div_96_mag_0.JK_FF_mag_4.Q.n8 CLK_div_96_mag_0.JK_FF_mag_4.Q.t10 25.4744
R18034 CLK_div_96_mag_0.JK_FF_mag_4.Q.n7 CLK_div_96_mag_0.JK_FF_mag_4.Q.t4 18.1962
R18035 CLK_div_96_mag_0.JK_FF_mag_4.Q.n6 CLK_div_96_mag_0.JK_FF_mag_4.Q.t11 18.1962
R18036 CLK_div_96_mag_0.JK_FF_mag_4.Q.n3 CLK_div_96_mag_0.JK_FF_mag_4.Q.t7 18.1962
R18037 CLK_div_96_mag_0.JK_FF_mag_4.Q.n4 CLK_div_96_mag_0.JK_FF_mag_4.Q.t5 15.3826
R18038 CLK_div_96_mag_0.JK_FF_mag_4.Q.n8 CLK_div_96_mag_0.JK_FF_mag_4.Q.t9 14.1417
R18039 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.JK_FF_mag_4.Q.t1 7.09905
R18040 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.JK_FF_mag_4.Q.n4 6.86029
R18041 CLK_div_96_mag_0.JK_FF_mag_4.Q.n9 CLK_div_96_mag_0.JK_FF_mag_4.Q 6.35399
R18042 CLK_div_96_mag_0.JK_FF_mag_4.Q.n5 CLK_div_96_mag_0.JK_FF_mag_4.Q 5.01077
R18043 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.JK_FF_mag_4.Q.n2 3.25053
R18044 CLK_div_96_mag_0.JK_FF_mag_4.Q.n2 CLK_div_96_mag_0.JK_FF_mag_4.Q.t0 2.2755
R18045 CLK_div_96_mag_0.JK_FF_mag_4.Q.n2 CLK_div_96_mag_0.JK_FF_mag_4.Q.n1 2.2755
R18046 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.JK_FF_mag_4.Q.n7 2.13265
R18047 CLK_div_96_mag_0.JK_FF_mag_4.Q.n0 CLK_div_96_mag_0.JK_FF_mag_4.Q 2.63776
R18048 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.JK_FF_mag_4.Q.n9 2.3405
R18049 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.JK_FF_mag_4.Q.n3 2.13459
R18050 CLK_div_96_mag_0.JK_FF_mag_4.Q.n6 CLK_div_96_mag_0.JK_FF_mag_4.Q 2.13261
R18051 CLK_div_96_mag_0.JK_FF_mag_4.Q.n9 CLK_div_96_mag_0.JK_FF_mag_4.Q.n5 1.54877
R18052 CLK_div_96_mag_0.JK_FF_mag_4.Q.n0 CLK_div_96_mag_0.JK_FF_mag_4.Q 2.1039
R18053 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.JK_FF_mag_4.Q.n8 1.62425
R18054 CLK_div_96_mag_0.JK_FF_mag_4.Q.n5 CLK_div_96_mag_0.JK_FF_mag_4.Q 1.12067
R18055 CLK_div_96_mag_0.JK_FF_mag_4.Q.n0 CLK_div_96_mag_0.JK_FF_mag_4.Q 1.11863
R18056 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n17 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t13 36.935
R18057 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n18 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t11 36.935
R18058 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n12 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t5 36.935
R18059 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n19 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t3 31.4332
R18060 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n14 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t7 31.4332
R18061 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n20 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t12 30.9379
R18062 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n22 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t10 25.4744
R18063 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n20 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t15 21.6422
R18064 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n17 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t8 18.1962
R18065 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n18 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t9 18.1962
R18066 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n12 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t4 18.1962
R18067 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n19 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t16 15.3826
R18068 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n14 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t6 15.3826
R18069 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n22 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t14 14.1417
R18070 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n11 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t1 7.09905
R18071 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n15 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n14 6.86029
R18072 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n16 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n13 5.01077
R18073 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n2 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n4 0.0219501
R18074 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n1 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n0 0.0360559
R18075 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n19 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 5.69501
R18076 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n4 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n1 2.23369
R18077 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n2 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n0 1.11499
R18078 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n23 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n8 2.2429
R18079 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n8 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n7 0.0171915
R18080 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n11 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n10 3.25053
R18081 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n10 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t2 2.2755
R18082 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n10 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n9 2.2755
R18083 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n25 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n24 2.2505
R18084 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n7 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n6 2.24196
R18085 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n13 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n12 2.13459
R18086 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n3 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n20 2.13074
R18087 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n4 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n17 2.12093
R18088 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n1 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n5 2.64237
R18089 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n0 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n21 4.95192
R18090 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n21 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 4.19069
R18091 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n24 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n16 1.52773
R18092 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n18 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n5 2.13281
R18093 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n7 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n22 1.42118
R18094 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n16 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n15 1.12067
R18095 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n6 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n0 0.960138
R18096 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n23 0.646487
R18097 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n8 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 0.187192
R18098 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n25 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n11 0.0905
R18099 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n15 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 0.0857632
R18100 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n25 0.0834687
R18101 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n13 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 0.0800273
R18102 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n3 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 0.0980715
R18103 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n2 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 0.0672526
R18104 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n5 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 0.0771461
R18105 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n24 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 0.0322045
R18106 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n23 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n6 0.0238218
R18107 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n21 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n3 2.08419
R18108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.n3 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.t4 36.935
R18109 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.n4 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.t6 31.4332
R18110 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.n2 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.t5 29.8635
R18111 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.n2 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.t7 27.7543
R18112 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.n3 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.t8 18.1962
R18113 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.n4 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.t3 15.3826
R18114 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.t2 7.09905
R18115 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.n4 6.86134
R18116 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.n5 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 5.0096
R18117 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.n6 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 3.41823
R18118 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.n1 3.25226
R18119 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.n1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.t0 2.2755
R18120 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.n1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.n0 2.2755
R18121 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.n6 2.2505
R18122 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.n3 2.13479
R18123 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.n2 1.7371
R18124 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.n6 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.n5 1.50498
R18125 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.n5 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 1.12056
R18126 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.n5 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.t5 37.1984
R18127 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.n4 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.t7 31.4332
R18128 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.n3 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.t3 30.5184
R18129 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.n3 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.t2 24.7029
R18130 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.n5 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.t6 17.6618
R18131 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.n4 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.t4 15.3826
R18132 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.n0 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K 12.0839
R18133 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.n0 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.n4 9.86691
R18134 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.n6 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K 6.09789
R18135 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.n7 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.n2 2.99416
R18136 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.n2 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.t0 2.2755
R18137 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.n2 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.n1 2.2755
R18138 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.n7 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.n6 2.2505
R18139 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.n0 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K 2.24134
R18140 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.n6 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.n0 1.93723
R18141 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.n3 1.81224
R18142 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.n5 1.43718
R18143 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.n7 0.4325
R18144 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n7 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t2 36.935
R18145 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n6 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t9 36.935
R18146 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n11 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t11 36.935
R18147 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n10 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t8 36.935
R18148 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n8 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t6 30.6315
R18149 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n15 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t4 25.5361
R18150 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n12 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t14 25.5361
R18151 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n8 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t10 21.7275
R18152 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n7 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t5 18.1962
R18153 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n6 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t13 18.1962
R18154 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n11 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t15 18.1962
R18155 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n10 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t3 18.1962
R18156 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n15 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t12 14.0734
R18157 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n12 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t7 14.0734
R18158 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n5 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t1 9.33985
R18159 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n0 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n9 7.41366
R18160 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n14 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n13 5.37352
R18161 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n5 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t0 5.17836
R18162 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n7 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK 2.13258
R18163 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n0 1.11745
R18164 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n11 2.13258
R18165 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n9 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n8 1.80525
R18166 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK 2.63808
R18167 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n0 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK 2.51975
R18168 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n10 2.13055
R18169 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n6 2.13055
R18170 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n3 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n12 1.43653
R18171 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n4 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n15 1.43653
R18172 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n3 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK 0.196042
R18173 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n4 0.196042
R18174 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n5 0.115328
R18175 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n9 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK 0.108371
R18176 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK 0.0763652
R18177 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n13 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n3 1.19546
R18178 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n4 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n14 1.19546
R18179 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n1 1.11745
R18180 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n13 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n0 1.01362
R18181 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n14 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n1 0.895294
R18182 Vdiv99.n2 Vdiv99.t3 30.9379
R18183 Vdiv99.n2 Vdiv99.t2 21.6422
R18184 Vdiv99 Vdiv99.n7 15.3654
R18185 Vdiv99.n10 Vdiv99.n9 9.33985
R18186 Vdiv99.n10 Vdiv99.n8 5.17836
R18187 Vdiv99.n5 Vdiv99.n0 4.5097
R18188 Vdiv99.n5 Vdiv99.n4 4.5005
R18189 Vdiv99 Vdiv99.n2 2.8805
R18190 Vdiv99 Vdiv99.n3 2.26066
R18191 Vdiv99.n3 Vdiv99.n0 2.25077
R18192 Vdiv99 Vdiv99.n1 1.5005
R18193 Vdiv99.n7 Vdiv99.n6 1.49782
R18194 Vdiv99 Vdiv99.n10 0.115328
R18195 Vdiv99.n4 Vdiv99 0.0281136
R18196 Vdiv99.n6 Vdiv99.n5 0.0270909
R18197 Vdiv99.n7 Vdiv99.n0 0.0118561
R18198 Vdiv99.n3 Vdiv99.n1 0.0101206
R18199 Vdiv99.n4 Vdiv99 0.00868182
R18200 Vdiv99.n6 Vdiv99.n1 0.00152273
R18201 Vdiv93.n0 Vdiv93.t2 30.9379
R18202 Vdiv93.n0 Vdiv93.t3 21.6422
R18203 Vdiv93.n3 Vdiv93.n2 9.33985
R18204 Vdiv93.n3 Vdiv93.n1 5.17836
R18205 Vdiv93 Vdiv93.n0 4.00478
R18206 Vdiv93 Vdiv93.n3 0.0749828
R18207 F1.n20 F1.t7 36.935
R18208 F1.n14 F1.t10 36.935
R18209 F1.n8 F1.t11 36.859
R18210 F1.n29 F1.t5 36.8284
R18211 F1.n44 F1.t8 31.528
R18212 F1.n50 F1.t4 31.528
R18213 F1.n58 F1.t0 25.7638
R18214 F1.n48 F1.t1 25.7638
R18215 F1.n2 F1.t16 25.515
R18216 F1.n20 F1.t3 18.1962
R18217 F1.n14 F1.t6 18.1962
R18218 F1.n7 F1.t9 17.5837
R18219 F1.n28 F1.t2 17.2177
R18220 F1.n44 F1.t13 15.3826
R18221 F1.n50 F1.t14 15.3826
R18222 F1.n58 F1.t15 13.2969
R18223 F1.n48 F1.t12 13.2969
R18224 F1.n1 F1.t17 12.3792
R18225 F1.n62 F1.n61 9.60207
R18226 F1 F1.n8 8.03007
R18227 F1 F1.n29 8.02697
R18228 F1.n14 F1 8.02621
R18229 F1.n45 F1.n44 7.62076
R18230 F1.n51 F1.n50 7.62076
R18231 F1.n57 F1.n56 6.90126
R18232 F1.n39 F1.n19 5.77472
R18233 F1.n46 F1.n43 4.54699
R18234 F1.n53 F1.n52 4.54699
R18235 F1.n60 F1 4.52833
R18236 F1.n54 F1 4.52833
R18237 F1.n35 F1.n34 4.5005
R18238 F1.n32 F1.n27 4.5005
R18239 F1.n32 F1.n31 4.5005
R18240 F1.n35 F1.n26 4.5005
R18241 F1.n3 F1.n2 4.5005
R18242 F1.n42 F1.n41 4.5005
R18243 F1 F1.n62 3.66527
R18244 F1.n30 F1.n28 3.61051
R18245 F1.n23 F1.n22 2.99669
R18246 F1.n40 F1.n39 2.96288
R18247 F1.n15 F1.n14 2.88073
R18248 F1.n39 F1.n38 2.64379
R18249 F1.n62 F1.n42 2.53643
R18250 F1 F1.n0 2.2713
R18251 F1.n59 F1.n57 2.25478
R18252 F1.n19 F1.n18 2.25429
R18253 F1.n56 F1.n49 2.25386
R18254 F1.n36 F1.n35 2.2505
R18255 F1.n55 F1.n49 2.2505
R18256 F1.n59 F1.n47 2.2505
R18257 F1.n11 F1.n10 2.24478
R18258 F1.n40 F1.n4 2.24169
R18259 F1.n1 F1 2.20908
R18260 F1.n21 F1.n20 2.1208
R18261 F1.n59 F1.n58 2.11815
R18262 F1.n49 F1.n48 2.11815
R18263 F1.n9 F1.n7 1.81009
R18264 F1.n12 F1.n11 1.63145
R18265 F1.n54 F1.n53 1.33991
R18266 F1.n61 F1.n60 1.28387
R18267 F1.n18 F1.n17 1.12663
R18268 F1.n46 F1.n45 1.12145
R18269 F1.n53 F1.n51 1.12145
R18270 F1.n29 F1.n28 0.857233
R18271 F1.n2 F1.n1 0.775233
R18272 F1.n8 F1.n7 0.435263
R18273 F1.n43 F1 0.0780197
R18274 F1.n52 F1 0.0780197
R18275 F1.n6 F1 0.0768393
R18276 F1.n22 F1 0.0752567
R18277 F1.n34 F1 0.0719706
R18278 F1.n61 F1.n46 0.0551093
R18279 F1.n17 F1 0.0464863
R18280 F1.n52 F1 0.0359098
R18281 F1 F1.n43 0.032959
R18282 F1.n38 F1.n37 0.0320584
R18283 F1.n10 F1.n6 0.0300714
R18284 F1.n55 F1.n54 0.0289694
R18285 F1.n60 F1.n47 0.0289694
R18286 F1.n35 F1.n24 0.0273831
R18287 F1.n42 F1.n4 0.0249444
R18288 F1 F1.n40 0.0237688
R18289 F1.n17 F1.n16 0.0215918
R18290 F1.n11 F1.n5 0.0177728
R18291 F1.n57 F1 0.0169815
R18292 F1.n56 F1 0.0160631
R18293 F1.n22 F1.n21 0.0144304
R18294 F1.n10 F1.n9 0.00692857
R18295 F1.n24 F1.n23 0.00517532
R18296 F1.n4 F1.n3 0.00494444
R18297 F1.n18 F1.n13 0.00484133
R18298 F1.n31 F1.n30 0.00447059
R18299 F1.n26 F1.n25 0.00314706
R18300 F1.n15 F1 0.00291681
R18301 F1.n33 F1.n32 0.00283766
R18302 F1 F1.n55 0.00233673
R18303 F1 F1.n47 0.00233673
R18304 F1.n21 F1 0.00212278
R18305 F1.n45 F1 0.00197541
R18306 F1 F1.n51 0.00197541
R18307 F1.n41 F1 0.00188462
R18308 F1.n30 F1 0.00182353
R18309 F1.n9 F1 0.00178571
R18310 F1.n35 F1.n33 0.00166883
R18311 F1.n37 F1.n36 0.00166883
R18312 F1.n3 F1 0.00161111
R18313 F1.n13 F1.n12 0.00159756
R18314 F1 F1.n59 0.00142783
R18315 F1 F1.n49 0.00142783
R18316 F1.n16 F1.n15 0.00142074
R18317 F2.n10 F2.t11 36.7069
R18318 F2.n24 F2.t12 36.5548
R18319 F2.n35 F2.t0 31.528
R18320 F2.n16 F2.t5 30.9379
R18321 F2.n2 F2.t6 30.4206
R18322 F2.n39 F2.t13 25.7638
R18323 F2.n2 F2.t8 24.7698
R18324 F2.n16 F2.t7 24.5101
R18325 F2.n30 F2.t1 23.4411
R18326 F2.n23 F2.t10 17.4145
R18327 F2.n9 F2.t9 17.3258
R18328 F2.n35 F2.t2 15.3826
R18329 F2.n43 F2.n42 13.8981
R18330 F2.n39 F2.t4 13.2969
R18331 F2.n31 F2.t3 10.8912
R18332 F2.n19 F2.n13 10.468
R18333 F2 F2.n29 8.62191
R18334 F2.n31 F2 8.0298
R18335 F2.n10 F2 8.02962
R18336 F2.n24 F2 8.02588
R18337 F2.n36 F2.n35 7.6289
R18338 F2.n41 F2 4.52833
R18339 F2.n7 F2.n6 4.5005
R18340 F2.n11 F2.n6 4.5005
R18341 F2.n11 F2.n10 4.5005
R18342 F2 F2.n1 4.5005
R18343 F2.n3 F2.n1 4.5005
R18344 F2.n28 F2.n27 4.5005
R18345 F2.n28 F2.n25 4.5005
R18346 F2.n25 F2.n24 4.5005
R18347 F2.n23 F2.n22 3.66972
R18348 F2.n9 F2.n8 3.63801
R18349 F2 F2.n43 3.02778
R18350 F2 F2.n16 2.8805
R18351 F2.n43 F2.n34 2.81046
R18352 F2.n32 F2.n31 2.40618
R18353 F2.n32 F2.n30 2.32323
R18354 F2 F2.n0 2.27492
R18355 F2.n38 F2 2.26613
R18356 F2.n17 F2 2.25751
R18357 F2.n18 F2.n14 2.251
R18358 F2.n40 F2.n37 2.2505
R18359 F2.n13 F2.n12 2.24496
R18360 F2.n5 F2.n4 2.2444
R18361 F2.n17 F2.n15 2.24399
R18362 F2.n33 F2.n32 2.11815
R18363 F2.n40 F2.n39 2.11815
R18364 F2.n21 F2.n20 1.66028
R18365 F2.n33 F2 1.50158
R18366 F2.n26 F2.n21 1.49405
R18367 F2 F2.n2 1.42163
R18368 F2.n42 F2.n41 1.28387
R18369 F2.n24 F2.n23 1.04377
R18370 F2.n10 F2.n9 0.955106
R18371 F2.n42 F2.n36 0.948428
R18372 F2.n20 F2.n19 0.575955
R18373 F2.n27 F2 0.484751
R18374 F2.n20 F2.n5 0.381035
R18375 F2.n19 F2.n18 0.296719
R18376 F2.n3 F2 0.192359
R18377 F2.n36 F2 0.108522
R18378 F2.n15 F2 0.0938405
R18379 F2.n7 F2 0.041692
R18380 F2.n12 F2.n7 0.0309412
R18381 F2.n41 F2.n37 0.0289694
R18382 F2.n4 F2.n3 0.0275
R18383 F2.n27 F2.n26 0.0270385
R18384 F2.n29 F2.n21 0.0255368
R18385 F2.n13 F2.n6 0.0200059
R18386 F2.n5 F2.n1 0.017373
R18387 F2.n18 F2.n17 0.0152683
R18388 F2.n15 F2.n14 0.0150187
R18389 F2.n4 F2 0.00725
R18390 F2.n26 F2.n25 0.00626923
R18391 F2.n40 F2.n38 0.00563331
R18392 F2.n12 F2.n11 0.00447059
R18393 F2.n29 F2.n28 0.00284618
R18394 F2 F2.n37 0.00233673
R18395 F2.n38 F2 0.00193332
R18396 F2.n11 F2.n8 0.00182353
R18397 F2 F2.n8 0.00182353
R18398 F2.n25 F2.n22 0.00165385
R18399 F2 F2.n22 0.00165385
R18400 F2 F2.n14 0.001625
R18401 F2.n34 F2.n33 0.00154651
R18402 F2.n33 F2 0.00154651
R18403 F2 F2.n40 0.00142783
R18404 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n2 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t5 37.1981
R18405 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n4 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t3 31.528
R18406 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n3 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t8 30.4613
R18407 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n3 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t7 24.7562
R18408 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n2 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t6 17.6611
R18409 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n4 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t4 15.3826
R18410 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n0 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 12.0856
R18411 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n0 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n4 9.86714
R18412 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n5 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 6.09789
R18413 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n7 2.99416
R18414 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n7 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t0 2.2755
R18415 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n7 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n6 2.2755
R18416 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n5 2.2505
R18417 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n0 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 2.24173
R18418 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n5 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n0 1.93771
R18419 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n3 1.81589
R18420 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n2 1.43706
R18421 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n1 0.281955
R18422 Vdiv90.n0 Vdiv90.t5 31.528
R18423 Vdiv90.n0 Vdiv90.t4 15.3826
R18424 Vdiv90 Vdiv90.n11 13.6025
R18425 Vdiv90.n9 Vdiv90.n8 9.28675
R18426 Vdiv90 Vdiv90.n0 7.62076
R18427 Vdiv90.n7 Vdiv90.n6 6.01414
R18428 Vdiv90.n7 Vdiv90.t3 6.01414
R18429 Vdiv90.n12 Vdiv90 4.73174
R18430 Vdiv90.n15 Vdiv90 4.53864
R18431 Vdiv90 Vdiv90.n16 4.5005
R18432 Vdiv90.n10 Vdiv90.n5 3.88449
R18433 Vdiv90.n9 Vdiv90.n7 3.74699
R18434 Vdiv90.n4 Vdiv90.n3 1.5005
R18435 Vdiv90.n14 Vdiv90.n13 1.5005
R18436 Vdiv90.n11 Vdiv90 0.0927551
R18437 Vdiv90.n11 Vdiv90 0.0814453
R18438 Vdiv90.n2 Vdiv90 0.0633894
R18439 Vdiv90.n3 Vdiv90.n2 0.040161
R18440 Vdiv90.n13 Vdiv90.n12 0.036125
R18441 Vdiv90.n10 Vdiv90.n9 0.0331087
R18442 Vdiv90.n16 Vdiv90.n15 0.0236683
R18443 Vdiv90.n3 Vdiv90 0.0127034
R18444 Vdiv90.n4 Vdiv90.n1 0.0124954
R18445 Vdiv90.n16 Vdiv90.n14 0.00673762
R18446 Vdiv90 Vdiv90.n10 0.00269512
R18447 Vdiv90.n14 Vdiv90.n4 0.00228218
R18448 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t4 30.9379
R18449 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t5 30.664
R18450 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t3 24.5385
R18451 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t2 24.5101
R18452 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n2 7.46763
R18453 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n3 5.28703
R18454 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n1 4.09208
R18455 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 3.12156
R18456 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 1.86016
R18457 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n0 1.4252
C0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.198f
C1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 1.33e-19
C2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.CLK 0.123f
C3 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 a_46777_1671# 0.00118f
C4 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_48712_n17599# 0.0036f
C5 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN 2.39e-20
C6 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 2.01e-19
C7 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT a_55019_7683# 0.0294f
C8 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT 0.16f
C9 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_53738_n1102# 1.43e-19
C10 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.27f
C11 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K Vdiv100 4.19e-19
C12 VDD96 a_28577_n2996# 0.00108f
C13 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.16f
C14 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.113f
C15 VDD105 a_45006_10154# 2.21e-19
C16 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.IN2 0.49f
C17 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_28093_n18723# 3.33e-19
C18 RST a_23019_5018# 8.64e-19
C19 Vdiv100 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 0.0265f
C20 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT a_25318_6115# 0.0203f
C21 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00118f
C22 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_54669_2768# 0.0202f
C23 CLK_div_96_mag_0.JK_FF_mag_4.Q a_23703_n287# 0.00939f
C24 VDD110 a_44625_n15583# 3.14e-19
C25 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 0.122f
C26 a_47030_n16726# a_47190_n16726# 0.0504f
C27 VDD105 a_45724_9057# 2.21e-19
C28 VDD110 a_47030_n16726# 2.21e-19
C29 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0156f
C30 RST CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.067f
C31 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 0.00335f
C32 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 0.215f
C33 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.159f
C34 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_30315_n15493# 0.00118f
C35 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 a_22711_n14504# 0.0177f
C36 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_96_mag_0.JK_FF_mag_0.Q 7.24e-19
C37 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 a_47187_2768# 0.0036f
C38 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT 5.76e-22
C39 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00243f
C40 RST a_35943_n10028# 0.00218f
C41 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_53973_n6862# 0.0733f
C42 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 3.81e-19
C43 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 a_46867_7960# 0.0084f
C44 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 5.11e-19
C45 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.0543f
C46 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_50304_n16724# 0.00789f
C47 F1 Vdiv100 0.074f
C48 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0129f
C49 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB a_21995_n7106# 2.96e-19
C50 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB a_52657_2768# 0.0811f
C51 CLK_div_96_mag_0.JK_FF_mag_5.Q a_23703_n287# 2.79e-20
C52 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 2.57e-20
C53 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 2.11e-20
C54 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 a_28010_n9876# 1.46e-19
C55 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 dec3x8_ibr_mag_0.and_3_ibr_1.nand3_mag_ibr_0.OUT 0.32f
C56 RST a_44436_9057# 0.0011f
C57 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.IN1 a_22575_n287# 0.0059f
C58 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.11f
C59 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.00975f
C60 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 2.81e-20
C61 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.231f
C62 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_53008_n2243# 0.0202f
C63 a_43751_n5176# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1.5e-20
C64 a_44315_n5176# a_44475_n5176# 0.0504f
C65 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_30244_398# 0.00372f
C66 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_23289_n6009# 0.0202f
C67 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.0635f
C68 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.215f
C69 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.884f
C70 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_33744_n17626# 0.00378f
C71 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.107f
C72 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.361f
C73 dec3x8_ibr_mag_0.and_3_ibr_3.nand3_mag_ibr_0.OUT a_39580_6821# 0.0779f
C74 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 0.00238f
C75 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0187f
C76 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.25f
C77 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.122f
C78 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_96_mag_0.JK_FF_mag_2.Q 0.107f
C79 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_30881_n18723# 2.96e-19
C80 CLK CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 1.22e-19
C81 CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 a_54978_6284# 0.069f
C82 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_42521_n13474# 0.00186f
C83 RST CLK_div_90_mag_0.CLK_div_10_mag_0.CLK 5.44e-19
C84 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 0.0286f
C85 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 a_45815_n1102# 8.17e-21
C86 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 0.0138f
C87 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.768f
C88 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB 0.25f
C89 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_26036_5018# 0.00695f
C90 RST CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.11f
C91 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN 0.0116f
C92 VDD110 a_48558_n18696# 3.14e-19
C93 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 0.00488f
C94 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 CLK_div_96_mag_0.JK_FF_mag_0.Q 0.00107f
C95 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN 0.316f
C96 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 0.149f
C97 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_37391_n9984# 0.00378f
C98 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_50441_n17599# 0.00789f
C99 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_26099_398# 1.43e-19
C100 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_23743_5062# 0.0036f
C101 RST CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 4.25e-20
C102 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 2.77e-19
C103 Vdiv96 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT 0.282f
C104 RST a_53221_2768# 9.41e-19
C105 CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 4.52e-20
C106 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.00118f
C107 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.765f
C108 RST a_26208_n2996# 0.00193f
C109 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_30727_n17626# 0.069f
C110 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_2x1_ibr_0.I0 0.234f
C111 VDD a_38294_6821# 2.21e-19
C112 a_28329_5018# a_28489_5018# 0.0504f
C113 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 1.82e-19
C114 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT a_48475_2768# 1.5e-20
C115 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT 0.306f
C116 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.0106f
C117 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_4.IN2 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_1.IN2 8.16e-20
C118 RST a_53309_n15631# 9.41e-19
C119 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.0725f
C120 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C121 VDD99 a_23948_n18723# 3.56e-19
C122 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 6.71e-19
C123 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_47086_5143# 2.81e-19
C124 RST a_53463_n16728# 0.00256f
C125 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.00183f
C126 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.11f
C127 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 7.08e-20
C128 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.0718f
C129 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00264f
C130 RST a_54456_n2199# 9.41e-19
C131 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 a_36024_n15495# 0.069f
C132 CLK_div_96_mag_0.JK_FF_mag_5.Q a_22988_n1789# 6.43e-21
C133 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 0.00586f
C134 CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0175f
C135 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_44282_10154# 0.069f
C136 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 9.98e-19
C137 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 7.24e-19
C138 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00166f
C139 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 4.42e-19
C140 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K a_45612_1671# 8.64e-19
C141 CLK_div_90_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.144f
C142 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_27180_n15491# 0.00118f
C143 F1 dec3x8_ibr_mag_0.and_3_ibr_3.nand3_mag_ibr_0.OUT 0.24f
C144 dec3x8_ibr_mag_0.and_3_ibr_0.nand3_mag_ibr_0.OUT a_37168_6821# 6.08e-20
C145 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 1.27f
C146 RST CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 0.00594f
C147 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.283f
C148 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.343f
C149 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 1.54e-21
C150 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.25f
C151 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 0.0146f
C152 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK a_39690_n8887# 6.43e-21
C153 VDD100 a_53785_2768# 0.00101f
C154 RST a_44324_1671# 0.0011f
C155 VDD90 a_22461_6115# 2.66e-19
C156 CLK a_22405_n6009# 0.00133f
C157 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.159f
C158 CLK a_49098_5187# 5.03e-19
C159 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 a_48098_n10160# 1.01e-20
C160 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT a_50922_1671# 0.0202f
C161 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 2f
C162 VDD110 a_41124_n16098# 3.14e-19
C163 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_29307_n1855# 0.0202f
C164 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.414f
C165 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 6.08e-19
C166 CLK CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 7.81e-19
C167 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C168 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.359f
C169 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN a_55197_n20487# 2.85e-20
C170 CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.11f
C171 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB a_24784_n8778# 1.4e-20
C172 VDD100 a_55020_n2199# 3.14e-19
C173 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I1 a_36873_n1822# 0.069f
C174 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 2.04e-19
C175 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.233f
C176 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 0.00975f
C177 a_51487_n10161# m3_20882_n11188# 0.00102f
C178 VDD108 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.653f
C179 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00161f
C180 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 a_29241_7256# 0.0105f
C181 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 3.88e-20
C182 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 a_25646_n17626# 6.04e-19
C183 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.654f
C184 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_26984_10099# 0.0732f
C185 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.0685f
C186 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.231f
C187 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 1.41e-20
C188 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 a_32750_n7675# 1.78e-19
C189 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 6.11e-20
C190 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0134f
C191 VDD108 a_50232_n7685# 0.165f
C192 VDD mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT 0.655f
C193 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.395f
C194 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0209f
C195 VDD100 a_44888_1671# 3.14e-19
C196 a_23948_n13382# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 2.69e-22
C197 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 0.0781f
C198 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 a_45458_2768# 0.00789f
C199 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK a_44253_n18696# 0.0101f
C200 RST CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.391f
C201 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.00183f
C202 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0129f
C203 CLK_div_96_mag_0.JK_FF_mag_5.Q CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.426f
C204 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN m3_20882_n11188# 0.00133f
C205 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00183f
C206 VDD110 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 8.33e-20
C207 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 0.0376f
C208 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.121f
C209 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB 0.103f
C210 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 2.89e-19
C211 RST a_44799_n7920# 4.71e-19
C212 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C213 VDD90 a_32076_6159# 3.14e-19
C214 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 0.415f
C215 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_50151_n2243# 1.46e-19
C216 RST CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 0.00628f
C217 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 3.43e-19
C218 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN 0.0758f
C219 Vdiv99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT 0.126f
C220 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN 1.02e-20
C221 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_47988_n17599# 9.1e-19
C222 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 F2 9.64e-20
C223 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_33519_11196# 1.17e-20
C224 RST CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.00657f
C225 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_53375_1671# 4.52e-20
C226 CLK a_44061_n15627# 0.0105f
C227 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0626f
C228 RST a_45541_n18696# 6.14e-19
C229 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0334f
C230 a_25482_n16632# CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 6.19e-21
C231 VDD100 a_55067_297# 0.0407f
C232 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 a_25625_n6010# 9.09e-19
C233 VDD99 a_31577_n15535# 2.21e-19
C234 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_54187_n16728# 0.0101f
C235 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0948f
C236 CLK_div_105_mag_0.CLK_div_10_mag_1.CLK a_54775_9057# 0.0101f
C237 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 0.128f
C238 VDD96 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_1.IN2 0.408f
C239 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.11f
C240 CLK_div_108_new_mag_0.JK_FF_mag_1.Q a_51957_n6821# 0.0157f
C241 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_32640_6159# 0.0059f
C242 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.0126f
C243 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0622f
C244 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.69f
C245 VDD VDD93 0.314f
C246 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 0.294f
C247 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C248 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 9.67e-20
C249 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_48623_n13424# 0.00747f
C250 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 7.98e-20
C251 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 a_53120_5143# 2.55e-20
C252 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_53850_6284# 1.43e-19
C253 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 8.81e-20
C254 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_22295_5018# 0.0202f
C255 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_48258_n10160# 0.0202f
C256 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 0.00586f
C257 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_54568_5187# 0.0036f
C258 CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 a_53892_n2243# 0.0101f
C259 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 9.62e-20
C260 VDD F0 6.8f
C261 RST CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 4.17e-20
C262 mux_8x1_ibr_0.mux_2x1_ibr_0.I1 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 5.19e-19
C263 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.391f
C264 RST a_23184_n9840# 9.46e-19
C265 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_96_mag_0.JK_FF_mag_3.QB 4.41e-19
C266 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 m3_20882_n11188# 1.63e-21
C267 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_30336_10099# 0.00119f
C268 RST CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 0.044f
C269 RST CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.305f
C270 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 2.81e-20
C271 RST CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 0.293f
C272 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 5.08e-20
C273 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.106f
C274 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 1.71e-21
C275 CLK_div_108_new_mag_0.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.IN2 9.3e-20
C276 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 a_47299_10154# 0.069f
C277 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT a_52385_n13362# 0.198f
C278 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00183f
C279 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_23403_10099# 0.0697f
C280 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 a_23956_n14213# 1.78e-20
C281 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT a_51983_7381# 0.00138f
C282 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.399f
C283 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_53174_n1146# 0.00119f
C284 Vdiv108 a_53255_n5765# 2.79e-20
C285 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 6.82e-19
C286 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_24512_n18723# 0.069f
C287 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 2.61e-19
C288 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 1.53e-19
C289 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.00183f
C290 CLK_div_100_mag_0.CLK_div_10_mag_1.CLK CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 1.48e-20
C291 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0274f
C292 VDD96 a_27496_n2952# 3.14e-19
C293 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.768f
C294 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 1.33e-19
C295 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 4.42e-19
C296 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 3.3e-19
C297 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_54028_n18696# 6.43e-21
C298 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.321f
C299 CLK_div_96_mag_0.JK_FF_mag_3.Q a_29116_398# 6.43e-21
C300 Vdiv100 a_35747_280# 0.00293f
C301 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.999f
C302 CLK_div_96_mag_0.JK_FF_mag_4.Q a_23139_n287# 6.43e-21
C303 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_54509_2768# 0.0731f
C304 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 1f
C305 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.125f
C306 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.122f
C307 RST a_25806_n17626# 0.00549f
C308 RST CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.027f
C309 VDD110 a_45907_n16680# 3.14e-19
C310 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 6.82e-19
C311 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 1.29e-19
C312 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.752f
C313 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 0.00458f
C314 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_29751_n15493# 0.011f
C315 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0948f
C316 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 a_22551_n14504# 0.00765f
C317 a_51486_1671# a_51646_1671# 0.0504f
C318 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 8.16e-20
C319 RST a_29270_n743# 0.00121f
C320 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00544f
C321 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 7.08e-20
C322 a_27939_n17626# a_28099_n17626# 0.0504f
C323 RST CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 0.129f
C324 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_53813_n6862# 0.0203f
C325 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C326 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0343f
C327 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.352f
C328 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 0.892f
C329 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00434f
C330 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 a_50768_2768# 8.64e-19
C331 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00183f
C332 RST a_54978_6284# 6.14e-19
C333 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K 1.41e-20
C334 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_50144_n16724# 0.00335f
C335 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 m3_20882_n11188# 0.00338f
C336 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.76e-19
C337 RST CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 0.188f
C338 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.133f
C339 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 5.13e-19
C340 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB a_21431_n7106# 0.0114f
C341 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 7.55e-19
C342 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00157f
C343 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 2.23e-19
C344 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB a_26636_n8734# 0.0114f
C345 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 9.98e-19
C346 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 4.08f
C347 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 a_46867_7960# 1.29e-22
C348 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.394f
C349 RST a_43872_9057# 4.42e-19
C350 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT a_47760_n15585# 0.00378f
C351 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 1.89e-19
C352 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 a_52951_7381# 0.0096f
C353 RST CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00544f
C354 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.186f
C355 Vdiv108 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.338f
C356 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.321f
C357 a_43591_n5176# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1.17e-20
C358 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 4.33e-19
C359 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_23129_n6009# 0.0731f
C360 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_29680_398# 0.069f
C361 CLK_div_96_mag_0.JK_FF_mag_4.Q a_25122_1919# 0.069f
C362 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 2.29e-19
C363 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 F1 0.413f
C364 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.527f
C365 CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.IN2 a_50353_n9020# 4.9e-20
C366 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00356f
C367 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.013f
C368 dec3x8_ibr_mag_0.and_3_ibr_3.nand3_mag_ibr_0.OUT a_39420_6821# 0.0249f
C369 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB 1.97f
C370 RST CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN 0.0233f
C371 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 6.43e-20
C372 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.122f
C373 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_30317_n18723# 0.012f
C374 RST CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.IN1 0.218f
C375 CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 a_55132_5187# 0.0157f
C376 RST CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00675f
C377 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT a_47905_1671# 0.0202f
C378 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.198f
C379 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_54866_n1102# 0.00372f
C380 CLK_div_96_mag_0.JK_FF_mag_4.Q a_26980_3016# 0.00335f
C381 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 0.631f
C382 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0032f
C383 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT m3_20882_n11188# 0.00434f
C384 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT 0.00183f
C385 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C386 Vdiv99 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I1 0.00437f
C387 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB 0.221f
C388 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 a_45787_574# 0.01f
C389 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 0.0693f
C390 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00169f
C391 VDD110 a_47994_n18696# 3.14e-19
C392 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 a_23956_n14213# 0.0205f
C393 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_48629_1671# 0.00111f
C394 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.0285f
C395 CLK CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.235f
C396 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_36827_n10028# 0.0733f
C397 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_50281_n17599# 0.00335f
C398 CLK_div_90_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 4.85e-20
C399 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_25535_354# 0.00119f
C400 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.00359f
C401 a_54028_n18696# CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 5.94e-20
C402 RST a_52657_2768# 9.66e-19
C403 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.VOUT CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.IN1 0.0103f
C404 RST a_25644_n2996# 0.00243f
C405 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_30163_n17626# 0.00372f
C406 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT 0.16f
C407 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0018f
C408 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0894f
C409 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.994f
C410 Vdiv100 CLK_div_100_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00229f
C411 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT a_47911_2768# 0.0203f
C412 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 0.0998f
C413 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_41284_n14596# 8.95e-19
C414 VDD99 CLK_div_90_mag_0.CLK_div_10_mag_0.CLK 1.08e-20
C415 CLK_div_96_mag_0.JK_FF_mag_4.QB CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 1.34e-19
C416 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00952f
C417 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_44799_n7920# 4.98e-20
C418 RST a_53303_n16728# 0.00256f
C419 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 5.23e-20
C420 CLK_div_96_mag_0.JK_FF_mag_5.Q a_22424_n1833# 0.00939f
C421 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.739f
C422 RST a_53892_n2243# 0.00186f
C423 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT a_51652_2768# 0.0202f
C424 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_41117_n13911# 0.00572f
C425 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 7.97e-19
C426 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_32071_11196# 0.0036f
C427 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_43718_10154# 0.00372f
C428 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.298f
C429 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 0.396f
C430 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.215f
C431 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.0384f
C432 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_26616_n15491# 0.011f
C433 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 9.82e-20
C434 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.0275f
C435 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 4.69e-20
C436 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 1.17f
C437 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.038f
C438 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 1.48e-20
C439 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 8.16e-20
C440 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT 0.266f
C441 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 0.58f
C442 a_22405_n6009# a_22565_n6009# 0.0504f
C443 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK a_39126_n8931# 0.00939f
C444 VDD100 a_53221_2768# 0.00152f
C445 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.333f
C446 RST a_43760_1671# 4.42e-19
C447 RST CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.633f
C448 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.097f
C449 VDD90 a_22301_6115# 0.00752f
C450 CLK a_21841_n6009# 0.00194f
C451 CLK a_48534_5187# 4.86e-19
C452 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 3.84e-20
C453 Vdiv93 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.0555f
C454 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT a_50358_1671# 4.52e-20
C455 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 0.0409f
C456 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.103f
C457 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 CLK 0.149f
C458 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 a_55310_n17599# 0.0157f
C459 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB a_34468_n17626# 0.00695f
C460 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K a_53014_n1146# 8.64e-19
C461 VDD96 a_29801_1733# 0.165f
C462 CLK_div_90_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 1.4e-19
C463 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 a_21431_n7106# 0.069f
C464 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 0.00889f
C465 Vdiv110 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT 2.57e-21
C466 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 0.881f
C467 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.352f
C468 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.235f
C469 VDD100 a_54456_n2199# 3.14e-19
C470 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 2.44e-20
C471 a_50923_n10161# m3_20882_n11188# 4.3e-19
C472 a_26990_11196# a_27150_11196# 0.0504f
C473 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.913f
C474 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_26420_10099# 0.00378f
C475 VDD108 a_48023_n7840# 0.165f
C476 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00183f
C477 VDD100 a_44324_1671# 3.14e-19
C478 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_27227_398# 0.00372f
C479 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_26984_10099# 0.00119f
C480 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 a_44894_2768# 0.0102f
C481 RST CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 0.445f
C482 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 Vdiv110 0.0011f
C483 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_29270_n743# 2.88e-20
C484 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 8.27e-19
C485 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 3.4e-19
C486 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_54781_10154# 1.17e-20
C487 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 2.81e-20
C488 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 a_28267_n7033# 0.0108f
C489 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.0685f
C490 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT 0.00132f
C491 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.291f
C492 a_55310_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0811f
C493 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K a_33583_n16588# 2.75e-21
C494 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.103f
C495 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0129f
C496 CLK_div_96_mag_0.JK_FF_mag_0.QB CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 1.7e-19
C497 CLK_div_108_new_mag_0.CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K 0.00384f
C498 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 a_29144_n8735# 0.0059f
C499 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT a_45899_7960# 0.00138f
C500 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT m3_20882_n11188# 0.00187f
C501 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_47424_n17599# 0.0731f
C502 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.744f
C503 CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 0.0445f
C504 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 Vdiv110 1.96e-19
C505 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_33359_11196# 1.5e-20
C506 RST a_28267_n7033# 3.99e-19
C507 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.159f
C508 VDD a_39420_6265# 2.21e-19
C509 CLK a_43901_n15627# 0.0114f
C510 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.122f
C511 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.742f
C512 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 8.02e-20
C513 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00183f
C514 RST a_44977_n18696# 2.66e-19
C515 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_23706_n2886# 0.0036f
C516 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT 2.57e-20
C517 Vdiv108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT 7.02e-21
C518 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_49488_n13383# 3.04e-20
C519 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 1.85e-19
C520 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_53469_n15631# 2.79e-20
C521 RST CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00412f
C522 VDD100 a_54907_297# 0.234f
C523 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 a_25465_n6010# 9.09e-19
C524 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_54027_n16728# 0.0102f
C525 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.395f
C526 CLK_div_105_mag_0.CLK_div_10_mag_1.CLK a_54615_9057# 0.00939f
C527 CLK_div_108_new_mag_0.JK_FF_mag_1.Q a_51393_n6821# 0.00859f
C528 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_32076_6159# 0.0697f
C529 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.398f
C530 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 0.0343f
C531 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 0.00115f
C532 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.0758f
C533 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K 6.21e-20
C534 RST CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0606f
C535 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 8.56e-20
C536 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 2.92f
C537 F1 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 2.05e-19
C538 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_53286_6240# 0.00119f
C539 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 a_52115_5187# 0.0157f
C540 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.397f
C541 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_48098_n10160# 0.0731f
C542 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C543 CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 a_53732_n2243# 0.0102f
C544 a_51165_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0733f
C545 RST a_22620_n9884# 0.00186f
C546 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.122f
C547 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K 3.03e-20
C548 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_29772_10099# 1.43e-19
C549 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00213f
C550 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.362f
C551 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.999f
C552 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_50447_n18696# 1.41e-20
C553 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.00335f
C554 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0995f
C555 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 0.104f
C556 RST CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 0.00594f
C557 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.103f
C558 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 a_46735_10154# 0.00372f
C559 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0346f
C560 RST CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 0.432f
C561 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 9.37e-19
C562 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I1 0.328f
C563 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT a_52225_n13362# 0.0135f
C564 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB 0.307f
C565 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_22839_10099# 0.0059f
C566 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT a_35747_880# 0.00949f
C567 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_50829_n6865# 2.88e-20
C568 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 CLK_div_96_mag_0.JK_FF_mag_2.QB 0.00139f
C569 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 a_45730_10154# 0.00117f
C570 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_23948_n18723# 0.00372f
C571 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.0659f
C572 VDD96 a_26932_n2952# 3.14e-19
C573 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 0.25f
C574 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.0957f
C575 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 8.16e-20
C576 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.653f
C577 VDD105 a_44282_10154# 3.14e-19
C578 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.16f
C579 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_26965_n18723# 0.0112f
C580 CLK_div_96_mag_0.JK_FF_mag_3.Q a_28552_354# 0.00959f
C581 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0702f
C582 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 9.07e-20
C583 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_53945_2768# 9.1e-19
C584 VDD99 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 0.00114f
C585 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 4.52e-20
C586 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 1.32e-19
C587 VDD110 a_43901_n15627# 2.21e-19
C588 VDD110 a_45343_n16680# 3.14e-19
C589 VDD105 a_45000_9057# 3.14e-19
C590 VDD99 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 2.15e-20
C591 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_0.Q 0.00335f
C592 RST a_25646_n17626# 0.00513f
C593 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.00118f
C594 CLK CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.00364f
C595 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_29187_n15493# 1.43e-19
C596 a_47698_n2243# a_47858_n2243# 0.0504f
C597 VDD96 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.751f
C598 RST a_29110_n743# 0.00141f
C599 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 1.28e-19
C600 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00164f
C601 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.0345f
C602 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB a_54503_1671# 0.00392f
C603 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 3.34e-21
C604 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0718f
C605 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 7.08e-20
C606 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.OUT 0.12f
C607 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_53249_n6862# 1.5e-20
C608 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 1.29e-19
C609 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.66f
C610 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_55020_n2199# 0.0811f
C611 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT 0.00718f
C612 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_46774_n6273# 0.00392f
C613 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0343f
C614 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 1.3e-19
C615 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 2.25e-21
C616 CLK_div_93_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 3.67e-20
C617 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_47134_n2243# 1.46e-19
C618 RST a_54414_6284# 6.14e-19
C619 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 0.244f
C620 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.215f
C621 RST a_55132_5187# 9.66e-19
C622 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN a_42083_n15712# 1.14e-19
C623 CLK Vdiv90 1.28f
C624 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 8.02e-20
C625 CLK_div_96_mag_0.JK_FF_mag_3.Q a_25529_n743# 0.00164f
C626 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 a_51871_n5# 0.0112f
C627 VDD105 a_47835_7960# 6e-19
C628 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB a_26072_n8734# 2.96e-19
C629 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K 9.55e-19
C630 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 0.0011f
C631 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT a_47196_n15629# 0.0732f
C632 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K m3_20882_n11188# 0.00468f
C633 VDD99 a_25806_n17626# 0.00743f
C634 RST CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.312f
C635 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_54978_6284# 0.00372f
C636 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 9.94e-21
C637 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00107f
C638 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 1.58e-20
C639 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 1.82e-19
C640 F0 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I1 0.0112f
C641 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.0147f
C642 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_51205_n7921# 1.82e-21
C643 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_22565_n6009# 9.1e-19
C644 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN 6.88e-21
C645 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 0.124f
C646 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00425f
C647 Vdiv108 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 0.0191f
C648 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_45405_n2199# 0.00378f
C649 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 a_51481_n9064# 2.79e-20
C650 CLK_div_90_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_23691_9000# 0.069f
C651 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.664f
C652 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 4.52e-20
C653 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.466f
C654 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 0.0664f
C655 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 6.51e-19
C656 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 Vdiv110 0.0223f
C657 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 0.0886f
C658 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.398f
C659 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.0485f
C660 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 2.48e-20
C661 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.00864f
C662 VDD99 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 0.00177f
C663 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 0.425f
C664 CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 a_54568_5187# 0.00859f
C665 RST a_24127_10099# 0.00222f
C666 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT a_47341_1671# 4.52e-20
C667 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 a_49276_n17599# 0.00372f
C668 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_54302_n1102# 0.069f
C669 CLK_div_96_mag_0.JK_FF_mag_4.Q a_26820_3016# 0.00789f
C670 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.21f
C671 RST CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.0541f
C672 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_29214_n6271# 3.85e-20
C673 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 0.578f
C674 RST CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0686f
C675 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN 2.47e-20
C676 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 a_26096_3016# 8.64e-19
C677 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.651f
C678 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C679 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_48469_1671# 9.32e-19
C680 a_55067_297# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 3.02e-19
C681 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_36667_n10028# 0.0203f
C682 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_1.IN2 Vdiv99 0.0173f
C683 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C684 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB 9.14e-19
C685 Vdiv99 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK 0.21f
C686 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT 2.18e-21
C687 CLK_div_108_new_mag_0.CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 3.67e-20
C688 RST a_25484_n2996# 0.00243f
C689 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_53333_10154# 0.0036f
C690 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 8.26e-20
C691 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 2.08f
C692 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.122f
C693 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00164f
C694 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_1.IN2 0.00975f
C695 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN 0.00529f
C696 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 9.52e-19
C697 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT a_47751_2768# 0.0733f
C698 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.236f
C699 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.648f
C700 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 1.21e-19
C701 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 8.58e-20
C702 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 0.3f
C703 RST a_52156_n16680# 0.0013f
C704 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 7.24e-19
C705 CLK_div_96_mag_0.JK_FF_mag_5.Q a_22264_n1833# 0.0101f
C706 RST a_53732_n2243# 0.00169f
C707 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT a_51492_2768# 0.0731f
C708 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 0.0131f
C709 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_47430_n18696# 0.00939f
C710 RST CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.0843f
C711 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.105f
C712 F1 a_36042_6821# 4.46e-19
C713 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_26052_n15491# 1.43e-19
C714 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 6.3e-20
C715 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.16f
C716 CLK CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 0.00343f
C717 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_43872_9057# 4.52e-20
C718 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.359f
C719 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 7.72e-21
C720 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.16f
C721 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK a_38966_n8931# 0.0101f
C722 VDD100 a_52657_2768# 0.00152f
C723 RST a_28828_1497# 4.93e-19
C724 VDD96 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 1.21f
C725 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.359f
C726 RST a_45603_n5176# 0.00173f
C727 RST CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 3.69e-19
C728 CLK CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.272f
C729 CLK a_21277_n6009# 0.00207f
C730 CLK a_47970_5143# 4.68e-19
C731 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT a_53738_n1102# 5.94e-20
C732 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_52161_n19793# 0.0112f
C733 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.109f
C734 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_31731_n16632# 1.46e-19
C735 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00157f
C736 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 0.00195f
C737 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.321f
C738 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB a_34308_n17626# 0.00696f
C739 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 a_54746_n17599# 0.00859f
C740 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB 0.25f
C741 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 4.2e-19
C742 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 6.87e-20
C743 CLK CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.00293f
C744 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 1.74e-19
C745 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K a_47030_n16726# 8.64e-19
C746 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 a_34896_n15539# 2.79e-20
C747 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.00129f
C748 CLK dec3x8_ibr_mag_0.and_3_ibr_4.nand3_mag_ibr_0.OUT 0.00278f
C749 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0995f
C750 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB m3_20882_n11188# 0.00466f
C751 CLK CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.414f
C752 CLK_div_90_mag_0.CLK_div_10_mag_0.CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.419f
C753 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 0.0703f
C754 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00174f
C755 a_50763_n10161# m3_20882_n11188# 4.3e-19
C756 a_46400_n9019# CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 4.52e-20
C757 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.103f
C758 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.VOUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.0017f
C759 dec3x8_ibr_mag_0.and_3_ibr_3.nand3_mag_ibr_0.OUT dec3x8_ibr_mag_0.and_3_ibr_7.nand3_mag_ibr_0.OUT 0.00141f
C760 VDD108 a_44799_n7920# 5.92e-19
C761 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT 0.999f
C762 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 6.57e-19
C763 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00541f
C764 VDD100 a_43760_1671# 3.56e-19
C765 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_26663_398# 0.069f
C766 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 8.02e-19
C767 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_26420_10099# 1.43e-19
C768 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 a_44734_2768# 0.0101f
C769 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.741f
C770 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.647f
C771 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C772 VDD96 CLK_div_96_mag_0.JK_FF_mag_0.QB 0.926f
C773 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_52951_7381# 8.17e-21
C774 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_29110_n743# 9.1e-19
C775 Vdiv96 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 0.0995f
C776 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_54621_10154# 1.5e-20
C777 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_47430_n18696# 1.41e-20
C778 CLK_div_108_new_mag_0.JK_FF_mag_1.Q CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K 0.0372f
C779 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.122f
C780 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 1e-19
C781 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_26770_n16588# 0.00378f
C782 a_54746_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.00964f
C783 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 4.84e-19
C784 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K a_33019_n16588# 5.58e-22
C785 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.00154f
C786 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_0.OUT CLK_div_96_mag_0.JK_FF_mag_3.Q 1.45e-19
C787 VDD96 a_30398_n699# 3.14e-19
C788 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 a_28580_n8735# 0.0697f
C789 VDD90 a_31352_6115# 2.21e-19
C790 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN 0.00326f
C791 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_47264_n17599# 0.0202f
C792 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT 0.00132f
C793 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C794 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_32795_11196# 0.0203f
C795 RST a_26343_n7107# 8.67e-19
C796 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN a_52839_n5# 0.069f
C797 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 5.74e-20
C798 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.768f
C799 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.IN2 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_1.IN2 0.00212f
C800 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 a_54669_2768# 0.00335f
C801 a_45458_2768# a_45618_2768# 0.0504f
C802 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_48783_n13424# 8.5e-20
C803 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT a_45927_6284# 2.05e-19
C804 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN 4.29e-20
C805 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 a_24901_n6010# 0.00108f
C806 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_53463_n16728# 0.00789f
C807 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.442f
C808 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.398f
C809 CLK_div_105_mag_0.CLK_div_10_mag_1.CLK a_54051_9057# 6.43e-21
C810 CLK_div_108_new_mag_0.JK_FF_mag_1.Q a_50829_n6865# 0.0101f
C811 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 m3_20882_n11188# 8.8e-19
C812 CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C813 a_43831_7266# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00239f
C814 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 2.81e-20
C815 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB a_51486_1671# 0.00392f
C816 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT a_26250_1919# 0.0202f
C817 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_50105_n6865# 1.46e-19
C818 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 3.27e-20
C819 VDD90 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 0.106f
C820 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C821 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.0205f
C822 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0042f
C823 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 a_50903_n5# 0.0105f
C824 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 a_50269_6240# 2.79e-20
C825 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_0.OUT 0.0884f
C826 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 a_25122_1919# 4.52e-20
C827 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 a_51551_5187# 0.00859f
C828 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0343f
C829 a_27342_n1855# CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 4.52e-20
C830 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_47534_n10160# 9.1e-19
C831 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_43757_n6273# 0.00392f
C832 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.0685f
C833 CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 a_53168_n2243# 0.00789f
C834 a_51005_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0203f
C835 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0106f
C836 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB 0.348f
C837 RST a_22460_n9884# 8.64e-19
C838 RST CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.155f
C839 RST a_29307_n1855# 3.83e-19
C840 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_29208_10099# 0.011f
C841 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.122f
C842 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_50287_n18696# 1.86e-20
C843 VDD93 a_37801_n8887# 3.6e-19
C844 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C845 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 0.0215f
C846 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 Vdiv90 0.274f
C847 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0346f
C848 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 0.0512f
C849 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 0.622f
C850 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 a_45241_n10160# 0.00335f
C851 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_23748_n9840# 0.00372f
C852 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_50669_n6865# 9.1e-19
C853 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 a_45570_10154# 0.00164f
C854 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 8.98e-19
C855 a_25122_1919# CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 3.98e-19
C856 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 a_38454_6821# 0.00297f
C857 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.321f
C858 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.00395f
C859 CLK_div_108_new_mag_0.JK_FF_mag_1.Q CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0635f
C860 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_23249_11196# 8.64e-19
C861 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.768f
C862 VDD105 a_43718_10154# 3.14e-19
C863 CLK_div_100_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.00154f
C864 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 1.34f
C865 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 0.0215f
C866 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K 0.0685f
C867 CLK_div_96_mag_0.JK_FF_mag_3.Q a_28392_354# 0.0101f
C868 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C869 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.28f
C870 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_53785_2768# 2.88e-20
C871 VDD105 a_44436_9057# 3.14e-19
C872 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 0.133f
C873 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.431f
C874 RST a_25082_n17626# 0.00211f
C875 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.321f
C876 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 0.0444f
C877 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_28623_n15537# 0.00119f
C878 VDD93 CLK_div_90_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 2.2e-19
C879 CLK dec3x8_ibr_mag_0.and_3_ibr_5.IN3 0.00218f
C880 RST a_28546_n743# 0.00254f
C881 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 1.05e-20
C882 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB a_53939_1671# 3.33e-19
C883 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 0.442f
C884 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 2.4f
C885 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN 0.0104f
C886 RST a_23145_810# 0.00103f
C887 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00162f
C888 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 0.055f
C889 F1 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.OUT 0.00227f
C890 RST CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.255f
C891 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_55156_n18696# 0.00372f
C892 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_53089_n6862# 1.17e-20
C893 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K a_31451_n17626# 5.54e-20
C894 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_54456_n2199# 0.00964f
C895 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 8.16e-20
C896 RST CLK_div_96_mag_0.JK_FF_mag_4.Q 0.161f
C897 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00357f
C898 CLK_div_108_new_mag_0.JK_FF_mag_1.Q CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 1.48e-20
C899 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 0.0502f
C900 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_33204_6159# 0.00118f
C901 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.644f
C902 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.231f
C903 RST a_53850_6284# 2.78e-19
C904 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 2.81e-20
C905 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0857f
C906 RST a_54568_5187# 9.41e-19
C907 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.00254f
C908 CLK a_33405_7558# 1.88e-19
C909 CLK_div_96_mag_0.JK_FF_mag_5.Q a_22011_n287# 0.069f
C910 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00183f
C911 CLK_div_96_mag_0.JK_FF_mag_3.Q a_25369_n743# 0.00117f
C912 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB a_25508_n8734# 3.25e-19
C913 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.0622f
C914 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_54414_6284# 0.069f
C915 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT a_47036_n15629# 0.0203f
C916 VDD99 a_25646_n17626# 0.00305f
C917 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K 9.55e-19
C918 VDD99 a_30315_n15493# 3.56e-19
C919 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT Vdiv100 0.0251f
C920 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 a_47332_n5176# 3.6e-22
C921 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_22405_n6009# 2.88e-20
C922 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.00335f
C923 Vdiv108 a_37999_280# 0.0024f
C924 RST CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 0.592f
C925 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_44841_n2243# 0.0733f
C926 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 0.397f
C927 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00305f
C928 RST CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.00337f
C929 a_43760_1671# CLK_div_100_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 2.1e-20
C930 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 a_53168_n2243# 0.00164f
C931 RST CLK_div_96_mag_0.JK_FF_mag_5.Q 0.0201f
C932 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT a_48629_1671# 0.0203f
C933 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0228f
C934 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 6.05e-19
C935 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_26226_n9831# 0.00378f
C936 CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 a_53286_6240# 2.79e-20
C937 RST a_54057_10154# 8.64e-19
C938 CLK CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00461f
C939 CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 a_54004_5143# 0.0101f
C940 RST a_23967_10099# 0.00159f
C941 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 a_48712_n17599# 0.069f
C942 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00808f
C943 CLK_div_96_mag_0.JK_FF_mag_4.Q a_26256_3016# 0.0102f
C944 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.233f
C945 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C946 RST a_24133_11196# 0.00325f
C947 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.121f
C948 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 1.47e-19
C949 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 1.03f
C950 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_22466_n8743# 0.00378f
C951 CLK_div_108_new_mag_0.JK_FF_mag_1.Q CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 6.27e-22
C952 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00157f
C953 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_47905_1671# 3.12e-19
C954 a_54907_297# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 9.21e-20
C955 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_36103_n10028# 1.5e-20
C956 a_24116_n1789# CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 4.52e-20
C957 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0894f
C958 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 0.442f
C959 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_22455_5018# 1.46e-19
C960 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.529f
C961 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.182f
C962 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.179f
C963 a_45899_7960# CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN 5.1e-20
C964 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 0.0343f
C965 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C966 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.21f
C967 RST a_24270_n2886# 0.0013f
C968 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 3.9f
C969 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 a_30315_n15493# 0.00372f
C970 VDD93 Vdiv100 1.65e-19
C971 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT a_47187_2768# 0.00378f
C972 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 2.93e-20
C973 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 0.00152f
C974 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 4.42e-19
C975 RST a_50874_n15583# 3.68e-20
C976 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 a_31128_n7028# 0.00479f
C977 RST a_51592_n16680# 0.00129f
C978 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT 0.00157f
C979 VDD100 a_54663_1671# 0.00752f
C980 RST a_53168_n2243# 0.00186f
C981 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.88f
C982 F0 Vdiv100 0.0242f
C983 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT a_50928_2768# 9.1e-19
C984 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 a_23510_n15620# 0.00208f
C985 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.268f
C986 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT a_47914_n16726# 2.88e-20
C987 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_46081_5187# 0.00372f
C988 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_47270_n18696# 0.0101f
C989 CLK CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 0.0215f
C990 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 a_29087_8532# 0.0134f
C991 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_25488_n15535# 0.00119f
C992 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 1.83e-19
C993 a_47092_6240# a_47252_6240# 0.0504f
C994 CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 9.92e-20
C995 RST CLK_div_105_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.021f
C996 CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 a_30060_9000# 7.48e-20
C997 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.652f
C998 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 0.159f
C999 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 2.8e-19
C1000 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.109f
C1001 RST a_45039_n5176# 0.00113f
C1002 a_43751_n5176# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.46e-19
C1003 CLK a_47810_5143# 4.68e-19
C1004 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_44170_2768# 0.069f
C1005 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0147f
C1006 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT a_44779_n16724# 2.88e-20
C1007 CLK_div_96_mag_0.JK_FF_mag_2.Q CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.267f
C1008 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 1.4e-21
C1009 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB a_33744_n17626# 0.00964f
C1010 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 3.06f
C1011 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 0.388f
C1012 CLK a_53129_n19793# 2.22e-19
C1013 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 6.35e-19
C1014 Vdiv96 Vdiv108 0.00317f
C1015 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K a_45907_n16680# 1.44e-21
C1016 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0378f
C1017 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.107f
C1018 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.00183f
C1019 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_51193_n19793# 0.0105f
C1020 VDD100 a_53732_n2243# 2.21e-19
C1021 CLK CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT 1.46e-19
C1022 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 2.53f
C1023 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 4.01e-20
C1024 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB a_48469_1671# 0.00392f
C1025 a_50199_n10117# m3_20882_n11188# 4.41e-19
C1026 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_1.IN2 a_35747_n1822# 0.00372f
C1027 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 8.51e-22
C1028 VDD100 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 3.91e-19
C1029 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00167f
C1030 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 1.99e-21
C1031 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 6.72e-20
C1032 a_31291_n17626# a_31451_n17626# 0.0504f
C1033 VDD99 a_28828_1497# 2.13e-20
C1034 VDD99 a_36742_n16592# 3.14e-19
C1035 a_53780_n10161# a_53940_n10161# 0.0504f
C1036 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.916f
C1037 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.0758f
C1038 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 a_44170_2768# 0.00859f
C1039 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_25856_10099# 0.011f
C1040 CLK_div_100_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 4.85e-20
C1041 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_28546_n743# 0.0731f
C1042 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 6.12e-21
C1043 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.121f
C1044 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 0.0147f
C1045 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_47270_n18696# 1.86e-20
C1046 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_54057_10154# 0.0203f
C1047 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB 0.00541f
C1048 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_26206_n16632# 0.0733f
C1049 Vdiv108 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 1.04e-19
C1050 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_0.OUT a_26974_1919# 0.0203f
C1051 VDD96 a_29834_n699# 3.14e-19
C1052 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.359f
C1053 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT 1.2e-19
C1054 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 a_48023_n7840# 0.0134f
C1055 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0836f
C1056 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1f
C1057 dec3x8_ibr_mag_0.and_3_ibr_3.nand3_mag_ibr_0.OUT F0 0.00326f
C1058 CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.107f
C1059 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_32635_11196# 0.0733f
C1060 RST a_26183_n7107# 7.2e-19
C1061 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 7.24e-19
C1062 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00118f
C1063 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 a_27180_n15491# 0.00372f
C1064 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 a_50903_n5# 2.48e-19
C1065 CLK a_44619_n16724# 6.8e-19
C1066 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_36588_n15495# 0.0114f
C1067 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 a_54509_2768# 0.00789f
C1068 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_48623_n13424# 1.32e-19
C1069 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.0592f
C1070 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00233f
C1071 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.038f
C1072 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK a_36103_n10028# 0.00164f
C1073 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 a_31177_7256# 0.01f
C1074 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 a_24337_n6010# 0.00108f
C1075 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 4.2e-19
C1076 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 1.82e-19
C1077 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_53303_n16728# 0.00335f
C1078 VDD110 a_53129_n19793# 3.14e-19
C1079 CLK_div_108_new_mag_0.JK_FF_mag_1.Q a_50669_n6865# 0.0102f
C1080 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 9.22e-20
C1081 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.122f
C1082 a_43671_7266# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00261f
C1083 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 6.04e-20
C1084 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB a_29862_n9832# 0.0811f
C1085 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT a_25686_1919# 4.52e-20
C1086 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB a_50922_1671# 3.25e-19
C1087 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 0.018f
C1088 VDD Vdiv105 0.429f
C1089 CLK_div_96_mag_0.JK_FF_mag_5.QB CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 1.38e-19
C1090 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 8.26e-20
C1091 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 a_50987_5143# 0.0101f
C1092 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 8.59e-20
C1093 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_47374_n10160# 2.88e-20
C1094 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_53280_5143# 1.46e-19
C1095 CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 a_53008_n2243# 0.00335f
C1096 a_50441_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 1.5e-20
C1097 a_51005_n17599# a_51165_n17599# 0.0504f
C1098 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0013f
C1099 VDD90 a_33519_11196# 0.0132f
C1100 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.338f
C1101 RST a_28743_n1899# 0.00182f
C1102 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0017f
C1103 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_28644_10099# 0.00118f
C1104 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.1f
C1105 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.321f
C1106 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 1.29e-19
C1107 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 0.109f
C1108 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_49122_n18696# 0.0114f
C1109 VDD93 a_37237_n8887# 3.18e-19
C1110 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 1.03f
C1111 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 a_33405_7558# 0.019f
C1112 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 a_45612_1671# 0.0101f
C1113 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 a_23510_n15620# 0.0177f
C1114 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.0635f
C1115 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 a_45081_n10160# 0.00789f
C1116 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_23184_n9840# 0.069f
C1117 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_50105_n6865# 0.0731f
C1118 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 a_38294_6821# 0.00699f
C1119 VDD96 a_26208_n2996# 2.21e-19
C1120 VDD105 a_54978_6284# 3.56e-19
C1121 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00183f
C1122 a_50868_n16724# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 5.49e-20
C1123 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT m3_20882_n11188# 1.87e-19
C1124 a_43901_n15627# a_44061_n15627# 0.0504f
C1125 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 0.11f
C1126 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 a_45724_9057# 0.0101f
C1127 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 0.0777f
C1128 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 a_29708_n8735# 0.00118f
C1129 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_26368_n2996# 8.64e-19
C1130 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 0.00233f
C1131 CLK_div_105_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 6.89e-19
C1132 VDD105 a_43872_9057# 3.56e-19
C1133 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.VOUT 0.867f
C1134 RST a_24922_n17626# 0.0019f
C1135 VDD110 a_44619_n16724# 2.21e-19
C1136 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 0.343f
C1137 CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_99_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.124f
C1138 RST a_29187_n15493# 3.08e-20
C1139 RST a_28386_n743# 0.00359f
C1140 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB a_53375_1671# 2.96e-19
C1141 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0343f
C1142 RST a_22985_810# 0.00144f
C1143 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 m3_20882_n11188# 0.00141f
C1144 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN m3_20882_n11188# 4.94e-19
C1145 F2 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 3.66e-19
C1146 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0501f
C1147 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 7.08e-20
C1148 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_54592_n18696# 0.069f
C1149 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_53892_n2243# 0.00696f
C1150 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_32640_6159# 0.011f
C1151 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.00335f
C1152 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_53464_n18696# 1.41e-20
C1153 VDD105 a_54781_10154# 0.0132f
C1154 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.857f
C1155 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00668f
C1156 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.23f
C1157 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.0835f
C1158 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.122f
C1159 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C1160 RST a_54004_5143# 0.00186f
C1161 a_30342_11196# a_30502_11196# 0.0504f
C1162 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_55020_n2199# 0.00372f
C1163 CLK a_33245_7558# 1.4e-19
C1164 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.00568f
C1165 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.768f
C1166 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB a_24944_n8778# 0.00392f
C1167 RST CLK_div_108_new_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.00333f
C1168 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00776f
C1169 VDD99 a_25082_n17626# 2.21e-19
C1170 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 a_51983_7381# 0.0112f
C1171 VDD99 a_29751_n15493# 3.14e-19
C1172 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 3.28e-19
C1173 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.159f
C1174 VDD dec3x8_ibr_mag_0.and_3_ibr_2.nand3_mag_ibr_0.OUT 0.764f
C1175 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.00602f
C1176 CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN a_22718_8532# 0.132f
C1177 a_43591_n5176# a_43751_n5176# 0.0504f
C1178 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 a_46768_n5176# 1.86e-20
C1179 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 1.82e-19
C1180 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 0.00152f
C1181 a_30060_9000# CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 1.71e-20
C1182 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C1183 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_44681_n2243# 0.0203f
C1184 RST CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 0.428f
C1185 VDD99 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 2.2e-20
C1186 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 1.08f
C1187 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_0.QB 4.51e-20
C1188 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT 0.00157f
C1189 RST CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.IN1 0.226f
C1190 Vdiv110 CLK_div_100_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 4.61e-19
C1191 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00732f
C1192 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 a_53008_n2243# 0.00117f
C1193 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT a_48469_1671# 0.0732f
C1194 VDD99 CLK_div_96_mag_0.JK_FF_mag_4.Q 0.301f
C1195 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_45449_n6273# 0.00372f
C1196 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.322f
C1197 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_25662_n9875# 0.0733f
C1198 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 8.64e-20
C1199 RST a_53897_10154# 0.00186f
C1200 Vdiv96 Vdiv93 0.00698f
C1201 CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 a_53844_5143# 0.0102f
C1202 RST a_23403_10099# 5.71e-19
C1203 CLK_div_96_mag_0.JK_FF_mag_4.Q a_26096_3016# 0.0101f
C1204 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 0.313f
C1205 VDD96 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.999f
C1206 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.16f
C1207 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C1208 RST a_23973_11196# 0.00302f
C1209 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_28093_n18723# 0.0697f
C1210 CLK_div_108_new_mag_0.JK_FF_mag_0.QB CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K 5.16e-20
C1211 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_21902_n8787# 0.0732f
C1212 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_47341_1671# 7.4e-19
C1213 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.654f
C1214 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_35943_n10028# 1.17e-20
C1215 CLK CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 1.05e-19
C1216 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_31737_n15535# 1.16e-20
C1217 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 0.875f
C1218 RST a_52293_n17599# 0.00122f
C1219 dec3x8_ibr_mag_0.and_3_ibr_7.nand3_mag_ibr_0.OUT Vdiv 0.00224f
C1220 CLK_div_96_mag_0.JK_FF_mag_5.QB CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_0.OUT 0.343f
C1221 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0319f
C1222 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 1.96f
C1223 RST a_23706_n2886# 0.00131f
C1224 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.647f
C1225 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.802f
C1226 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.109f
C1227 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 a_29751_n15493# 0.069f
C1228 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 a_51486_1671# 2.79e-20
C1229 VDD99 CLK_div_96_mag_0.JK_FF_mag_5.Q 0.0839f
C1230 RST CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.0172f
C1231 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00262f
C1232 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN 5.47e-20
C1233 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 8.28e-20
C1234 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_52003_n2199# 0.0811f
C1235 a_33652_n13270# a_33812_n13270# 0.186f
C1236 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 2.48e-20
C1237 Vdiv90 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 2.08e-19
C1238 CLK CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00433f
C1239 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C1240 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C1241 RST a_51028_n16724# 0.00216f
C1242 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.338f
C1243 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 2.37f
C1244 VDD100 a_54503_1671# 2.66e-19
C1245 RST a_53008_n2243# 0.00186f
C1246 VDD108 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.392f
C1247 VDD108 a_45603_n5176# 0.00149f
C1248 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT a_50768_2768# 2.88e-20
C1249 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0894f
C1250 RST a_48148_n17599# 0.00211f
C1251 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT a_47754_n16726# 9.1e-19
C1252 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_45517_5187# 0.069f
C1253 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_46105_n18696# 0.069f
C1254 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_47902_n6273# 4.52e-20
C1255 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 0.124f
C1256 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_32794_5062# 0.00378f
C1257 VDD93 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 0.12f
C1258 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00118f
C1259 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.002f
C1260 a_30187_6159# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 4.52e-20
C1261 CLK a_44799_6284# 6.43e-21
C1262 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 F0 0.0552f
C1263 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0698f
C1264 RST a_35614_n16636# 0.00162f
C1265 a_39684_n10028# a_39844_n10028# 0.0504f
C1266 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.104f
C1267 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.00252f
C1268 CLK a_47246_5143# 0.00111f
C1269 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.122f
C1270 a_25375_354# a_25535_354# 0.0504f
C1271 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_43606_2768# 0.00372f
C1272 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB 1.76e-21
C1273 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 0.00637f
C1274 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 3.61e-20
C1275 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT a_44619_n16724# 9.1e-19
C1276 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 1.16f
C1277 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB a_33180_n17626# 0.0811f
C1278 VDD96 a_30435_n1855# 3.56e-19
C1279 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 1.23f
C1280 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.012f
C1281 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.25f
C1282 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K a_45343_n16680# 4.96e-22
C1283 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 a_27144_10099# 3.69e-19
C1284 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 2.48e-19
C1285 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.0622f
C1286 VDD100 a_53168_n2243# 0.00299f
C1287 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 1.94f
C1288 CLK a_51647_n10161# 0.00117f
C1289 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB a_47905_1671# 3.25e-19
C1290 a_49635_n10117# m3_20882_n11188# 4.57e-19
C1291 VDD mux_8x1_ibr_0.mux_2x1_ibr_0.I1 0.422f
C1292 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_1.IN2 a_35184_n1822# 0.069f
C1293 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 0.109f
C1294 a_21995_n7106# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB 5e-20
C1295 VDD100 a_39580_6821# 4.47e-19
C1296 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 0.857f
C1297 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 2.76e-19
C1298 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 0.00173f
C1299 VDD100 CLK_div_105_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00149f
C1300 VDD99 a_36178_n16592# 3.14e-19
C1301 RST CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.112f
C1302 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 6.63e-19
C1303 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_53939_1671# 0.0697f
C1304 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.3f
C1305 VDD110 a_49276_n17599# 0.00152f
C1306 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_51758_9057# 0.00876f
C1307 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_2.OUT CLK_div_96_mag_0.JK_FF_mag_4.QB 0.103f
C1308 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_36827_n10028# 8.64e-19
C1309 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 3.83e-19
C1310 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_23184_n9840# 0.00378f
C1311 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_25292_10099# 0.00118f
C1312 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 a_43606_2768# 0.0157f
C1313 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_51011_n18696# 1.25e-20
C1314 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_28386_n743# 0.0202f
C1315 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_53897_10154# 0.0733f
C1316 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_46105_n18696# 0.0114f
C1317 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 2.89e-19
C1318 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 1.65f
C1319 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.121f
C1320 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_26046_n16632# 0.0203f
C1321 VDD93 a_36202_6821# 0.00167f
C1322 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB a_47911_2768# 0.00695f
C1323 CLK_div_96_mag_0.JK_FF_mag_4.QB CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00182f
C1324 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_0.OUT a_26814_1919# 0.0732f
C1325 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 6.62e-20
C1326 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.122f
C1327 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 0.00586f
C1328 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 9.5e-19
C1329 VDD96 a_23869_810# 0.00108f
C1330 VDD110 a_45131_n17599# 0.00101f
C1331 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 0.647f
C1332 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_32071_11196# 0.00378f
C1333 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 2.21e-20
C1334 RST a_25619_n7107# 3.98e-19
C1335 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN a_54907_297# 2.85e-20
C1336 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT 6.2e-20
C1337 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0147f
C1338 RST CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 0.0232f
C1339 CLK_div_108_new_mag_0.JK_FF_mag_0.QB CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.0592f
C1340 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 a_26616_n15491# 0.069f
C1341 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 1.23e-19
C1342 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 2.51e-19
C1343 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_51803_n5724# 0.00372f
C1344 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.00123f
C1345 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_36024_n15495# 2.96e-19
C1346 CLK a_44055_n16724# 0.00253f
C1347 VDD96 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 0.656f
C1348 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 a_53945_2768# 0.0102f
C1349 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_22418_n2930# 1.46e-19
C1350 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.343f
C1351 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 1.54e-21
C1352 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.283f
C1353 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 0.397f
C1354 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK a_35943_n10028# 0.00117f
C1355 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB 0.179f
C1356 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.768f
C1357 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 0.0138f
C1358 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 3.7f
C1359 CLK_div_108_new_mag_0.JK_FF_mag_1.Q a_50105_n6865# 0.00789f
C1360 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.129f
C1361 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_24307_5062# 0.00372f
C1362 VDD99 F1 0.342f
C1363 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.647f
C1364 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB a_29298_n9832# 0.00964f
C1365 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB a_50358_1671# 2.96e-19
C1366 CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 9.83e-19
C1367 VDD100 F1 0.00799f
C1368 VDD93 a_29862_n9832# 3.14e-19
C1369 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 7.3e-19
C1370 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 8.51e-22
C1371 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 a_50827_5143# 0.0102f
C1372 a_48832_n1102# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 4.52e-20
C1373 a_50281_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 1.17e-20
C1374 CLK_div_96_mag_0.JK_FF_mag_4.QB a_26663_398# 2.05e-20
C1375 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 0.0275f
C1376 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_29054_11196# 0.069f
C1377 VDD90 a_33359_11196# 0.00888f
C1378 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.107f
C1379 RST CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.305f
C1380 RST a_28583_n1899# 0.00242f
C1381 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.00139f
C1382 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 2.52e-20
C1383 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT a_26980_3016# 1.17e-20
C1384 VDD96 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.IN1 0.661f
C1385 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_48558_n18696# 2.96e-19
C1386 VDD93 a_36673_n8887# 3.18e-19
C1387 Vdiv93 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 7.46e-20
C1388 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 0.275f
C1389 RST CLK_div_100_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.021f
C1390 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 a_45452_1671# 0.00939f
C1391 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 6.62e-20
C1392 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.392f
C1393 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN 0.00162f
C1394 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 a_44517_n10160# 0.0102f
C1395 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT Vdiv110 0.00562f
C1396 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 0.0693f
C1397 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_49945_n6865# 0.0202f
C1398 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 a_45730_10154# 0.00335f
C1399 CLK_div_105_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 4.85e-20
C1400 VDD105 a_54414_6284# 3.14e-19
C1401 VDD105 a_55132_5187# 3.14e-19
C1402 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 a_45564_9057# 0.00939f
C1403 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 1.3f
C1404 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 2.81e-20
C1405 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 a_29144_n8735# 0.011f
C1406 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 1.99e-19
C1407 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_53897_10154# 8.64e-19
C1408 VDD93 a_28268_n6266# 3.14e-19
C1409 RST a_24358_n17626# 7.06e-19
C1410 a_53813_n6862# a_53973_n6862# 0.0504f
C1411 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_53819_n5721# 0.00378f
C1412 RST a_27381_n699# 0.00186f
C1413 a_53463_n16728# CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 7.56e-21
C1414 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.321f
C1415 a_51604_10154# a_51764_10154# 0.0504f
C1416 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB a_52811_1671# 0.0114f
C1417 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT Vdiv99 0.0331f
C1418 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.429f
C1419 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.00975f
C1420 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.231f
C1421 a_47835_7960# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 7.43e-22
C1422 a_29862_n9832# m3_20882_n11188# 2.96e-19
C1423 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 2.03e-20
C1424 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_53732_n2243# 0.00695f
C1425 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 Vdiv110 0.00536f
C1426 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 3.84e-20
C1427 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_32076_6159# 1.43e-19
C1428 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 0.0314f
C1429 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_53304_n18696# 1.86e-20
C1430 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 2.45e-22
C1431 VDD105 a_54621_10154# 0.00892f
C1432 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB 1.96f
C1433 RST a_53844_5143# 0.00169f
C1434 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 0.9f
C1435 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 0.00212f
C1436 CLK a_30209_7256# 1.71e-20
C1437 F0 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 2.08e-19
C1438 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_54456_n2199# 0.069f
C1439 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 5.7e-19
C1440 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 3.79e-19
C1441 Vdiv105 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I1 1.08e-19
C1442 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.0248f
C1443 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB 2f
C1444 CLK_div_96_mag_0.JK_FF_mag_3.QB CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.343f
C1445 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 a_51015_7381# 0.00929f
C1446 VDD99 a_29187_n15493# 3.14e-19
C1447 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.26f
C1448 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 0.648f
C1449 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 a_46608_n5176# 2.55e-20
C1450 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_44885_n6273# 4.52e-20
C1451 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.289f
C1452 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 0.622f
C1453 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB 1.34e-19
C1454 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_29772_10099# 0.0202f
C1455 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 a_55156_n18696# 0.069f
C1456 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.0948f
C1457 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.652f
C1458 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 a_49789_n9020# 0.069f
C1459 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_44117_n2243# 1.5e-20
C1460 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 1.99e-19
C1461 Vdiv105 CLK_div_105_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 0.0301f
C1462 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.018f
C1463 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 Vdiv110 0.0434f
C1464 CLK CLK_div_96_mag_0.JK_FF_mag_3.Q 0.0187f
C1465 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT a_47905_1671# 0.00378f
C1466 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_44885_n6273# 0.069f
C1467 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_25502_n9875# 0.0203f
C1468 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.00403f
C1469 RST a_53333_10154# 9.41e-19
C1470 RST a_53375_1671# 6.14e-19
C1471 CLK CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 0.0013f
C1472 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 a_31506_5018# 0.00164f
C1473 CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 a_53280_5143# 0.00789f
C1474 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.397f
C1475 RST a_22839_10099# 5.16e-19
C1476 CLK_div_96_mag_0.JK_FF_mag_4.Q a_25532_3016# 0.00859f
C1477 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT 0.00157f
C1478 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 0.0379f
C1479 RST a_23409_11196# 0.00232f
C1480 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_27529_n18723# 0.0059f
C1481 VDD90 RST 3.32f
C1482 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN a_47835_7960# 0.069f
C1483 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT 2.74e-20
C1484 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_21742_n8787# 0.0203f
C1485 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C1486 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.233f
C1487 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_46777_1671# 7.4e-19
C1488 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.92f
C1489 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 0.275f
C1490 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 2.14e-21
C1491 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 0.00761f
C1492 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT 6.99e-20
C1493 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN 0.124f
C1494 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_31577_n15535# 1.49e-20
C1495 RST a_51729_n17599# 0.00119f
C1496 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.652f
C1497 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_54781_10154# 0.0202f
C1498 RST a_23142_n2930# 0.00215f
C1499 CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN a_24391_n20290# 0.132f
C1500 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_55156_n18696# 0.0114f
C1501 VDD108 a_39580_6821# 2.34e-19
C1502 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00118f
C1503 RST CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 0.105f
C1504 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_51439_n2199# 0.00964f
C1505 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 8.11e-19
C1506 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 0.0126f
C1507 CLK CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 0.417f
C1508 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 4.73e-19
C1509 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 9.62e-20
C1510 RST a_50868_n16724# 0.00199f
C1511 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0064f
C1512 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0622f
C1513 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 1.7e-19
C1514 VDD100 a_53939_1671# 3.14e-19
C1515 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT 0.00243f
C1516 VDD108 a_45039_n5176# 0.00149f
C1517 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00356f
C1518 RST a_52003_n2199# 9.66e-19
C1519 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 0.0582f
C1520 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN 0.423f
C1521 RST a_47988_n17599# 0.00195f
C1522 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT a_47190_n16726# 0.0731f
C1523 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_45541_n18696# 6.06e-21
C1524 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_47338_n6273# 0.0202f
C1525 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.642f
C1526 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 0.116f
C1527 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_32230_5018# 0.0733f
C1528 VDD108 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 5.23e-19
C1529 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 3.84e-20
C1530 F0 Vdiv 0.794f
C1531 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.105f
C1532 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 0.391f
C1533 RST CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 0.59f
C1534 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 a_30881_n18723# 0.069f
C1535 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0881f
C1536 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K a_30915_n13291# 2.5e-19
C1537 CLK a_44235_6240# 0.00939f
C1538 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 2.96e-19
C1539 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 2.03e-20
C1540 RST a_35454_n16636# 0.00176f
C1541 CLK_div_96_mag_0.JK_FF_mag_2.Q CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 9.71e-20
C1542 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_35949_n8931# 8.64e-19
C1543 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00164f
C1544 RST CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.254f
C1545 CLK a_47086_5143# 0.00111f
C1546 Vdiv110 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 2.4e-20
C1547 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.IN2 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT 0.12f
C1548 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0399f
C1549 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT a_44055_n16724# 0.0731f
C1550 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 0.00761f
C1551 VDD96 a_29871_n1855# 3.14e-19
C1552 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT 0.122f
C1553 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 1.48e-19
C1554 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0231f
C1555 CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 0.0445f
C1556 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 3.88e-20
C1557 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 a_32009_n18723# 2.79e-20
C1558 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_55179_7683# 0.00261f
C1559 CLK a_33204_6159# 4.6e-20
C1560 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_34308_n17626# 8.64e-19
C1561 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 1.49e-21
C1562 F2 F1 2.87f
C1563 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_29623_6159# 4.52e-20
C1564 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00243f
C1565 VDD100 a_53008_n2243# 0.00727f
C1566 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.313f
C1567 a_26984_10099# a_27144_10099# 0.0504f
C1568 CLK a_51487_n10161# 0.00164f
C1569 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.321f
C1570 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB a_47341_1671# 2.96e-19
C1571 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 0.647f
C1572 a_48258_n10160# m3_20882_n11188# 0.00102f
C1573 RST CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 0.288f
C1574 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 3.55e-20
C1575 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 0.0108f
C1576 VDD108 F1 0.00936f
C1577 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.0147f
C1578 VDD100 a_39420_6821# 6.05e-19
C1579 RST CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.166f
C1580 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN 0.112f
C1581 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT 2.59e-20
C1582 a_26266_11196# a_26426_11196# 0.0504f
C1583 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 1.17f
C1584 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 a_27180_n15491# 0.069f
C1585 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_53375_1671# 0.0059f
C1586 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 a_28267_n7033# 0.00353f
C1587 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C1588 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C1589 VDD110 a_48712_n17599# 0.00152f
C1590 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_51598_9057# 9.32e-19
C1591 CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN a_30760_n20290# 0.132f
C1592 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_22620_n9884# 0.0733f
C1593 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT a_37436_n1822# 9.43e-19
C1594 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT 0.103f
C1595 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 0.027f
C1596 VDD90 a_33358_5062# 3.14e-19
C1597 CLK_div_108_new_mag_0.CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 6.02e-20
C1598 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_53333_10154# 0.00378f
C1599 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_45541_n18696# 2.96e-19
C1600 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00301f
C1601 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0894f
C1602 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00118f
C1603 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.00481f
C1604 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_25482_n16632# 1.5e-20
C1605 VDD93 a_36042_6821# 0.00218f
C1606 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB a_47751_2768# 0.00696f
C1607 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN 0.146f
C1608 RST CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0914f
C1609 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_0.OUT a_26250_1919# 0.00378f
C1610 a_52923_9057# CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 8.17e-21
C1611 VDD96 a_29110_n743# 2.21e-19
C1612 a_47914_n16726# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 1.04e-19
C1613 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 0.00212f
C1614 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 1.83e-19
C1615 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 1.96e-19
C1616 VDD110 a_44971_n17599# 0.00123f
C1617 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 9.24e-20
C1618 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 m3_20882_n11188# 0.041f
C1619 RST a_25055_n7107# 0.00173f
C1620 CLK_div_105_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_55179_7683# 5.39e-20
C1621 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 7.86e-19
C1622 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN 0.512f
C1623 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_51239_n5724# 0.069f
C1624 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_35460_n15495# 3.33e-19
C1625 CLK a_43895_n16724# 0.00224f
C1626 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 a_53785_2768# 0.0101f
C1627 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 0.339f
C1628 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_48986_n2199# 0.0811f
C1629 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_35026_n18723# 0.00119f
C1630 CLK_div_108_new_mag_0.JK_FF_mag_1.Q a_49945_n6865# 0.00335f
C1631 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_23743_5062# 0.069f
C1632 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_33180_n17626# 2.58e-20
C1633 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB a_28734_n9876# 0.00696f
C1634 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB a_49794_1671# 0.0114f
C1635 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 2.34e-19
C1636 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00118f
C1637 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 1.01e-19
C1638 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB 0.308f
C1639 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 8.16e-20
C1640 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.122f
C1641 VDD93 a_29298_n9832# 3.14e-19
C1642 CLK_div_90_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 4.39e-19
C1643 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 8.51e-22
C1644 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 a_50263_5143# 0.00789f
C1645 CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.338f
C1646 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 0.00165f
C1647 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.266f
C1648 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.0014f
C1649 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00162f
C1650 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_35192_n17626# 0.0202f
C1651 CLK CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 0.0114f
C1652 RST CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.0123f
C1653 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 0.554f
C1654 CLK CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 1.48e-20
C1655 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_28490_11196# 0.00372f
C1656 VDD99 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 0.00933f
C1657 VDD90 a_32795_11196# 0.0012f
C1658 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 a_29801_1733# 6.83e-19
C1659 CLK_div_90_mag_0.CLK_div_10_mag_0.CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 1.48e-20
C1660 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 1.32e-19
C1661 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 8.04e-19
C1662 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00264f
C1663 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT a_26820_3016# 1.5e-20
C1664 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB 0.11f
C1665 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_47994_n18696# 3.25e-19
C1666 VDD93 a_36109_n8931# 2.65e-19
C1667 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 2.84e-19
C1668 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 1.05e-20
C1669 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 a_44888_1671# 6.43e-21
C1670 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB 0.911f
C1671 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 3.48e-19
C1672 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0306f
C1673 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN 5.57e-20
C1674 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 7.24e-19
C1675 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 1.07f
C1676 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K 6.19e-22
C1677 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_26420_10099# 0.0202f
C1678 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 a_44357_n10160# 0.0101f
C1679 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C1680 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_26606_6159# 4.52e-20
C1681 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 a_45570_10154# 0.00789f
C1682 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.0463f
C1683 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.00183f
C1684 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 3.38e-19
C1685 VDD96 a_25484_n2996# 0.00108f
C1686 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 1.5e-20
C1687 VDD105 a_53850_6284# 3.14e-19
C1688 RST CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 0.00222f
C1689 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 6.11e-19
C1690 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_27227_398# 0.0112f
C1691 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00101f
C1692 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_27144_10099# 8.64e-19
C1693 a_46980_n1146# a_47140_n1146# 0.0504f
C1694 VDD105 a_54568_5187# 3.14e-19
C1695 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 a_45000_9057# 6.43e-21
C1696 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN 6.85e-19
C1697 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 0.0376f
C1698 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 a_28580_n8735# 1.43e-19
C1699 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_54383_n5721# 0.0059f
C1700 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 9.75e-21
C1701 a_39124_880# Vdiv108 7.52e-19
C1702 VDD110 a_43895_n16724# 2.21e-19
C1703 RST a_23794_n17626# 7.28e-19
C1704 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 0.203f
C1705 dec3x8_ibr_mag_0.and_3_ibr_1.nand3_mag_ibr_0.OUT a_37328_6821# 0.0779f
C1706 a_23510_n15620# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 0.132f
C1707 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB a_32795_11196# 0.00695f
C1708 a_46974_n2243# a_47134_n2243# 0.0504f
C1709 VDD CLK 0.547f
C1710 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_53255_n5765# 0.0732f
C1711 RST a_26817_n699# 8.5e-19
C1712 CLK a_43719_n120# 6.43e-19
C1713 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_46964_n9019# 0.069f
C1714 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.514f
C1715 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT 1.2e-19
C1716 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00183f
C1717 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.159f
C1718 VDD93 a_30164_n7017# 3.14e-19
C1719 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.469f
C1720 a_52811_1671# CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 8.17e-21
C1721 a_29298_n9832# m3_20882_n11188# 2.84e-19
C1722 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.122f
C1723 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K F2 0.00315f
C1724 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT 2.67e-20
C1725 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_24116_n1789# 0.00372f
C1726 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 1.53e-20
C1727 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT 0.00157f
C1728 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 8.64e-20
C1729 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 m3_20882_n11188# 0.00101f
C1730 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_31512_6115# 0.00119f
C1731 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_52139_n18696# 0.0114f
C1732 VDD105 a_54057_10154# 0.00123f
C1733 Vdiv108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB 5.82e-21
C1734 RST a_53280_5143# 0.00186f
C1735 VDD96 a_28828_1497# 5.92e-19
C1736 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 3.47f
C1737 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_33812_n13270# 1.9e-19
C1738 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C1739 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1.77e-19
C1740 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 1.37e-20
C1741 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_43993_n13477# 0.015f
C1742 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00335f
C1743 CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN a_50232_n7685# 0.132f
C1744 VDD99 a_24358_n17626# 3.14e-19
C1745 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 3.28e-21
C1746 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 1.86e-19
C1747 CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 2f
C1748 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0052f
C1749 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_44321_n6273# 0.0202f
C1750 a_46774_n6273# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0732f
C1751 RST CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.109f
C1752 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_29208_10099# 4.52e-20
C1753 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.321f
C1754 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0894f
C1755 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.911f
C1756 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_43957_n2243# 1.17e-20
C1757 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 a_48252_n9063# 3.51e-19
C1758 CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_90_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 3.34e-19
C1759 CLK_div_100_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 4.39e-19
C1760 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.161f
C1761 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB 1.99f
C1762 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.076f
C1763 CLK a_26974_1919# 0.0101f
C1764 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.00739f
C1765 RST CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.194f
C1766 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 0.0506f
C1767 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_24938_n9875# 1.5e-20
C1768 RST a_52769_10154# 9.66e-19
C1769 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT 8.51e-22
C1770 RST a_52811_1671# 6.14e-19
C1771 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 a_31346_5018# 0.00117f
C1772 CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 a_53120_5143# 0.00335f
C1773 RST a_22275_10099# 5.16e-19
C1774 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 0.119f
C1775 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00183f
C1776 CLK_div_96_mag_0.JK_FF_mag_4.Q a_24968_3016# 0.0157f
C1777 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00335f
C1778 CLK a_51393_n6821# 3.54e-21
C1779 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT a_23869_810# 1.17e-20
C1780 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 8.16e-20
C1781 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.0126f
C1782 RST a_23249_11196# 0.00221f
C1783 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 9.8e-20
C1784 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_32015_n17626# 1.46e-19
C1785 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_48098_n10160# 1.46e-19
C1786 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00393f
C1787 VDD VDD110 0.404f
C1788 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0592f
C1789 VDD105 a_39580_6821# 7.36e-19
C1790 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.0151f
C1791 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.745f
C1792 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 3.67e-20
C1793 F2 a_39420_6821# 0.00692f
C1794 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 a_24938_n9875# 0.00216f
C1795 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.514f
C1796 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_54621_10154# 0.0731f
C1797 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT a_35747_n1822# 0.00949f
C1798 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.0263f
C1799 CLK a_23025_6159# 2.18e-20
C1800 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 6.28e-19
C1801 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 1.48e-20
C1802 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 a_33204_6159# 0.069f
C1803 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 4.92e-19
C1804 RST a_22982_n2930# 0.00106f
C1805 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.122f
C1806 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 0.179f
C1807 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 1.73e-20
C1808 CLK_div_99_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_25364_n19822# 0.069f
C1809 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.235f
C1810 F1 dec3x8_ibr_mag_0.and_3_ibr_5.nand3_mag_ibr_0.OUT 0.259f
C1811 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.27f
C1812 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_54592_n18696# 2.96e-19
C1813 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 Vdiv110 0.00436f
C1814 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 a_50358_1671# 6.06e-21
C1815 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_45570_10154# 1.46e-19
C1816 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_50875_n2243# 0.00696f
C1817 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 0.198f
C1818 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT 0.266f
C1819 RST CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.152f
C1820 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C1821 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C1822 Vdiv110 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 5.47e-19
C1823 RST a_50304_n16724# 0.00257f
C1824 VDD100 a_53375_1671# 3.14e-19
C1825 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB 0.00258f
C1826 RST a_51439_n2199# 9.41e-19
C1827 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0969f
C1828 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 a_44324_1671# 0.069f
C1829 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 a_23948_n13382# 0.00718f
C1830 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.VOUT 0.122f
C1831 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_33204_6159# 0.00372f
C1832 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT a_47030_n16726# 0.0202f
C1833 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 a_50880_10154# 8.64e-19
C1834 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN 0.112f
C1835 VDD90 VDD99 0.045f
C1836 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00118f
C1837 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.765f
C1838 RST a_47424_n17599# 0.00247f
C1839 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 0.0044f
C1840 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_32070_5018# 0.0203f
C1841 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 4.44e-20
C1842 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB 0.141f
C1843 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 0.0112f
C1844 CLK CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.0215f
C1845 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK 2.53e-19
C1846 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 a_43947_n9019# 0.069f
C1847 CLK a_44407_n17599# 4.62e-19
C1848 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C1849 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_2.OUT CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 0.00118f
C1850 CLK_div_96_mag_0.JK_FF_mag_5.Q CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_4.IN2 0.0635f
C1851 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT 0.768f
C1852 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 a_39124_280# 0.00372f
C1853 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.00388f
C1854 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 a_30317_n18723# 0.00372f
C1855 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.038f
C1856 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K 0.0156f
C1857 CLK a_44075_6240# 0.0101f
C1858 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT a_50903_n5# 7.43e-22
C1859 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.272f
C1860 RST a_34890_n16636# 0.00201f
C1861 RST a_23594_n8743# 0.00221f
C1862 CLK a_46081_5187# 5.03e-19
C1863 CLK_div_90_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_22718_8532# 3.25e-19
C1864 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00152f
C1865 Vdiv90 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 0.00411f
C1866 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT a_43895_n16724# 0.0202f
C1867 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_44841_n2243# 8.64e-19
C1868 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00306f
C1869 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 2.86f
C1870 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 Vdiv110 0.00131f
C1871 VDD96 a_29307_n1855# 3.14e-19
C1872 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 5.57e-19
C1873 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00183f
C1874 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_55019_7683# 0.00239f
C1875 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.108f
C1876 VDD105 F1 0.0132f
C1877 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.419f
C1878 CLK a_32640_6159# 4.6e-20
C1879 VDD100 a_52003_n2199# 0.00152f
C1880 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_29059_6159# 0.0202f
C1881 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT a_44625_n15583# 0.00378f
C1882 F1 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT 4.77e-19
C1883 CLK CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00131f
C1884 VDD99 a_38454_6821# 0.00126f
C1885 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB a_46777_1671# 0.0114f
C1886 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 CLK_div_96_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.305f
C1887 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 2.01e-19
C1888 a_48098_n10160# m3_20882_n11188# 0.00102f
C1889 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT 1.48e-19
C1890 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 1.34e-19
C1891 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 0.741f
C1892 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 9.98e-19
C1893 RST CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 0.134f
C1894 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00158f
C1895 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C1896 CLK_div_108_new_mag_0.JK_FF_mag_1.Q CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 1.4e-20
C1897 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 0.492f
C1898 VDD99 a_35454_n16636# 2.21e-19
C1899 mux_8x1_ibr_0.mux_2x1_ibr_0.I0 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 3.43e-19
C1900 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0957f
C1901 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_51034_9057# 3.12e-19
C1902 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT a_36873_n1822# 0.00949f
C1903 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_22460_n9884# 0.0203f
C1904 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 9.9e-19
C1905 a_24512_n18723# CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 4.9e-20
C1906 CLK_div_100_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 CLK_div_100_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.11f
C1907 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.215f
C1908 Vdiv110 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 0.374f
C1909 VDD90 a_32794_5062# 3.14e-19
C1910 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT 7.24e-19
C1911 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_44977_n18696# 3.33e-19
C1912 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 0.104f
C1913 Vdiv90 dec3x8_ibr_mag_0.and_3_ibr_5.IN3 2.68e-19
C1914 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 2.61e-19
C1915 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_25322_n16632# 1.17e-20
C1916 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C1917 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 4.76e-19
C1918 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB a_47187_2768# 0.00964f
C1919 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 7.84e-19
C1920 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 0.235f
C1921 VDD96 a_28546_n743# 3.1e-20
C1922 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00718f
C1923 RST CLK_div_108_new_mag_0.CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 0.00746f
C1924 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 0.00396f
C1925 CLK CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT 0.235f
C1926 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0759f
C1927 VDD96 a_23145_810# 2.21e-19
C1928 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_23025_6159# 0.00378f
C1929 VDD110 a_44407_n17599# 0.00892f
C1930 VDD96 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 7.04e-22
C1931 RST CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT 0.284f
C1932 RST a_24491_n7107# 0.00252f
C1933 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT a_51764_10154# 0.0202f
C1934 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0573f
C1935 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_48466_n6273# 0.00118f
C1936 CLK_div_105_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_55019_7683# 9.16e-20
C1937 CLK_div_96_mag_0.JK_FF_mag_0.QB CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.343f
C1938 VDD96 CLK_div_96_mag_0.JK_FF_mag_4.Q 2.21f
C1939 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.36f
C1940 VDD93 a_26636_n8734# 3.56e-19
C1941 a_33405_7558# Vdiv90 0.198f
C1942 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_34896_n15539# 0.00392f
C1943 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 8.59e-20
C1944 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 a_30589_n2952# 0.00372f
C1945 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 a_53221_2768# 0.00859f
C1946 a_44734_2768# a_44894_2768# 0.0504f
C1947 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_48252_n9063# 8.64e-19
C1948 dec3x8_ibr_mag_0.and_3_ibr_0.nand3_mag_ibr_0.OUT dec3x8_ibr_mag_0.and_3_ibr_1.nand3_mag_ibr_0.OUT 6.9e-19
C1949 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT 0.00123f
C1950 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.122f
C1951 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_48422_n2199# 0.00964f
C1952 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN a_52951_7381# 5.1e-20
C1953 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_34462_n18723# 1.43e-19
C1954 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB 0.28f
C1955 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.802f
C1956 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.359f
C1957 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT a_52225_n13362# 8.09e-22
C1958 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 1.18e-19
C1959 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0622f
C1960 Vdiv110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.00185f
C1961 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB a_28574_n9876# 0.00695f
C1962 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.21f
C1963 RST CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.0498f
C1964 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT 4.36e-19
C1965 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 3.04f
C1966 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 m3_20882_n11188# 3.33e-19
C1967 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.28f
C1968 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 a_50103_5143# 0.00335f
C1969 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.746f
C1970 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 a_37999_n1822# 0.00372f
C1971 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_35032_n17626# 0.0731f
C1972 VDD96 CLK_div_96_mag_0.JK_FF_mag_5.Q 2.19f
C1973 VDD90 a_32635_11196# 9.82e-19
C1974 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 a_48587_10154# 1.46e-19
C1975 RST CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.161f
C1976 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT a_26256_3016# 0.0203f
C1977 VDD93 a_35949_n8931# 6.05e-19
C1978 VDD93 RST 7f
C1979 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K Vdiv 1.75e-19
C1980 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 a_25532_3016# 0.069f
C1981 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_25800_n18723# 0.0203f
C1982 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 8.33e-20
C1983 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_37391_n9984# 0.0036f
C1984 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 a_43757_n6273# 2.79e-20
C1985 CLK_div_99_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN a_30760_n20290# 3.25e-19
C1986 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 m3_20882_n11188# 3.21e-19
C1987 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 a_43793_n10116# 0.00859f
C1988 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 a_37999_n1822# 2.44e-19
C1989 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_25856_10099# 4.52e-20
C1990 a_30398_n699# CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 4.58e-20
C1991 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 0.103f
C1992 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_26042_6159# 0.0202f
C1993 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 a_45006_10154# 0.0102f
C1994 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB a_54057_10154# 0.00695f
C1995 VDD99 dec3x8_ibr_mag_0.and_3_ibr_7.nand3_mag_ibr_0.OUT 6.02e-19
C1996 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_44977_n18696# 0.00378f
C1997 VDD96 a_24270_n2886# 3.54e-19
C1998 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 a_26206_n16632# 8.64e-19
C1999 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 0.12f
C2000 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_24307_5062# 0.0811f
C2001 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C2002 VDD100 dec3x8_ibr_mag_0.and_3_ibr_7.nand3_mag_ibr_0.OUT 8.19e-20
C2003 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 1f
C2004 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 0.0314f
C2005 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 a_28016_n8779# 0.00119f
C2006 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.273f
C2007 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.0661f
C2008 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 0.0113f
C2009 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 0.321f
C2010 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_53819_n5721# 0.0697f
C2011 a_38561_880# Vdiv108 5.59e-19
C2012 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 8.2e-19
C2013 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.31f
C2014 CLK_div_96_mag_0.JK_FF_mag_2.Q CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.0635f
C2015 dec3x8_ibr_mag_0.and_3_ibr_2.nand3_mag_ibr_0.OUT dec3x8_ibr_mag_0.and_3_ibr_3.nand3_mag_ibr_0.OUT 6.97e-19
C2016 dec3x8_ibr_mag_0.and_3_ibr_1.nand3_mag_ibr_0.OUT a_37168_6821# 0.0249f
C2017 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB a_32635_11196# 0.00696f
C2018 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 3.14f
C2019 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_53095_n5765# 0.0203f
C2020 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 8.16e-20
C2021 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 2.61e-19
C2022 CLK a_43559_n120# 0.00136f
C2023 RST a_26253_n743# 0.00147f
C2024 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.122f
C2025 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_46400_n9019# 0.00372f
C2026 CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 8.98e-19
C2027 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 3.8e-20
C2028 a_28734_n9876# m3_20882_n11188# 2.89e-19
C2029 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 m3_20882_n11188# 0.0195f
C2030 dec3x8_ibr_mag_0.and_3_ibr_5.IN3 dec3x8_ibr_mag_0.and_3_ibr_4.nand3_mag_ibr_0.OUT 0.289f
C2031 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 2.11e-19
C2032 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.28f
C2033 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_23552_n1789# 0.069f
C2034 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K a_45724_9057# 8.64e-19
C2035 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.313f
C2036 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_51575_n18696# 2.96e-19
C2037 VDD105 a_53897_10154# 0.00101f
C2038 RST a_53120_5143# 0.00186f
C2039 mux_8x1_ibr_0.mux_2x1_ibr_0.I1 Vdiv100 9.62e-20
C2040 CLK_div_96_mag_0.JK_FF_mag_3.QB CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.0387f
C2041 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 0.0343f
C2042 CLK CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K 2.2f
C2043 a_25318_6115# a_25478_6115# 0.0504f
C2044 VDD99 a_23794_n17626# 3.14e-19
C2045 RST m3_20882_n11188# 1.81f
C2046 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.0635f
C2047 VDD99 a_28463_n15537# 2.21e-19
C2048 RST CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.00289f
C2049 a_50441_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 1.46e-19
C2050 VDD90 F2 0.204f
C2051 F1 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.367f
C2052 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_29772_10099# 0.0697f
C2053 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 8.65e-20
C2054 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT a_31177_7256# 0.00138f
C2055 a_46614_n6273# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0203f
C2056 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.348f
C2057 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 0.36f
C2058 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 8.16e-20
C2059 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 0.109f
C2060 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.397f
C2061 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.305f
C2062 CLK a_26814_1919# 0.00939f
C2063 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 8.04e-19
C2064 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_24778_n9875# 1.17e-20
C2065 a_31731_n16632# CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 5.98e-19
C2066 CLK a_54658_n9064# 0.0101f
C2067 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 a_50470_9057# 0.069f
C2068 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN 0.00323f
C2069 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT a_23709_810# 1.5e-20
C2070 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT a_54033_n15587# 0.00378f
C2071 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 0.109f
C2072 RST a_22685_11196# 0.00123f
C2073 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 0.0979f
C2074 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT 8.51e-22
C2075 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 2.34e-19
C2076 VDD96 F1 0.0836f
C2077 VDD105 a_39420_6821# 0.00124f
C2078 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 a_29708_n8735# 0.00372f
C2079 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_0.OUT a_23863_n287# 0.0203f
C2080 F2 a_38454_6821# 0.0115f
C2081 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 a_24778_n9875# 0.00185f
C2082 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_54057_10154# 9.1e-19
C2083 CLK a_22461_6115# 1.32e-19
C2084 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 2.86f
C2085 RST a_22418_n2930# 4.58e-19
C2086 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.00243f
C2087 F1 a_37328_6265# 0.0102f
C2088 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 2.27e-20
C2089 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 a_49794_1671# 0.069f
C2090 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_54028_n18696# 3.25e-19
C2091 a_45618_2768# Vdiv110 0.00138f
C2092 F1 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I1 0.0593f
C2093 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.655f
C2094 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT Vdiv99 0.00214f
C2095 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_50715_n2243# 0.00695f
C2096 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.00335f
C2097 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.00586f
C2098 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 3.38e-19
C2099 Vdiv110 a_37999_280# 2.66e-19
C2100 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 m3_20882_n11188# 8.77e-19
C2101 RST a_50144_n16724# 0.00257f
C2102 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00152f
C2103 VDD100 a_52811_1671# 3.56e-19
C2104 RST a_50875_n2243# 0.00186f
C2105 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK 0.253f
C2106 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 a_43760_1671# 0.00372f
C2107 RST a_47264_n17599# 0.00247f
C2108 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_32640_6159# 0.069f
C2109 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 0.98f
C2110 CLK CLK_div_105_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 2.42e-19
C2111 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0854f
C2112 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.0215f
C2113 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00154f
C2114 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_31506_5018# 1.5e-20
C2115 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT a_35747_280# 0.0964f
C2116 CLK a_32169_n18723# 0.0101f
C2117 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.00153f
C2118 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 1.82e-19
C2119 a_45753_n15583# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 4.52e-20
C2120 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 0.0725f
C2121 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 a_43383_n9019# 0.00372f
C2122 CLK a_44247_n17599# 4.62e-19
C2123 CLK CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 2.59e-19
C2124 a_42521_n13474# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 2.69e-22
C2125 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 1.36e-19
C2126 a_47810_5143# a_47970_5143# 0.0504f
C2127 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.122f
C2128 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 9.41e-19
C2129 RST a_34730_n16636# 0.00201f
C2130 RST a_23030_n8743# 0.00165f
C2131 CLK a_45517_5187# 4.86e-19
C2132 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_45449_n6273# 0.00118f
C2133 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 2.52f
C2134 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_30336_10099# 0.00392f
C2135 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 0.235f
C2136 VDD99 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 1.08e-20
C2137 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.653f
C2138 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 2.44e-20
C2139 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.0881f
C2140 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 6.22e-20
C2141 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN a_48023_n7840# 0.132f
C2142 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN 0.424f
C2143 a_53129_n19793# CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.069f
C2144 CLK_div_96_mag_0.JK_FF_mag_0.Q CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.338f
C2145 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_25662_n9875# 8.64e-19
C2146 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT a_44061_n15627# 0.0732f
C2147 VDD100 a_51439_n2199# 0.00152f
C2148 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.04e-19
C2149 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.321f
C2150 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB 0.904f
C2151 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK CLK_div_108_new_mag_0.CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 1.73e-19
C2152 VDD99 a_38294_6821# 0.0016f
C2153 CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 a_55179_7683# 0.019f
C2154 a_47534_n10160# m3_20882_n11188# 4.29e-19
C2155 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 1.89e-20
C2156 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 a_39580_6821# 0.00244f
C2157 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_27342_n1855# 1.71e-20
C2158 a_36202_6265# dec3x8_ibr_mag_0.and_3_ibr_4.nand3_mag_ibr_0.OUT 0.0779f
C2159 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 4.69e-20
C2160 VDD90 a_30496_10099# 2.21e-19
C2161 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 a_24901_n6010# 0.069f
C2162 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.233f
C2163 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C2164 VDD108 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.3f
C2165 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_41124_n16098# 0.00347f
C2166 VDD99 a_34890_n16636# 7.37e-19
C2167 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 2.81e-20
C2168 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.22f
C2169 CLK_div_96_mag_0.JK_FF_mag_0.Q CLK_div_96_mag_0.JK_FF_mag_2.QB 0.307f
C2170 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_50470_9057# 7.4e-19
C2171 F1 mux_8x1_ibr_0.mux_2x1_ibr_0.I0 0.0118f
C2172 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN 0.514f
C2173 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 8.16e-20
C2174 CLK CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 1.29e-19
C2175 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_21896_n9884# 1.5e-20
C2176 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.00518f
C2177 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.199f
C2178 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.25f
C2179 CLK_div_99_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_24391_n20290# 3.25e-19
C2180 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.0864f
C2181 RST CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 0.0893f
C2182 RST CLK_div_108_new_mag_0.JK_FF_mag_1.Q 0.178f
C2183 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN 2.63e-20
C2184 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.768f
C2185 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB a_46623_2768# 0.0811f
C2186 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT 1.61e-19
C2187 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0951f
C2188 VDD96 a_28386_n743# 0.00743f
C2189 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.235f
C2190 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.122f
C2191 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C2192 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 0.027f
C2193 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_30315_n15493# 0.0114f
C2194 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.748f
C2195 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_45081_n10160# 1.46e-19
C2196 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 0.144f
C2197 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_22461_6115# 0.0732f
C2198 VDD110 a_44247_n17599# 0.0132f
C2199 RST CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0134f
C2200 VDD99 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 1.08e-20
C2201 F2 dec3x8_ibr_mag_0.and_3_ibr_7.nand3_mag_ibr_0.OUT 0.108f
C2202 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K 5.7e-19
C2203 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT a_51604_10154# 0.0731f
C2204 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_47902_n6273# 0.011f
C2205 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_100_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00154f
C2206 VDD93 a_26072_n8734# 3.14e-19
C2207 a_33245_7558# Vdiv90 0.0132f
C2208 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 3.08e-19
C2209 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN a_51871_n5# 0.069f
C2210 VDD108 dec3x8_ibr_mag_0.and_3_ibr_7.nand3_mag_ibr_0.OUT 3.42e-19
C2211 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB a_30496_10099# 1.86e-20
C2212 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 a_30025_n2952# 0.069f
C2213 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 a_52657_2768# 0.0157f
C2214 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_47858_n2243# 0.00696f
C2215 CLK a_44117_n2243# 0.00164f
C2216 CLK CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 0.471f
C2217 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.1f
C2218 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT a_49488_n13383# 2.05e-19
C2219 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 dec3x8_ibr_mag_0.and_3_ibr_2.nand3_mag_ibr_0.OUT 0.127f
C2220 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_33898_n18723# 0.011f
C2221 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 1.36e-19
C2222 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB 0.198f
C2223 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 a_50199_n10117# 0.069f
C2224 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 0.0112f
C2225 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 F1 0.427f
C2226 VDD93 a_28574_n9876# 2.21e-19
C2227 VDD96 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 0.00128f
C2228 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0378f
C2229 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 2.57e-19
C2230 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 a_37436_n1822# 0.069f
C2231 VDD99 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT 0.0122f
C2232 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.00729f
C2233 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_34468_n17626# 9.1e-19
C2234 a_50281_n17599# a_50441_n17599# 0.0504f
C2235 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN 0.303f
C2236 VDD90 a_32071_11196# 0.00149f
C2237 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 0.768f
C2238 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN m3_20882_n11188# 0.0064f
C2239 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 0.00121f
C2240 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT a_26096_3016# 0.0733f
C2241 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 6.22e-20
C2242 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_25662_n9875# 2.88e-20
C2243 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT 0.00395f
C2244 CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 9.34e-19
C2245 RST a_29116_398# 3.41e-19
C2246 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 a_24968_3016# 0.00372f
C2247 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 a_45452_1671# 2.79e-20
C2248 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_25640_n18723# 0.0732f
C2249 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT a_32301_n15491# 0.00378f
C2250 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00229f
C2251 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 0.00376f
C2252 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.105f
C2253 VDD96 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.0224f
C2254 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 a_37436_n1822# 1.04e-19
C2255 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 a_43229_n10116# 0.0157f
C2256 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB a_53897_10154# 0.00696f
C2257 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 a_44846_10154# 0.0101f
C2258 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 0.00542f
C2259 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 9.64e-19
C2260 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 6.02e-20
C2261 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT a_47723_574# 3.38e-20
C2262 VDD96 a_23706_n2886# 3.14e-19
C2263 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 0.741f
C2264 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00156f
C2265 VDD105 a_53126_6240# 2.21e-19
C2266 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.0615f
C2267 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_26099_398# 3.33e-19
C2268 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 1.89e-19
C2269 VDD105 a_53844_5143# 2.21e-19
C2270 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.122f
C2271 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_23743_5062# 0.00964f
C2272 VDD100 a_39580_6265# 7.22e-20
C2273 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 a_45564_9057# 2.79e-20
C2274 CLK_div_96_mag_0.JK_FF_mag_4.QB CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 1.32e-19
C2275 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 1.49e-21
C2276 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT a_37999_280# 0.0964f
C2277 a_44619_n16724# a_44779_n16724# 0.0504f
C2278 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 2.61e-19
C2279 a_37999_880# Vdiv108 7.52e-19
C2280 VDD93 VDD99 0.302f
C2281 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.109f
C2282 a_47902_n6273# CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 4.9e-20
C2283 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB a_32071_11196# 0.00964f
C2284 RST a_26093_n743# 8.64e-19
C2285 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0626f
C2286 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.21f
C2287 CLK_div_100_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 a_55067_297# 2.44e-20
C2288 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 9.24e-20
C2289 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_44517_n10160# 0.00695f
C2290 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN a_31177_7256# 0.069f
C2291 a_28574_n9876# m3_20882_n11188# 2.89e-19
C2292 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.00481f
C2293 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 3.43e-19
C2294 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.0592f
C2295 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00233f
C2296 dec3x8_ibr_mag_0.and_3_ibr_5.IN3 a_36202_6265# 0.0104f
C2297 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 2.4e-19
C2298 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 a_54781_10154# 0.00335f
C2299 VDD99 F0 0.104f
C2300 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 0.36f
C2301 Vdiv105 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 1.08e-19
C2302 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 1.53e-20
C2303 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.IN1 0.091f
C2304 VDD100 F0 0.0749f
C2305 RST a_50833_6284# 1.23e-20
C2306 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_51011_n18696# 3.25e-19
C2307 VDD105 a_53333_10154# 0.00152f
C2308 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.103f
C2309 RST a_52115_5187# 9.66e-19
C2310 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0622f
C2311 a_29618_11196# a_29778_11196# 0.0504f
C2312 RST CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0299f
C2313 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 0.198f
C2314 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.122f
C2315 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 9.52e-19
C2316 VDD99 a_27180_n15491# 3.56e-19
C2317 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 0.0165f
C2318 RST a_28817_n18723# 6.26e-19
C2319 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT 1.29e-19
C2320 VDD90 a_31177_7256# 3.14e-19
C2321 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_29208_10099# 0.0059f
C2322 a_46614_n6273# a_46774_n6273# 0.0504f
C2323 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.122f
C2324 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 5.45e-20
C2325 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 5.42e-20
C2326 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 1.7e-20
C2327 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 0.285f
C2328 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 0.01f
C2329 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 2.54e-20
C2330 CLK a_26250_1919# 6.43e-21
C2331 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0622f
C2332 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00158f
C2333 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.00586f
C2334 a_36588_n15495# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 4.52e-20
C2335 a_31571_n16632# CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 5.98e-19
C2336 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_26984_10099# 0.00392f
C2337 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 a_49906_9057# 0.00372f
C2338 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB Vdiv110 0.0101f
C2339 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.00183f
C2340 CLK a_54498_n9064# 0.00939f
C2341 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT a_35747_n1222# 0.0964f
C2342 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 1.9e-19
C2343 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT a_23145_810# 0.0203f
C2344 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT a_53469_n15631# 0.0732f
C2345 VDD99 m3_20882_n11188# 0.938f
C2346 RST a_22121_11196# 0.00114f
C2347 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.398f
C2348 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 3.31e-20
C2349 VDD mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 0.456f
C2350 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_4.IN2 a_22421_810# 0.069f
C2351 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT 6.64e-19
C2352 VDD105 a_38454_6821# 0.00174f
C2353 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.0205f
C2354 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 a_29144_n8735# 0.069f
C2355 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 8.94e-19
C2356 F2 a_38294_6821# 0.00241f
C2357 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_0.OUT a_23703_n287# 0.0732f
C2358 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 a_23748_n9840# 0.0157f
C2359 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_27342_n1855# 0.00118f
C2360 CLK a_22301_6115# 1.63e-19
C2361 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_53897_10154# 2.88e-20
C2362 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_52839_n5# 8.17e-21
C2363 RST a_22258_n2930# 4.58e-19
C2364 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C2365 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 0.0979f
C2366 F1 a_37168_6265# 0.00731f
C2367 a_26036_5018# a_26196_5018# 0.0504f
C2368 a_45458_2768# Vdiv110 0.00138f
C2369 a_48888_n15585# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 4.52e-20
C2370 a_49951_n5768# a_50111_n5768# 0.0504f
C2371 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.109f
C2372 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_47970_5143# 2.88e-20
C2373 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 0.139f
C2374 RST a_47760_n15585# 3.08e-20
C2375 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0622f
C2376 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN 8.53e-19
C2377 VDD96 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 0.391f
C2378 CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 CLK_div_100_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00357f
C2379 RST a_49042_n16682# 0.00129f
C2380 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 2.35e-19
C2381 Vdiv105 Vdiv 0.906f
C2382 RST a_50715_n2243# 0.00169f
C2383 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_45564_9057# 0.00119f
C2384 CLK_div_100_mag_0.CLK_div_10_mag_1.CLK Vdiv110 0.0222f
C2385 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.235f
C2386 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_31346_5018# 1.17e-20
C2387 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 3.06f
C2388 CLK_div_96_mag_0.JK_FF_mag_5.Q CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT 0.0345f
C2389 CLK a_32009_n18723# 0.00939f
C2390 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 2.04e-19
C2391 CLK a_35192_n17626# 0.00117f
C2392 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 0.0177f
C2393 RST CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.0545f
C2394 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 2.6e-20
C2395 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 8.58e-20
C2396 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 0.391f
C2397 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN a_43831_7266# 2.85e-20
C2398 Vdiv99 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 8.44e-19
C2399 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.00602f
C2400 RST a_22466_n8743# 3.21e-19
C2401 a_38960_n10028# a_39120_n10028# 0.0504f
C2402 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_44885_n6273# 0.011f
C2403 CLK a_44953_5143# 4.68e-19
C2404 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_29772_10099# 1.75e-19
C2405 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT a_28734_n9876# 2.88e-20
C2406 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 9.62e-20
C2407 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.291f
C2408 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT 0.235f
C2409 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 1.07f
C2410 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 2.58f
C2411 VDD96 a_28583_n1899# 0.00535f
C2412 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.108f
C2413 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.121f
C2414 CLK_div_108_new_mag_0.JK_FF_mag_1.QB CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.28f
C2415 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK CLK_div_108_new_mag_0.JK_FF_mag_1.Q 0.161f
C2416 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0334f
C2417 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 0.209f
C2418 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 a_30317_n18723# 0.069f
C2419 VDD110 a_42529_n14305# 3.85e-19
C2420 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 4.78e-20
C2421 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT a_43901_n15627# 0.0203f
C2422 VDD100 a_50875_n2243# 0.00101f
C2423 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0309f
C2424 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 0.0116f
C2425 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_44841_n2243# 2.88e-20
C2426 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN 0.0042f
C2427 a_47374_n10160# m3_20882_n11188# 4.29e-19
C2428 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT 0.0826f
C2429 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 a_39420_6821# 0.00175f
C2430 CLK Vdiv100 0.249f
C2431 a_36042_6265# dec3x8_ibr_mag_0.and_3_ibr_4.nand3_mag_ibr_0.OUT 0.0249f
C2432 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 a_24337_n6010# 0.00372f
C2433 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.289f
C2434 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_30398_n699# 0.00372f
C2435 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_32175_n17626# 1.17e-20
C2436 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 a_25488_n15535# 3.43e-19
C2437 VDD99 a_34730_n16636# 9.58e-19
C2438 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C2439 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 0.465f
C2440 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_49906_9057# 7.4e-19
C2441 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.00447f
C2442 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 0.00825f
C2443 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 0.98f
C2444 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_21736_n9884# 1.17e-20
C2445 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.802f
C2446 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 1.97f
C2447 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 a_43947_n9019# 4.9e-20
C2448 VDD90 a_32070_5018# 2.21e-19
C2449 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.00335f
C2450 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT a_50721_n1102# 0.00378f
C2451 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_48148_n17599# 8.64e-19
C2452 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_45730_10154# 1.17e-20
C2453 CLK_div_90_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 4.25e-20
C2454 VDD96 a_27381_n699# 0.00149f
C2455 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 1.29e-20
C2456 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 3.28e-19
C2457 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 0.122f
C2458 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 1.53e-19
C2459 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_29751_n15493# 2.96e-19
C2460 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0635f
C2461 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 8.58e-20
C2462 VDD96 a_22421_810# 3.14e-19
C2463 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0228f
C2464 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_22301_6115# 0.0203f
C2465 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.346f
C2466 CLK_div_96_mag_0.JK_FF_mag_0.QB CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.0388f
C2467 VDD105 dec3x8_ibr_mag_0.and_3_ibr_7.nand3_mag_ibr_0.OUT 0.0241f
C2468 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 0.321f
C2469 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 0.434f
C2470 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.00568f
C2471 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT a_51040_10154# 9.1e-19
C2472 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_47338_n6273# 1.43e-19
C2473 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_32230_5018# 8.64e-19
C2474 VDD108 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.756f
C2475 Vdiv110 Vdiv108 1.03f
C2476 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 0.0502f
C2477 VDD93 a_25508_n8734# 3.14e-19
C2478 a_33245_7558# a_33405_7558# 0.186f
C2479 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB a_30336_10099# 1.41e-20
C2480 Vdiv108 a_44687_n1102# 1.08e-19
C2481 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.768f
C2482 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_47698_n2243# 0.00695f
C2483 CLK a_43957_n2243# 0.00117f
C2484 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.833f
C2485 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.101f
C2486 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_47430_n18696# 9.32e-19
C2487 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 1.24f
C2488 VDD93 F2 1.06f
C2489 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 a_30435_n1855# 0.00372f
C2490 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_33334_n18723# 0.00118f
C2491 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT a_48783_n13424# 0.0731f
C2492 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 6.24e-20
C2493 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 3.44e-20
C2494 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 1.01f
C2495 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 a_49635_n10117# 0.00372f
C2496 Vdiv96 a_36873_n1822# 7.87e-19
C2497 RST CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.00511f
C2498 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN Vdiv96 0.131f
C2499 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 0.11f
C2500 Vdiv108 a_39124_280# 0.00237f
C2501 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_45405_n2199# 0.0036f
C2502 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT 1.26e-19
C2503 RST CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 0.045f
C2504 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 4.24e-20
C2505 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT 0.00183f
C2506 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 6.18e-19
C2507 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.08f
C2508 F2 F0 0.465f
C2509 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_0.OUT CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0017f
C2510 a_54947_n5721# CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 4.52e-20
C2511 mux_8x1_ibr_0.mux_2x1_ibr_0.I1 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 0.11f
C2512 VDD110 Vdiv100 0.114f
C2513 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_34308_n17626# 2.88e-20
C2514 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.00123f
C2515 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 4.42e-19
C2516 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_29623_6159# 0.0059f
C2517 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN 0.0012f
C2518 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.122f
C2519 VDD90 a_31507_11196# 0.00149f
C2520 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_48023_n7840# 0.00168f
C2521 VDD108 F0 0.089f
C2522 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 0.0276f
C2523 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 0.231f
C2524 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT a_25532_3016# 0.00378f
C2525 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 1.93f
C2526 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.215f
C2527 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_25502_n9875# 9.1e-19
C2528 RST CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.312f
C2529 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 4.21e-20
C2530 RST a_28552_354# 0.00156f
C2531 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 3.09e-19
C2532 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_25076_n18723# 0.00378f
C2533 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 0.397f
C2534 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.IN1 0.00501f
C2535 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT a_31737_n15535# 0.0732f
C2536 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 8.27e-19
C2537 VDD90 VDD96 0.982f
C2538 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C2539 a_54592_n18696# CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 5.94e-20
C2540 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 a_36873_n1822# 2.44e-19
C2541 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_22620_n9884# 8.64e-19
C2542 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 a_44282_10154# 0.00859f
C2543 CLK_div_108_new_mag_0.CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 6.11e-19
C2544 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB a_53333_10154# 0.00964f
C2545 CLK_div_100_mag_0.CLK_div_10_mag_1.CLK a_54669_2768# 0.00117f
C2546 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 8.26e-20
C2547 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 0.777f
C2548 a_53487_9057# CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 8.17e-21
C2549 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K a_34736_n15539# 0.00472f
C2550 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0129f
C2551 VDD105 a_51961_6284# 3.56e-19
C2552 RST CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.145f
C2553 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_25535_354# 0.00392f
C2554 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN 0.00382f
C2555 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_23179_5018# 0.00696f
C2556 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00137f
C2557 VDD100 a_39420_6265# 9.99e-20
C2558 VDD105 a_53280_5143# 0.00299f
C2559 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.019f
C2560 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 1.45e-19
C2561 a_26046_n16632# a_26206_n16632# 0.0504f
C2562 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.VOUT CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN 1.26e-19
C2563 a_37436_880# Vdiv108 5.59e-19
C2564 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K a_28457_n16634# 8.64e-19
C2565 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 2.96e-19
C2566 a_29301_n2996# a_29461_n2996# 0.0504f
C2567 CLK CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 1.29e-19
C2568 a_53089_n6862# a_53249_n6862# 0.0504f
C2569 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB a_31507_11196# 0.0811f
C2570 CLK_div_90_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 0.00442f
C2571 a_50880_10154# a_51040_10154# 0.0504f
C2572 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 1.29e-19
C2573 CLK_div_100_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 a_54907_297# 9.02e-19
C2574 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_44357_n10160# 0.00696f
C2575 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0201f
C2576 a_28010_n9876# m3_20882_n11188# 6.86e-19
C2577 VDD108 m3_20882_n11188# 0.138f
C2578 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT a_47704_n1102# 0.00378f
C2579 a_48783_n13424# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 4.33e-21
C2580 dec3x8_ibr_mag_0.and_3_ibr_5.IN3 a_36042_6265# 0.00321f
C2581 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 a_54621_10154# 0.00789f
C2582 VDD mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 0.46f
C2583 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.00137f
C2584 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_48324_n15585# 4.52e-20
C2585 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 8.16e-20
C2586 VDD105 a_52769_10154# 0.00152f
C2587 RST a_51551_5187# 9.41e-19
C2588 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 1.77e-19
C2589 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.41f
C2590 CLK_div_90_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 7.14e-19
C2591 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.235f
C2592 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 m3_20882_n11188# 0.032f
C2593 RST CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.014f
C2594 RST a_55357_n20487# 4.79e-19
C2595 VDD99 a_26616_n15491# 3.14e-19
C2596 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 0.0127f
C2597 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.101f
C2598 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.177f
C2599 RST a_28657_n18723# 5.13e-19
C2600 VDD110 dec3x8_ibr_mag_0.and_3_ibr_3.nand3_mag_ibr_0.OUT 0.0338f
C2601 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0728f
C2602 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT a_48747_10154# 1.17e-20
C2603 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0836f
C2604 Vdiv93 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 6.64e-19
C2605 a_49276_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.0811f
C2606 CLK_div_105_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 a_54978_6284# 2.1e-20
C2607 RST CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 0.354f
C2608 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 6.23e-19
C2609 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT 0.999f
C2610 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_24944_n8778# 3.42e-20
C2611 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.VOUT 0.0102f
C2612 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_26420_10099# 3.33e-19
C2613 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT 0.1f
C2614 CLK a_53934_n9020# 6.43e-21
C2615 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C2616 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C2617 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_26606_6159# 0.0059f
C2618 CLK_div_96_mag_0.JK_FF_mag_0.Q CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 6.64e-19
C2619 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT a_22985_810# 0.0733f
C2620 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 a_22551_n16006# 4.44e-20
C2621 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT a_53309_n15631# 0.0203f
C2622 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.00158f
C2623 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.065f
C2624 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_26770_n16588# 0.0036f
C2625 VDD99 a_28817_n18723# 5.99e-19
C2626 RST CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 0.00258f
C2627 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_30727_n17626# 0.0036f
C2628 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.CLK 0.0262f
C2629 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 3.67e-20
C2630 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_4.IN2 a_21857_810# 0.00372f
C2631 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.101f
C2632 VDD100 m1_42708_4265# 0.00929f
C2633 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_46810_n10116# 0.0036f
C2634 RST CLK_div_108_new_mag_0.JK_FF_mag_0.QB 0.107f
C2635 CLK CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 1.22e-19
C2636 VDD105 a_38294_6821# 0.00139f
C2637 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 0.11f
C2638 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 0.648f
C2639 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 0.516f
C2640 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_0.OUT a_23139_n287# 0.00378f
C2641 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 a_23184_n9840# 0.00859f
C2642 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_26778_n1855# 0.011f
C2643 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 a_31512_6115# 2.79e-20
C2644 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 6.13e-20
C2645 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00136f
C2646 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT Vdiv108 0.0404f
C2647 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 a_31129_n6271# 0.00347f
C2648 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 8.98e-19
C2649 a_44894_2768# Vdiv110 5.84e-19
C2650 a_53375_1671# CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 8.17e-21
C2651 a_51871_n5# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 1.29e-22
C2652 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 0.0905f
C2653 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT Vdiv108 0.037f
C2654 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.00975f
C2655 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.231f
C2656 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_44282_10154# 0.0036f
C2657 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_47810_5143# 9.1e-19
C2658 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0343f
C2659 RST a_48478_n16682# 0.00129f
C2660 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN 0.769f
C2661 Vdiv110 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 1.83e-19
C2662 a_45131_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0733f
C2663 RST a_50151_n2243# 0.00186f
C2664 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_45000_9057# 1.43e-19
C2665 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.25f
C2666 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT m3_20882_n11188# 0.00167f
C2667 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 2.15e-20
C2668 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 0.00119f
C2669 VDD90 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 0.0583f
C2670 CLK a_31445_n18723# 6.43e-21
C2671 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.0592f
C2672 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.106f
C2673 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 6.95e-19
C2674 CLK a_35032_n17626# 0.00164f
C2675 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_45458_2768# 1.46e-19
C2676 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0177f
C2677 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.305f
C2678 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 0.00542f
C2679 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00367f
C2680 CLK CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.272f
C2681 RST a_21902_n8787# 7.68e-19
C2682 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_44321_n6273# 1.43e-19
C2683 CLK a_44793_5143# 4.68e-19
C2684 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.122f
C2685 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 1.11e-19
C2686 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.122f
C2687 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT a_28574_n9876# 9.1e-19
C2688 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_29208_10099# 2.96e-19
C2689 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT a_45787_574# 3.92e-20
C2690 VDD96 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.402f
C2691 CLK_div_100_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 7.14e-19
C2692 a_38454_6265# dec3x8_ibr_mag_0.and_3_ibr_6.nand3_mag_ibr_0.OUT 0.0779f
C2693 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 6.95e-19
C2694 CLK_div_108_new_mag_0.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 4.37e-20
C2695 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 7.03e-21
C2696 Vdiv96 Vdiv99 0.0578f
C2697 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 a_53014_n1146# 6.36e-19
C2698 RST CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.0568f
C2699 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 3.77e-20
C2700 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 m3_20882_n11188# 1.57e-20
C2701 VDD96 a_30244_398# 3.56e-19
C2702 VDD100 a_50715_n2243# 0.00123f
C2703 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT a_50833_6284# 0.00378f
C2704 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.374f
C2705 a_23594_n8743# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 4.52e-20
C2706 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT a_36873_n1222# 0.0964f
C2707 a_46810_n10116# m3_20882_n11188# 4.4e-19
C2708 VDD108 CLK_div_108_new_mag_0.JK_FF_mag_1.Q 2.25f
C2709 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.792f
C2710 VDD93 dec3x8_ibr_mag_0.and_3_ibr_5.nand3_mag_ibr_0.OUT 0.0206f
C2711 Vdiv99 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.00136f
C2712 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_44681_n2243# 9.1e-19
C2713 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 9.58e-19
C2714 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 3.09e-19
C2715 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 0.0285f
C2716 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 a_38454_6821# 8.64e-19
C2717 a_36042_6265# a_36202_6265# 0.0504f
C2718 VDD90 a_29772_10099# 3.14e-19
C2719 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.857f
C2720 RST CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_0.OUT 0.00942f
C2721 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_29834_n699# 0.069f
C2722 CLK_div_108_new_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 0.124f
C2723 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 9.67e-20
C2724 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_32015_n17626# 1.5e-20
C2725 Vdiv110 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 0.118f
C2726 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 a_25328_n15535# 4.47e-19
C2727 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_32789_10099# 0.0697f
C2728 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.111f
C2729 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.121f
C2730 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 6.11e-19
C2731 F0 dec3x8_ibr_mag_0.and_3_ibr_5.nand3_mag_ibr_0.OUT 0.344f
C2732 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.0345f
C2733 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 1.06e-19
C2734 Vdiv108 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 7.24e-19
C2735 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN m3_20882_n11188# 0.00612f
C2736 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 a_45075_n9063# 2.79e-20
C2737 VDD90 a_31506_5018# 0.00299f
C2738 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 0.198f
C2739 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN 0.00527f
C2740 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.25f
C2741 CLK dec3x8_ibr_mag_0.and_3_ibr_6.IN3 0.00298f
C2742 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 1.9e-21
C2743 CLK_div_108_new_mag_0.JK_FF_mag_1.QB CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.103f
C2744 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 7.07e-19
C2745 VDD Vdiv90 0.425f
C2746 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT a_50157_n1146# 0.0732f
C2747 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 3.84e-20
C2748 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_26817_n699# 0.00378f
C2749 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 Vdiv99 0.0867f
C2750 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_45570_10154# 1.5e-20
C2751 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 a_54503_1671# 2.79e-20
C2752 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00444f
C2753 VDD96 a_26817_n699# 0.00149f
C2754 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB 0.179f
C2755 RST CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00237f
C2756 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_29187_n15493# 3.12e-19
C2757 VDD96 a_21857_810# 3.14e-19
C2758 VDD105 a_39580_6265# 7.87e-19
C2759 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.273f
C2760 F2 a_39420_6265# 0.00692f
C2761 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT a_50880_10154# 2.88e-20
C2762 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 0.198f
C2763 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.0147f
C2764 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.121f
C2765 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 9.62e-20
C2766 VDD108 a_48466_n6273# 3.73e-19
C2767 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB 0.321f
C2768 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 3.12e-19
C2769 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_26196_5018# 2.88e-20
C2770 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 0.299f
C2771 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.0894f
C2772 Vdiv108 a_44123_n1146# 3e-19
C2773 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_47270_n18696# 0.00876f
C2774 CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_90_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.124f
C2775 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0502f
C2776 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN a_51983_7381# 0.069f
C2777 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB 1.98f
C2778 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 a_29871_n1855# 0.069f
C2779 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT a_48623_n13424# 0.0202f
C2780 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 9.28e-20
C2781 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 Vdiv110 0.0191f
C2782 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.447f
C2783 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_0.Q 0.00211f
C2784 Vdiv96 a_36310_n1822# 5.86e-19
C2785 RST a_47338_n6273# 2.95e-19
C2786 VDD93 a_27850_n9876# 0.00108f
C2787 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT Vdiv110 0.00521f
C2788 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.471f
C2789 VDD105 F0 0.564f
C2790 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.994f
C2791 F0 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT 0.0522f
C2792 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 5.55e-21
C2793 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 2.86e-19
C2794 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_26226_n9831# 0.0036f
C2795 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_29059_6159# 0.0697f
C2796 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00174f
C2797 VDD mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 1.4f
C2798 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 8.16e-20
C2799 CLK CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00118f
C2800 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_44799_n7920# 3.16e-19
C2801 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 5.96e-22
C2802 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 a_47299_10154# 0.0036f
C2803 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 1.05e-20
C2804 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT 0.343f
C2805 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.121f
C2806 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_24938_n9875# 0.0731f
C2807 RST a_28392_354# 0.00217f
C2808 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00118f
C2809 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 1.65f
C2810 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.36f
C2811 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 0.857f
C2812 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.0654f
C2813 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 0.00132f
C2814 CLK_div_108_new_mag_0.JK_FF_mag_1.Q CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 4.18e-21
C2815 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT a_31577_n15535# 0.0203f
C2816 RST Vdiv105 0.00765f
C2817 VDD110 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 1.86e-20
C2818 CLK_div_100_mag_0.CLK_div_10_mag_1.CLK CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.267f
C2819 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_36103_n10028# 1.46e-19
C2820 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_31291_n17626# 8.64e-19
C2821 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 0.783f
C2822 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 a_36310_n1822# 0.00211f
C2823 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT a_47816_6284# 0.00378f
C2824 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 1e-19
C2825 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 a_43718_10154# 0.0157f
C2826 CLK_div_100_mag_0.CLK_div_10_mag_1.CLK a_54509_2768# 0.00164f
C2827 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB a_52769_10154# 0.0811f
C2828 RST a_29059_6159# 1.23e-20
C2829 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.109f
C2830 Vdiv96 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.IN2 0.0205f
C2831 VDD96 a_22982_n2930# 2.21e-19
C2832 VDD105 a_51397_6284# 3.14e-19
C2833 RST CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0633f
C2834 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.768f
C2835 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.391f
C2836 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 dec3x8_ibr_mag_0.and_3_ibr_7.nand3_mag_ibr_0.OUT 0.00277f
C2837 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 4.94e-20
C2838 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_23019_5018# 0.00695f
C2839 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.0286f
C2840 VDD105 a_53120_5143# 0.00727f
C2841 RST a_51652_2768# 0.00186f
C2842 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 0.179f
C2843 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 a_30187_6159# 0.069f
C2844 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0622f
C2845 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 6.69e-19
C2846 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 1.19e-19
C2847 VDD96 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 6.19e-20
C2848 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.0189f
C2849 a_33429_n15491# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 4.52e-20
C2850 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.0725f
C2851 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_48466_n6273# 4.52e-20
C2852 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 a_29110_n743# 3.6e-22
C2853 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 0.121f
C2854 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN 5.82e-21
C2855 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN 7.4e-22
C2856 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_43793_n10116# 0.00964f
C2857 VDD108 m1_42708_4265# 0.0109f
C2858 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT a_47140_n1146# 0.0732f
C2859 a_27850_n9876# m3_20882_n11188# 6.86e-19
C2860 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB a_28016_n8779# 1.33e-20
C2861 CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 3.99e-20
C2862 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_47988_n17599# 3.6e-22
C2863 a_45787_574# CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN 5.1e-20
C2864 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.313f
C2865 VDD dec3x8_ibr_mag_0.and_3_ibr_4.nand3_mag_ibr_0.OUT 0.672f
C2866 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 a_54057_10154# 0.0102f
C2867 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.514f
C2868 a_43719_n120# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00239f
C2869 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB 0.25f
C2870 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_34462_n18723# 0.0202f
C2871 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 a_33583_n16588# 0.0157f
C2872 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_47760_n15585# 0.0195f
C2873 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1f
C2874 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K a_32301_n15491# 1.39e-19
C2875 RST CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.279f
C2876 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.IN2 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 0.00394f
C2877 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT 0.12f
C2878 CLK_div_100_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_54302_n1102# 5.94e-20
C2879 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.205f
C2880 RST a_50987_5143# 0.00186f
C2881 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0576f
C2882 VDD99 a_25420_n13385# 0.165f
C2883 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.395f
C2884 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_35186_n18723# 8.64e-19
C2885 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 5.48e-20
C2886 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.0591f
C2887 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.0132f
C2888 VDD99 a_26052_n15491# 3.14e-19
C2889 RST a_28093_n18723# 1.8e-19
C2890 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.16f
C2891 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 0.00675f
C2892 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 a_28267_n7033# 0.00692f
C2893 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00183f
C2894 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT a_48587_10154# 1.5e-20
C2895 RST CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.213f
C2896 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 1.97e-19
C2897 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 2.1f
C2898 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 3.81e-19
C2899 RST CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.00337f
C2900 Vdiv110 a_39124_880# 6.06e-19
C2901 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.321f
C2902 a_48712_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.00964f
C2903 CLK CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.308f
C2904 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.0106f
C2905 a_52161_n19793# CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.069f
C2906 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 m3_20882_n11188# 0.00222f
C2907 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 7e-19
C2908 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 0.00586f
C2909 CLK_div_90_mag_0.CLK_div_10_mag_0.CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.307f
C2910 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.122f
C2911 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 0.00335f
C2912 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT m3_20882_n11188# 3.02e-19
C2913 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_32175_n17626# 0.0202f
C2914 CLK a_28268_n6266# 2.25e-19
C2915 CLK a_53370_n9020# 6.06e-21
C2916 VDD93 a_31129_n6271# 5.2e-19
C2917 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_26042_6159# 0.0697f
C2918 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.00395f
C2919 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT a_22421_810# 0.00378f
C2920 VDD99 a_28657_n18723# 2.65e-19
C2921 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 8.09e-19
C2922 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 7.11e-21
C2923 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 7.75e-19
C2924 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C2925 CLK_div_96_mag_0.JK_FF_mag_2.Q a_27342_n1855# 0.069f
C2926 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.653f
C2927 CLK a_26980_3016# 0.0017f
C2928 VDD105 a_52951_7381# 3.14e-19
C2929 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00183f
C2930 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 0.00188f
C2931 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_26214_n1855# 1.43e-19
C2932 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 a_22620_n9884# 0.0101f
C2933 CLK CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.013f
C2934 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.395f
C2935 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.0659f
C2936 CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_99_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 3.34e-19
C2937 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 a_30165_n6282# 8.97e-21
C2938 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN 2.97e-19
C2939 a_44734_2768# Vdiv110 5.84e-19
C2940 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.00154f
C2941 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 1.3f
C2942 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C2943 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00183f
C2944 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.107f
C2945 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 m3_20882_n11188# 5.1e-20
C2946 VDD96 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT 0.999f
C2947 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 a_49042_n16682# 0.00372f
C2948 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_47246_5143# 0.0731f
C2949 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.0205f
C2950 a_30050_n13332# a_30210_n13332# 0.0504f
C2951 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00183f
C2952 RST CLK_div_108_new_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.00146f
C2953 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 0.0275f
C2954 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.0592f
C2955 RST a_47914_n16726# 0.00216f
C2956 a_44971_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0203f
C2957 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 a_47835_7960# 2.36e-22
C2958 RST a_49991_n2243# 0.00186f
C2959 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_44436_9057# 0.011f
C2960 VDD mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 0.404f
C2961 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C2962 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0943f
C2963 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C2964 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 0.0302f
C2965 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB 1.96f
C2966 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.266f
C2967 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 a_47988_n17599# 1.04e-19
C2968 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 0.127f
C2969 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 a_45907_n16680# 0.00372f
C2970 F0 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 4.09e-19
C2971 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 a_28828_1497# 0.01f
C2972 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 2.23e-19
C2973 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 5.37e-19
C2974 RST a_21742_n8787# 9.22e-19
C2975 CLK a_44229_5143# 0.00275f
C2976 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_28644_10099# 0.012f
C2977 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT a_28010_n9876# 0.0731f
C2978 CLK_div_96_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN Vdiv96 1e-19
C2979 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.0445f
C2980 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 5.57e-19
C2981 CLK_div_108_new_mag_0.JK_FF_mag_1.QB CLK_div_108_new_mag_0.JK_FF_mag_1.Q 1.96f
C2982 CLK_div_90_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 2.25e-19
C2983 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 0.144f
C2984 a_38294_6265# dec3x8_ibr_mag_0.and_3_ibr_6.nand3_mag_ibr_0.OUT 0.0249f
C2985 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 0.00916f
C2986 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.109f
C2987 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 a_51849_n1102# 0.069f
C2988 VDD96 VDD93 0.591f
C2989 VDD96 a_29680_398# 3.14e-19
C2990 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 3.81e-19
C2991 VDD100 a_50151_n2243# 0.00891f
C2992 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT a_50269_6240# 0.0732f
C2993 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 7.08e-20
C2994 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 5.37e-19
C2995 Vdiv110 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK 0.295f
C2996 VDD dec3x8_ibr_mag_0.and_3_ibr_5.IN3 0.915f
C2997 a_46246_n10116# m3_20882_n11188# 4.57e-19
C2998 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_44117_n2243# 0.0731f
C2999 VDD93 a_37328_6265# 8.68e-19
C3000 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 a_38294_6821# 0.00175f
C3001 a_46755_574# CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN 5.1e-20
C3002 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_25312_5018# 2.81e-19
C3003 VDD90 a_29208_10099# 3.14e-19
C3004 a_47050_n7372# CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 7.48e-20
C3005 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 2.45e-22
C3006 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 3.94e-19
C3007 VDD96 F0 0.117f
C3008 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_31451_n17626# 0.0203f
C3009 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_32225_10099# 0.0059f
C3010 CLK Vdiv 0.284f
C3011 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB 3.49e-19
C3012 F0 a_37328_6265# 0.00193f
C3013 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.198f
C3014 F0 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I1 0.0109f
C3015 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0934f
C3016 VDD90 a_31346_5018# 0.00727f
C3017 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 1.89e-20
C3018 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 3.28e-19
C3019 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 0.109f
C3020 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.802f
C3021 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT a_49997_n1146# 0.0203f
C3022 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN 1.59e-19
C3023 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 m3_20882_n11188# 0.00141f
C3024 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.998f
C3025 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT Vdiv110 2.57e-21
C3026 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_26253_n743# 0.0733f
C3027 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_45006_10154# 0.0203f
C3028 VDD96 a_26253_n743# 9.82e-19
C3029 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB 0.308f
C3030 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.018f
C3031 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 6.69e-19
C3032 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_28623_n15537# 0.00392f
C3033 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 m3_20882_n11188# 0.00101f
C3034 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_43793_n10116# 0.0036f
C3035 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C3036 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 0.00213f
C3037 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1f
C3038 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.121f
C3039 VDD105 a_39420_6265# 0.00132f
C3040 CLK a_33519_11196# 0.00117f
C3041 VDD99 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_0.OUT 2.2e-21
C3042 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 8.16e-20
C3043 CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 8.88e-20
C3044 RST CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.276f
C3045 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 0.00146f
C3046 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00131f
C3047 VDD108 a_47902_n6273# 3.14e-19
C3048 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.792f
C3049 a_26093_n743# CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 9.78e-20
C3050 Vdiv96 a_37999_n1222# 1.35e-19
C3051 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_26036_5018# 9.1e-19
C3052 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN 4.48e-19
C3053 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.00137f
C3054 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.215f
C3055 VDD93 a_24784_n8778# 0.00519f
C3056 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT 0.00134f
C3057 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 1.17e-19
C3058 Vdiv108 a_43963_n1146# 3.71e-19
C3059 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_43760_1671# 4.52e-20
C3060 RST CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0981f
C3061 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB 0.311f
C3062 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_33429_n15491# 0.0114f
C3063 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 1.83e-20
C3064 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.321f
C3065 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.125f
C3066 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.648f
C3067 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 3.43f
C3068 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_90_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 3.38e-19
C3069 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0576f
C3070 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_45449_n6273# 4.52e-20
C3071 Vdiv96 a_35747_n1822# 7.87e-19
C3072 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.125f
C3073 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.0979f
C3074 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 0.0116f
C3075 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT a_39124_880# 0.00949f
C3076 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 0.089f
C3077 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_30342_11196# 1.46e-19
C3078 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.995f
C3079 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 2.02e-20
C3080 VDD99 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 2.2e-20
C3081 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C3082 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 4.42e-19
C3083 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 1.84e-21
C3084 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 8.62e-19
C3085 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.122f
C3086 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0871f
C3087 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.0378f
C3088 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 0.98f
C3089 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 0.407f
C3090 VDD110 Vdiv 0.333f
C3091 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 a_36873_880# 0.00372f
C3092 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 1.99e-20
C3093 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 a_37999_n1222# 0.00375f
C3094 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 a_50204_2768# 0.069f
C3095 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 1.96f
C3096 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 1.96f
C3097 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_24778_n9875# 0.0202f
C3098 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 4.66e-21
C3099 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.514f
C3100 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C3101 RST CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.0112f
C3102 CLK_div_96_mag_0.JK_FF_mag_2.QB CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.25f
C3103 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 a_43760_1671# 0.069f
C3104 F0 mux_8x1_ibr_0.mux_2x1_ibr_0.I0 6.5e-20
C3105 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT 0.745f
C3106 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.298f
C3107 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT m3_20882_n11188# 0.00341f
C3108 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.398f
C3109 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 0.00146f
C3110 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 0.397f
C3111 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 a_35747_n1822# 0.069f
C3112 RST CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.257f
C3113 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0384f
C3114 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT a_47252_6240# 0.0732f
C3115 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 1.31e-20
C3116 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.00335f
C3117 CLK_div_96_mag_0.JK_FF_mag_5.Q CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.269f
C3118 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 2.39e-21
C3119 VDD105 a_50833_6284# 3.14e-19
C3120 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.231f
C3121 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 1.03e-19
C3122 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00836f
C3123 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 a_39580_6265# 6.46e-19
C3124 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT 0.342f
C3125 VDD105 a_52115_5187# 0.00152f
C3126 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.768f
C3127 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 a_43872_9057# 0.069f
C3128 RST a_51492_2768# 0.00186f
C3129 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.321f
C3130 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C3131 RST CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.286f
C3132 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 m3_20882_n11188# 0.0187f
C3133 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 a_28546_n743# 1.86e-20
C3134 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 3.43e-19
C3135 VDD99 Vdiv105 0.348f
C3136 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_32794_5062# 0.0036f
C3137 VDD93 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 0.0388f
C3138 RST a_48017_9057# 1.23e-20
C3139 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_43229_n10116# 0.0811f
C3140 VDD100 Vdiv105 0.289f
C3141 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.0872f
C3142 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.00104f
C3143 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB a_27856_n8779# 1.72e-20
C3144 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT a_46980_n1146# 0.0203f
C3145 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_47424_n17599# 0.00166f
C3146 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 1.14e-19
C3147 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 a_53897_10154# 0.0101f
C3148 CLK CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 0.00254f
C3149 a_43559_n120# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00261f
C3150 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_33898_n18723# 4.52e-20
C3151 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 9.66e-19
C3152 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 1.99e-20
C3153 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 F0 0.368f
C3154 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 a_33019_n16588# 0.00859f
C3155 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K a_31737_n15535# 8.21e-19
C3156 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 0.00146f
C3157 RST a_23289_n6009# 9.7e-19
C3158 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_48478_n16682# 0.00378f
C3159 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.431f
C3160 CLK_div_96_mag_0.JK_FF_mag_4.QB CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 0.0592f
C3161 RST a_50827_5143# 0.00169f
C3162 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN 0.423f
C3163 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0346f
C3164 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 4.92e-21
C3165 RST CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.154f
C3166 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 a_55357_n20487# 2.44e-20
C3167 VDD100 a_51652_2768# 0.0123f
C3168 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.28f
C3169 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 7.16e-20
C3170 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 2.48e-19
C3171 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00153f
C3172 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1f
C3173 RST a_27529_n18723# 7.58e-19
C3174 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.109f
C3175 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_30187_6159# 0.00118f
C3176 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 5.06e-21
C3177 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 5.14e-20
C3178 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I1 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 0.00141f
C3179 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.208f
C3180 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 0.16f
C3181 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 7.04e-20
C3182 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT a_48023_10154# 0.0203f
C3183 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 0.129f
C3184 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 4.26e-19
C3185 a_52225_n13362# a_52385_n13362# 0.186f
C3186 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB 0.0615f
C3187 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 2.64e-19
C3188 Vdiv110 a_38561_880# 4.45e-19
C3189 VDD108 CLK_div_108_new_mag_0.JK_FF_mag_0.QB 0.982f
C3190 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 Vdiv105 3.1e-22
C3191 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.125f
C3192 RST CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.15f
C3193 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 2.33e-20
C3194 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK CLK_div_108_new_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 1e-19
C3195 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_23030_n8743# 4.52e-20
C3196 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_23184_n9840# 0.0036f
C3197 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_25292_10099# 0.0112f
C3198 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_32015_n17626# 0.0731f
C3199 CLK a_52806_n9020# 9.45e-19
C3200 VDD93 a_30165_n6282# 3.14e-19
C3201 CLK CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 0.0385f
C3202 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN 0.517f
C3203 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 1.9e-19
C3204 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.231f
C3205 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 4.27e-20
C3206 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00118f
C3207 Vdiv93 Vdiv99 0.607f
C3208 VDD99 a_28093_n18723# 3.14e-19
C3209 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_36827_n10028# 2.88e-20
C3210 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 1.65f
C3211 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C3212 CLK_div_96_mag_0.JK_FF_mag_2.Q a_26778_n1855# 5.39e-21
C3213 a_33513_10099# F2 3.07e-19
C3214 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.121f
C3215 CLK a_26820_3016# 0.00205f
C3216 VDD105 a_55179_7683# 0.0407f
C3217 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.321f
C3218 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_2.OUT 0.00167f
C3219 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.00252f
C3220 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 3.25e-19
C3221 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 a_22460_n9884# 0.0102f
C3222 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_25650_n1899# 0.00119f
C3223 a_44170_2768# Vdiv110 6.25e-19
C3224 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0343f
C3225 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0576f
C3226 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 6.62e-20
C3227 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00183f
C3228 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 a_48478_n16682# 0.069f
C3229 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_47086_5143# 0.0202f
C3230 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 4.41e-20
C3231 RST CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 0.0232f
C3232 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 1.3f
C3233 RST a_47050_n7372# 3.11e-19
C3234 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_2.OUT a_23869_810# 0.0202f
C3235 RST a_47754_n16726# 0.00199f
C3236 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 2.11e-19
C3237 VDD99 dec3x8_ibr_mag_0.and_3_ibr_2.nand3_mag_ibr_0.OUT 8.8e-19
C3238 a_44971_n17599# a_45131_n17599# 0.0504f
C3239 a_44407_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1.5e-20
C3240 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT m3_20882_n11188# 0.00137f
C3241 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 0.109f
C3242 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.103f
C3243 RST a_48986_n2199# 9.66e-19
C3244 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_43872_9057# 0.00118f
C3245 RST CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_0.OUT 0.0145f
C3246 VDD100 dec3x8_ibr_mag_0.and_3_ibr_2.nand3_mag_ibr_0.OUT 0.145f
C3247 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_32169_n18723# 0.0203f
C3248 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 a_28267_n7033# 0.00347f
C3249 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.122f
C3250 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 3.49e-19
C3251 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.00288f
C3252 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.122f
C3253 a_30164_n7017# CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 8.97e-21
C3254 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 a_45343_n16680# 0.069f
C3255 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.00169f
C3256 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 1.55e-19
C3257 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB 3.09e-19
C3258 a_47086_5143# a_47246_5143# 0.0504f
C3259 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.00252f
C3260 CLK_div_105_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_43831_7266# 9.16e-20
C3261 a_29213_n7028# CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 4.18e-21
C3262 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN a_30164_n7017# 1.05e-20
C3263 CLK a_44069_5143# 0.00228f
C3264 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT a_27850_n9876# 0.0202f
C3265 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 a_29801_1733# 8.64e-19
C3266 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN m3_20882_n11188# 0.00669f
C3267 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.186f
C3268 a_38294_6265# a_38454_6265# 0.0504f
C3269 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.163f
C3270 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.46e-20
C3271 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 9.64e-19
C3272 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT 0.00718f
C3273 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.122f
C3274 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 2.71e-21
C3275 VDD96 a_29116_398# 3.14e-19
C3276 VDD100 a_49991_n2243# 0.0132f
C3277 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT a_50109_6240# 0.0203f
C3278 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.198f
C3279 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.211f
C3280 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00183f
C3281 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_25508_n8734# 4.61e-20
C3282 a_22839_10099# CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 4.9e-20
C3283 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_2.OUT 0.00164f
C3284 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.913f
C3285 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_27170_6159# 0.00118f
C3286 VDD93 a_37168_6265# 0.00148f
C3287 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_43957_n2243# 0.0202f
C3288 a_45241_n10160# m3_20882_n11188# 0.00102f
C3289 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.999f
C3290 VDD90 a_28644_10099# 3.56e-19
C3291 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 7.22e-20
C3292 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_31291_n17626# 0.0733f
C3293 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 0.493f
C3294 VDD93 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_1.IN2 5.56e-19
C3295 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK 2.93f
C3296 Vdiv108 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00335f
C3297 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 7.08e-20
C3298 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_47374_n10160# 8.64e-19
C3299 a_51487_n10161# a_51647_n10161# 0.0504f
C3300 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 0.00205f
C3301 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 8.16e-20
C3302 F0 a_37168_6265# 0.00181f
C3303 VDD90 a_30341_5062# 0.00152f
C3304 F0 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_1.IN2 0.368f
C3305 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB a_29708_n8735# 0.0114f
C3306 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 7.57e-20
C3307 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_26093_n743# 0.0203f
C3308 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.359f
C3309 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 a_53375_1671# 6.06e-21
C3310 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_44846_10154# 0.0733f
C3311 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN 0.517f
C3312 VDD96 a_26093_n743# 0.0012f
C3313 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 6.82e-19
C3314 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 7.49e-20
C3315 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.16f
C3316 CLK a_33359_11196# 0.00164f
C3317 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0569f
C3318 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.11f
C3319 VDD108 a_47338_n6273# 3.14e-19
C3320 Vdiv96 a_36873_n1222# 0.00641f
C3321 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_25472_5018# 0.0731f
C3322 a_44475_n5176# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.00696f
C3323 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.001f
C3324 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_45618_2768# 1.17e-20
C3325 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 2.33e-20
C3326 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_96_mag_0.JK_FF_mag_2.Q 1.11e-19
C3327 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 2.22e-20
C3328 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.0894f
C3329 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_32865_n15491# 2.96e-19
C3330 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.JK_FF_mag_5.QB 2.73e-21
C3331 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.0615f
C3332 VDD96 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.391f
C3333 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT a_46755_574# 0.00138f
C3334 VDD93 a_23283_n7106# 0.00523f
C3335 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 0.0204f
C3336 Vdiv105 F2 0.092f
C3337 Vdiv96 a_35184_n1822# 5.86e-19
C3338 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 8.58e-20
C3339 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.397f
C3340 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_44117_n2243# 1.46e-19
C3341 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 0.00205f
C3342 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 a_48466_n6273# 0.069f
C3343 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN 3.08e-19
C3344 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_30209_7256# 5.1e-20
C3345 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00157f
C3346 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.768f
C3347 Vdiv99 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00154f
C3348 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT a_38561_880# 9.46e-19
C3349 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0432f
C3350 VDD108 Vdiv105 1.96f
C3351 VDD110 a_54022_n17599# 2.21e-19
C3352 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 0.11f
C3353 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 3.26e-20
C3354 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK m3_20882_n11188# 0.00276f
C3355 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 0.0285f
C3356 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_96_mag_0.JK_FF_mag_2.QB 2.7e-19
C3357 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 a_36310_880# 0.069f
C3358 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 a_36873_n1222# 8.2e-19
C3359 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 a_49640_2768# 0.00372f
C3360 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_52293_n17599# 0.0157f
C3361 CLK_div_90_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 Vdiv90 0.028f
C3362 a_53249_n6862# CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K 2.59e-19
C3363 RST CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN 0.147f
C3364 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 0.0593f
C3365 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.36f
C3366 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_48258_n10160# 1.17e-20
C3367 VDD105 a_48741_9057# 0.00746f
C3368 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.395f
C3369 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 0.0285f
C3370 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.25f
C3371 CLK CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 0.149f
C3372 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT a_47092_6240# 0.0203f
C3373 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.0758f
C3374 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK 0.0159f
C3375 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00152f
C3376 VDD96 a_22258_n2930# 0.00108f
C3377 VDD105 a_50269_6240# 2.66e-19
C3378 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 a_39420_6265# 5.51e-19
C3379 VDD105 a_51551_5187# 0.00152f
C3380 Vdiv96 a_35184_880# 2.98e-21
C3381 CLK_div_90_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 1.29e-19
C3382 RST a_50928_2768# 0.00169f
C3383 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 2.66e-19
C3384 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0894f
C3385 a_43895_n16724# a_44055_n16724# 0.0504f
C3386 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 a_39684_n10028# 3.6e-22
C3387 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 7.32e-20
C3388 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.108f
C3389 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN 0.00185f
C3390 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 4.27e-20
C3391 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT 0.122f
C3392 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00153f
C3393 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 a_28386_n743# 2.55e-20
C3394 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.00123f
C3395 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 8.58e-20
C3396 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 0.389f
C3397 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 0.391f
C3398 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 0.198f
C3399 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 a_44436_9057# 0.069f
C3400 CLK_div_96_mag_0.JK_FF_mag_0.Q CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.235f
C3401 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 1.56e-21
C3402 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_47264_n17599# 0.001f
C3403 VDD a_36042_6265# 2.21e-19
C3404 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 a_53333_10154# 0.00859f
C3405 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 4.84e-19
C3406 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.121f
C3407 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.806f
C3408 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_3.Q 0.00292f
C3409 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 a_32455_n16632# 0.0101f
C3410 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.656f
C3411 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K a_31577_n15535# 0.00598f
C3412 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_47914_n16726# 0.0733f
C3413 RST a_23129_n6009# 9.7e-19
C3414 RST a_50263_5143# 0.00186f
C3415 VDD99 a_23956_n14213# 3.14e-19
C3416 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.431f
C3417 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 a_55197_n20487# 9.02e-19
C3418 RST CLK 17.7f
C3419 CLK_div_108_new_mag_0.JK_FF_mag_1.QB CLK_div_108_new_mag_0.JK_FF_mag_0.QB 4.17e-22
C3420 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_54592_n18696# 0.0059f
C3421 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB 9.14e-19
C3422 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.JK_FF_mag_1.Q 0.0343f
C3423 VDD100 a_51492_2768# 0.00863f
C3424 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN 0.124f
C3425 F2 dec3x8_ibr_mag_0.and_3_ibr_2.nand3_mag_ibr_0.OUT 0.354f
C3426 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.995f
C3427 VDD99 a_25328_n15535# 2.21e-19
C3428 RST a_26965_n18723# 7.24e-19
C3429 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 0.447f
C3430 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00718f
C3431 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_29623_6159# 0.011f
C3432 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 0.175f
C3433 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.IN1 a_32750_n7675# 0.0144f
C3434 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.648f
C3435 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT a_47863_10154# 0.0733f
C3436 CLK_div_96_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 0.124f
C3437 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 0.00118f
C3438 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT 0.768f
C3439 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT 1.01e-19
C3440 RST a_54664_n10161# 0.00218f
C3441 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN a_25420_n13385# 2.4e-20
C3442 Vdiv93 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 0.00133f
C3443 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 1.16f
C3444 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT 0.0951f
C3445 Vdiv90 Vdiv100 0.0176f
C3446 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C3447 RST CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.00698f
C3448 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 6.25e-19
C3449 Vdiv110 a_37999_880# 6.06e-19
C3450 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN 0.0123f
C3451 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 0.0124f
C3452 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 2.34e-19
C3453 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C3454 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 0.122f
C3455 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 4.24e-20
C3456 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.0264f
C3457 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_22466_n8743# 0.0202f
C3458 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_31451_n17626# 9.1e-19
C3459 CLK_div_100_mag_0.CLK_div_10_mag_1.CLK a_55067_297# 0.198f
C3460 CLK a_51641_n9064# 0.0101f
C3461 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 1.17e-19
C3462 CLK_div_108_new_mag_0.CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT 2.34e-19
C3463 VDD93 a_29214_n6271# 3.14e-19
C3464 Vdiv93 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 2.91e-19
C3465 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.16f
C3466 Vdiv96 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 0.0775f
C3467 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 1.3f
C3468 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_25482_n16632# 8.66e-20
C3469 VDD99 a_27529_n18723# 3.14e-19
C3470 RST CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.336f
C3471 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00167f
C3472 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_36667_n10028# 9.1e-19
C3473 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.103f
C3474 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K a_49488_n13383# 2.5e-19
C3475 RST CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 0.00927f
C3476 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.469f
C3477 VDD105 a_55019_7683# 0.234f
C3478 a_48944_6284# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 4.52e-20
C3479 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT 1.19f
C3480 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 a_21896_n9884# 0.00789f
C3481 RST CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.00661f
C3482 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 4.22e-20
C3483 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 0.00145f
C3484 a_45000_9057# CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT 5.94e-20
C3485 a_25312_5018# a_25472_5018# 0.0504f
C3486 a_43606_2768# Vdiv110 6.45e-19
C3487 Vdiv108 a_55020_n2199# 7.51e-19
C3488 a_47723_574# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 7.43e-22
C3489 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_45612_1671# 0.0203f
C3490 CLK CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 1.32f
C3491 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_2.OUT a_23709_810# 0.0731f
C3492 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.00104f
C3493 RST a_47190_n16726# 0.00257f
C3494 a_44247_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1.17e-20
C3495 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 6.02e-20
C3496 VDD110 RST 2.78f
C3497 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 6.82e-19
C3498 RST a_48422_n2199# 9.41e-19
C3499 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB a_35026_n18723# 0.00392f
C3500 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN 5.7e-20
C3501 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 Vdiv100 0.217f
C3502 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 a_48324_n15585# 0.0059f
C3503 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_32009_n18723# 0.0732f
C3504 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 0.0112f
C3505 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 0.0189f
C3506 RST a_32225_10099# 3.62e-19
C3507 RST CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 0.0507f
C3508 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 a_26343_n7107# 5.54e-19
C3509 RST CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 0.00356f
C3510 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_44170_2768# 0.0036f
C3511 Vdiv93 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 0.00233f
C3512 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0568f
C3513 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT 0.338f
C3514 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 a_51034_9057# 0.0697f
C3515 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 3.4e-19
C3516 CLK_div_105_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_43671_7266# 5.39e-20
C3517 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 7.24e-19
C3518 CLK a_33358_5062# 6.21e-19
C3519 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 2.47e-20
C3520 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 8.2e-19
C3521 CLK CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 1.22e-19
C3522 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN 0.146f
C3523 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_2.Q 0.0179f
C3524 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 3.45e-19
C3525 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_30025_n2952# 0.0036f
C3526 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT 1.74e-19
C3527 VDD100 a_48986_n2199# 0.00152f
C3528 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 0.281f
C3529 F2 mux_8x1_ibr_0.mux_2x1_ibr_0.I1 0.0639f
C3530 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB 0.911f
C3531 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C3532 a_45081_n10160# m3_20882_n11188# 0.00102f
C3533 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_26606_6159# 0.011f
C3534 CLK a_53458_n17599# 1.84e-20
C3535 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.0172f
C3536 a_45570_10154# a_45730_10154# 0.0504f
C3537 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT 0.00183f
C3538 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_30727_n17626# 0.00378f
C3539 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_30760_n20290# 1.4e-19
C3540 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00252f
C3541 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 a_30315_n15493# 0.069f
C3542 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT m3_20882_n11188# 0.00134f
C3543 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 0.0655f
C3544 CLK CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 1.46e-19
C3545 Vdiv100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 8.11e-20
C3546 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN 0.0829f
C3547 VDD90 a_29777_5062# 0.00152f
C3548 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 a_43383_n9019# 0.069f
C3549 CLK_div_96_mag_0.JK_FF_mag_2.QB a_27496_n2952# 0.0811f
C3550 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN a_31129_n6271# 0.069f
C3551 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.304f
C3552 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 a_52161_n19793# 1.29e-22
C3553 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.348f
C3554 RST CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.0251f
C3555 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB a_29144_n8735# 2.96e-19
C3556 CLK_div_96_mag_0.JK_FF_mag_0.QB CLK_div_96_mag_0.JK_FF_mag_0.Q 1.95f
C3557 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 0.0334f
C3558 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_25529_n743# 1.5e-20
C3559 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.109f
C3560 VDD93 a_29708_n8735# 3.56e-19
C3561 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_44282_10154# 0.00378f
C3562 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 a_52811_1671# 0.069f
C3563 VDD96 a_25529_n743# 0.00888f
C3564 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00356f
C3565 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.313f
C3566 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT 1.29e-19
C3567 CLK CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.27f
C3568 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_45000_9057# 0.0202f
C3569 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.0378f
C3570 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 2.32e-19
C3571 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_27375_n17626# 0.069f
C3572 Vdiv96 a_35747_n1222# 0.00347f
C3573 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 8.59e-20
C3574 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_25312_5018# 0.0202f
C3575 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT a_51647_n10161# 0.0202f
C3576 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_45039_n5176# 0.00378f
C3577 a_44315_n5176# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.00695f
C3578 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT Vdiv90 6.02e-19
C3579 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.01e-19
C3580 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_45075_n9063# 0.00392f
C3581 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_45458_2768# 1.5e-20
C3582 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C3583 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_32301_n15491# 3.08e-19
C3584 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 2.45e-19
C3585 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 0.888f
C3586 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT a_43719_n120# 0.0294f
C3587 VDD105 Vdiv105 0.156f
C3588 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 9.58e-20
C3589 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 1.32e-19
C3590 VDD96 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.742f
C3591 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.00183f
C3592 Vdiv105 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT 1.33e-19
C3593 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 0.198f
C3594 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 Vdiv96 0.011f
C3595 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.338f
C3596 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_29241_7256# 0.069f
C3597 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 0.0635f
C3598 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT a_37999_880# 0.00949f
C3599 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0334f
C3600 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00243f
C3601 VDD110 a_53458_n17599# 0.00299f
C3602 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 2.86e-19
C3603 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_24938_n9875# 1.46e-19
C3604 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 0.203f
C3605 VDD108 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.997f
C3606 a_25640_n18723# a_25800_n18723# 0.0504f
C3607 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.36f
C3608 CLK_div_90_mag_0.CLK_div_10_mag_0.CLK CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.129f
C3609 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.257f
C3610 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 1.96f
C3611 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN 0.112f
C3612 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0596f
C3613 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 a_35747_n1222# 1.5e-19
C3614 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_51729_n17599# 0.00859f
C3615 CLK_div_90_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 a_33405_7558# 2.44e-20
C3616 a_53089_n6862# CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K 2.59e-19
C3617 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT 0.117f
C3618 Vdiv99 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN 3.87e-19
C3619 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.0215f
C3620 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN a_43383_n9019# 4.94e-20
C3621 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.209f
C3622 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 0.414f
C3623 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_54456_n2199# 0.00378f
C3624 RST CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 0.0395f
C3625 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_48098_n10160# 1.5e-20
C3626 VDD105 a_48581_9057# 2.66e-19
C3627 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.121f
C3628 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00164f
C3629 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.00384f
C3630 CLK_div_96_mag_0.JK_FF_mag_5.Q CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 3.64e-19
C3631 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 5.45e-20
C3632 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 2f
C3633 Vdiv100 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 0.0499f
C3634 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.431f
C3635 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_51005_n17599# 3.6e-22
C3636 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_52385_n13362# 1.9e-19
C3637 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K 6.15e-20
C3638 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 2.79e-20
C3639 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0385f
C3640 VDD105 a_50109_6240# 0.00746f
C3641 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 0.25f
C3642 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.00157f
C3643 VDD105 a_50987_5143# 0.00101f
C3644 RST a_50768_2768# 0.00186f
C3645 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 a_28495_6115# 2.79e-20
C3646 a_25322_n16632# a_25482_n16632# 0.0504f
C3647 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_48092_n9063# 0.00119f
C3648 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K 1.41e-20
C3649 Vdiv110 a_39124_280# 2.66e-19
C3650 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 a_39120_n10028# 1.86e-20
C3651 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_44357_n10160# 8.64e-19
C3652 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT m3_20882_n11188# 0.00187f
C3653 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.103f
C3654 a_28577_n2996# a_28737_n2996# 0.0504f
C3655 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB 0.186f
C3656 CLK_div_96_mag_0.JK_FF_mag_3.Q a_25490_n1899# 3.77e-20
C3657 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.103f
C3658 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN 0.515f
C3659 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 a_27381_n699# 0.0157f
C3660 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 8.58e-20
C3661 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 3.38e-19
C3662 VDD93 a_26349_n6010# 0.00108f
C3663 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.076f
C3664 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.161f
C3665 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 a_43872_9057# 0.00372f
C3666 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.768f
C3667 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.0622f
C3668 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 a_52769_10154# 0.0157f
C3669 a_25619_n7107# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 4.61e-20
C3670 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.395f
C3671 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_50829_n6865# 8.64e-19
C3672 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 a_32295_n16632# 0.0102f
C3673 RST a_47816_6284# 1.23e-20
C3674 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 1.89e-19
C3675 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 5.37e-19
C3676 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_47754_n16726# 0.0203f
C3677 a_25490_n1899# a_25650_n1899# 0.0504f
C3678 RST a_22565_n6009# 0.00155f
C3679 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 2.25e-19
C3680 RST a_50103_5143# 0.00186f
C3681 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0334f
C3682 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_30502_11196# 1.17e-20
C3683 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 a_21841_n6009# 0.069f
C3684 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 7.81e-19
C3685 VDD105 dec3x8_ibr_mag_0.and_3_ibr_2.nand3_mag_ibr_0.OUT 0.0274f
C3686 VDD100 a_50928_2768# 0.00123f
C3687 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT 0.00147f
C3688 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_54028_n18696# 0.0697f
C3689 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.14f
C3690 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 5.2e-20
C3691 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB 1.99f
C3692 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.103f
C3693 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_29059_6159# 1.43e-19
C3694 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00264f
C3695 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT a_47299_10154# 0.00378f
C3696 RST a_54504_n10161# 0.00218f
C3697 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN 0.00165f
C3698 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.026f
C3699 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 0.00209f
C3700 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 5.2e-20
C3701 a_47835_7960# CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 2.48e-19
C3702 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.107f
C3703 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00157f
C3704 Vdiv110 a_37436_880# 4.45e-19
C3705 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT a_51758_9057# 0.0203f
C3706 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.JK_FF_mag_2.Q 0.16f
C3707 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT 0.00395f
C3708 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_0.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 5.23e-20
C3709 CLK_div_108_new_mag_0.JK_FF_mag_1.Q CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT 9.01e-22
C3710 VDD96 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_0.OUT 0.746f
C3711 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 1.32e-19
C3712 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 a_29213_n7028# 0.0114f
C3713 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_31291_n17626# 2.88e-20
C3714 CLK_div_100_mag_0.CLK_div_10_mag_1.CLK a_54907_297# 0.0133f
C3715 CLK a_51481_n9064# 0.00939f
C3716 VDD99 CLK 6.14f
C3717 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 a_33358_5062# 0.0157f
C3718 VDD100 CLK 2.51f
C3719 Vdiv90 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 5.13e-20
C3720 RST CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.317f
C3721 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.0435f
C3722 VDD99 a_26965_n18723# 3.56e-19
C3723 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.092f
C3724 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 0.391f
C3725 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 CLK_div_105_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00357f
C3726 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_36103_n10028# 0.0731f
C3727 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN 7e-19
C3728 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_2.OUT CLK_div_96_mag_0.JK_FF_mag_4.Q 0.338f
C3729 VDD108 a_47050_n7372# 5.92e-19
C3730 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 2.11e-20
C3731 CLK_div_96_mag_0.JK_FF_mag_2.Q a_25650_n1899# 2.79e-20
C3732 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 0.0444f
C3733 RST CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.0758f
C3734 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 1.77e-19
C3735 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.122f
C3736 VDD105 a_51983_7381# 3.14e-19
C3737 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 3.18e-19
C3738 Vdiv99 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN 9.83e-19
C3739 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.00559f
C3740 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.103f
C3741 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 a_21736_n9884# 0.00335f
C3742 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_45241_n10160# 1.17e-20
C3743 RST a_29213_n7028# 3.66e-19
C3744 CLK CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.00364f
C3745 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 9.6e-19
C3746 Vdiv108 a_54456_n2199# 7.3e-19
C3747 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_45452_1671# 0.0732f
C3748 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_45753_n15583# 0.069f
C3749 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT a_51871_n5# 0.00138f
C3750 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.101f
C3751 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00229f
C3752 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.457f
C3753 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_2.OUT a_23145_810# 9.1e-19
C3754 RST a_47030_n16726# 0.00257f
C3755 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.321f
C3756 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.122f
C3757 RST a_47858_n2243# 0.00186f
C3758 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_45075_n9063# 0.00119f
C3759 RST CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 3.84e-20
C3760 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 3.76e-19
C3761 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 1.34e-19
C3762 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT 1.48e-19
C3763 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB a_34462_n18723# 3.33e-19
C3764 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.002f
C3765 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.0014f
C3766 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 a_47760_n15585# 0.0697f
C3767 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1f
C3768 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_2.OUT 0.235f
C3769 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_31445_n18723# 0.00378f
C3770 RST CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.145f
C3771 RST a_31661_10099# 7.24e-19
C3772 Vdiv105 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 1.08e-19
C3773 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 a_54504_n10161# 1.46e-19
C3774 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.0509f
C3775 F1 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT 0.112f
C3776 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 a_26183_n7107# 4.21e-19
C3777 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.16f
C3778 a_44075_6240# a_44235_6240# 0.0504f
C3779 CLK CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 6.62e-20
C3780 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 2.42f
C3781 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 4.44e-20
C3782 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 a_27334_n16588# 0.0157f
C3783 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_23594_n8743# 2.21e-19
C3784 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 1.31e-20
C3785 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 1.53e-19
C3786 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 a_50470_9057# 0.0059f
C3787 a_54669_2768# Vdiv110 0.00138f
C3788 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.103f
C3789 CLK a_32794_5062# 6.02e-19
C3790 RST CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.337f
C3791 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 0.0693f
C3792 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 5.97e-20
C3793 Vdiv110 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT 0.00565f
C3794 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.298f
C3795 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 0.149f
C3796 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 a_50157_n1146# 2.79e-20
C3797 VDD100 VDD110 0.085f
C3798 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_2.OUT CLK_div_96_mag_0.JK_FF_mag_5.Q 0.338f
C3799 VDD96 a_28392_354# 2.21e-19
C3800 VDD100 a_48422_n2199# 0.00152f
C3801 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.00183f
C3802 Vdiv93 a_35184_n1822# 0.00347f
C3803 Vdiv110 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT 0.00625f
C3804 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 6.24e-19
C3805 RST CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 0.163f
C3806 VDD96 Vdiv105 0.00374f
C3807 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.0654f
C3808 CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 0.00132f
C3809 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_26042_6159# 1.43e-19
C3810 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.0126f
C3811 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 0.00125f
C3812 a_44517_n10160# m3_20882_n11188# 4.29e-19
C3813 VDD100 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 0.0164f
C3814 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.00118f
C3815 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_37955_n9984# 0.0811f
C3816 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT a_39124_280# 0.0964f
C3817 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C3818 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C3819 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 1.03f
C3820 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 0.122f
C3821 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.00154f
C3822 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 Vdiv110 2.4e-20
C3823 CLK CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.235f
C3824 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 0.122f
C3825 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C3826 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 0.124f
C3827 VDD90 a_29213_5018# 0.00101f
C3828 CLK_div_96_mag_0.JK_FF_mag_2.QB a_26932_n2952# 0.00964f
C3829 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 4.44e-20
C3830 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 2.51e-19
C3831 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB a_28580_n8735# 3.33e-19
C3832 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT m3_20882_n11188# 1.22e-19
C3833 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 0.994f
C3834 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_25369_n743# 1.17e-20
C3835 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 1.49e-19
C3836 VDD93 a_29144_n8735# 3.14e-19
C3837 VDD96 a_25369_n743# 0.0133f
C3838 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 a_47835_7960# 0.0105f
C3839 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT 8.36e-19
C3840 F1 a_37328_6821# 0.00993f
C3841 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 dec3x8_ibr_mag_0.and_3_ibr_4.nand3_mag_ibr_0.OUT 0.133f
C3842 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN 0.112f
C3843 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00943f
C3844 CLK_div_96_mag_0.JK_FF_mag_2.QB CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.103f
C3845 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_44436_9057# 4.52e-20
C3846 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.25f
C3847 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C3848 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.395f
C3849 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_26811_n17626# 0.00372f
C3850 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT a_51487_n10161# 0.0731f
C3851 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.998f
C3852 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.177f
C3853 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_44511_n9019# 1.75e-19
C3854 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_44894_2768# 0.0203f
C3855 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_31737_n15535# 0.00392f
C3856 CLK_div_100_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 3.87e-19
C3857 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 a_37999_280# 0.00372f
C3858 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT a_43559_n120# 0.00894f
C3859 VDD93 a_22559_n7106# 3.14e-19
C3860 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.0072f
C3861 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_29054_11196# 0.0036f
C3862 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 0.00233f
C3863 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.0661f
C3864 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 9.64e-20
C3865 VDD110 a_53298_n17599# 0.00727f
C3866 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 4.49e-20
C3867 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 0.342f
C3868 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0834f
C3869 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 0.177f
C3870 CLK CLK_div_100_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 7.44e-19
C3871 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB a_26072_n8734# 4.61e-20
C3872 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 1.32f
C3873 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.414f
C3874 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 1.1e-19
C3875 Vdiv93 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 3.78e-20
C3876 CLK_div_90_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 a_33245_7558# 9.02e-19
C3877 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 a_22711_n14504# 1.75e-19
C3878 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 3.56e-19
C3879 VDD96 dec3x8_ibr_mag_0.and_3_ibr_2.nand3_mag_ibr_0.OUT 0.031f
C3880 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 a_50715_n2243# 3.6e-22
C3881 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.019f
C3882 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_31451_n17626# 0.00695f
C3883 VDD90 a_23691_9000# 5.92e-19
C3884 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_53892_n2243# 0.0733f
C3885 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_47534_n10160# 0.0203f
C3886 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_46105_n18696# 0.00372f
C3887 VDD105 a_48017_9057# 3.14e-19
C3888 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN 0.299f
C3889 CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.00124f
C3890 a_23948_n18723# CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 4.94e-20
C3891 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_50441_n17599# 0.00166f
C3892 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 3.89e-20
C3893 VDD105 a_48944_6284# 3.56e-19
C3894 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.655f
C3895 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_26253_n743# 8.64e-19
C3896 VDD105 a_50827_5143# 0.00123f
C3897 RST a_50204_2768# 9.41e-19
C3898 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.108f
C3899 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_47528_n9019# 1.43e-19
C3900 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_25076_n18723# 0.0697f
C3901 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.065f
C3902 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT m3_20882_n11188# 0.00166f
C3903 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 a_38960_n10028# 2.55e-20
C3904 CLK F2 0.472f
C3905 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.654f
C3906 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00169f
C3907 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 2.17e-21
C3908 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 Vdiv110 0.00367f
C3909 RST CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.143f
C3910 a_44681_n2243# a_44841_n2243# 0.0504f
C3911 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.338f
C3912 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 5.18e-20
C3913 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 a_26817_n699# 0.00859f
C3914 RST CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN 9.43e-19
C3915 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_31506_5018# 1.46e-19
C3916 VDD99 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 0.0151f
C3917 VDD108 CLK 3.88f
C3918 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 1.76e-20
C3919 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.21f
C3920 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 0.00586f
C3921 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00917f
C3922 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 4e-19
C3923 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 a_26814_1919# 0.00119f
C3924 a_25502_n9875# a_25662_n9875# 0.0504f
C3925 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 a_31731_n16632# 0.00789f
C3926 VDD108 a_54664_n10161# 0.0132f
C3927 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 0.00995f
C3928 RST a_22405_n6009# 0.00127f
C3929 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_47190_n16726# 1.5e-20
C3930 CLK CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 0.00361f
C3931 RST a_49098_5187# 9.66e-19
C3932 a_44888_1671# CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT 5.94e-20
C3933 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 0.564f
C3934 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 0.995f
C3935 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_30342_11196# 1.5e-20
C3936 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 1.23e-20
C3937 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.647f
C3938 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 a_21277_n6009# 0.00372f
C3939 VDD100 a_50768_2768# 0.00101f
C3940 CLK_div_108_new_mag_0.CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 3.34e-19
C3941 CLK_div_96_mag_0.JK_FF_mag_2.QB CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 3e-19
C3942 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK a_53469_n15631# 1.88e-19
C3943 RST CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.00289f
C3944 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 8.93e-19
C3945 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 2.95e-20
C3946 CLK_div_105_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 4.25e-20
C3947 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_28495_6115# 0.00119f
C3948 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 0.198f
C3949 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 0.0174f
C3950 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 mux_8x1_ibr_0.mux_2x1_ibr_0.I1 0.109f
C3951 VDD110 a_53304_n18696# 2.21e-19
C3952 RST a_53940_n10161# 0.00187f
C3953 dec3x8_ibr_mag_0.and_3_ibr_5.IN3 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 0.546f
C3954 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 0.231f
C3955 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.496f
C3956 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT a_51598_9057# 0.0732f
C3957 CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 4.44e-20
C3958 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_51646_1671# 0.00876f
C3959 Vdiv110 a_36873_880# 6.06e-19
C3960 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_51957_n6821# 0.00372f
C3961 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.36f
C3962 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 a_47698_n2243# 3.6e-22
C3963 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 m3_20882_n11188# 8.73e-19
C3964 CLK_div_96_mag_0.JK_FF_mag_0.QB CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.103f
C3965 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 0.0432f
C3966 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.303f
C3967 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_21896_n9884# 1.46e-19
C3968 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 7.24e-20
C3969 CLK a_50917_n9020# 6.43e-21
C3970 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0854f
C3971 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 9.55e-20
C3972 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.28f
C3973 F1 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 2.44e-19
C3974 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.321f
C3975 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.447f
C3976 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 1.82e-19
C3977 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN 2.39e-20
C3978 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 a_32794_5062# 0.00859f
C3979 VDD110 F2 0.0129f
C3980 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 0.177f
C3981 CLK_div_105_mag_0.CLK_div_10_mag_1.CLK a_54781_10154# 0.00117f
C3982 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_35943_n10028# 0.0202f
C3983 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 0.0145f
C3984 VDD108 a_43826_n7684# 0.165f
C3985 VDD105 a_51015_7381# 6e-19
C3986 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.321f
C3987 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_0.Q 0.0343f
C3988 CLK_div_96_mag_0.JK_FF_mag_0.QB CLK_div_96_mag_0.JK_FF_mag_2.QB 6.67e-20
C3989 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.122f
C3990 VDD108 VDD110 0.236f
C3991 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.0285f
C3992 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_45081_n10160# 1.5e-20
C3993 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.496f
C3994 RST CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.272f
C3995 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0835f
C3996 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 CLK_div_100_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00357f
C3997 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB 2.42e-20
C3998 Vdiv108 a_53892_n2243# 6.67e-19
C3999 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_44888_1671# 0.00378f
C4000 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 0.399f
C4001 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_47190_n16726# 4.52e-19
C4002 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 0.392f
C4003 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 0.396f
C4004 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_2.OUT a_22985_810# 2.88e-20
C4005 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 5.48f
C4006 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 8.04e-19
C4007 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 4.19e-20
C4008 RST a_45907_n16680# 0.00154f
C4009 CLK CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 0.00302f
C4010 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_44511_n9019# 1.43e-19
C4011 RST a_47698_n2243# 0.00169f
C4012 F0 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT 0.0515f
C4013 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 dec3x8_ibr_mag_0.and_3_ibr_2.nand3_mag_ibr_0.OUT 0.329f
C4014 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.643f
C4015 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.198f
C4016 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.25f
C4017 VDD99 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 1.08e-20
C4018 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0334f
C4019 dec3x8_ibr_mag_0.and_3_ibr_5.IN3 a_36202_6821# 0.00903f
C4020 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 0.0127f
C4021 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00397f
C4022 dec3x8_ibr_mag_0.and_3_ibr_0.nand3_mag_ibr_0.OUT F1 5.08e-19
C4023 CLK a_30496_10099# 0.0101f
C4024 RST CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 4.25e-20
C4025 Vdiv110 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 3.32e-19
C4026 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 5.55e-21
C4027 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT a_51011_n18696# 0.00378f
C4028 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 a_26770_n16588# 0.00859f
C4029 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.0591f
C4030 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.657f
C4031 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00137f
C4032 a_54509_2768# Vdiv110 0.00138f
C4033 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 a_30187_6159# 0.00372f
C4034 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K a_30315_n15493# 8.11e-19
C4035 CLK a_32230_5018# 5.65e-19
C4036 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 0.233f
C4037 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 0.00975f
C4038 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.00125f
C4039 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB a_48023_10154# 0.00695f
C4040 a_51592_n16680# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 4.81e-20
C4041 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 0.0655f
C4042 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_45189_n15583# 4.52e-20
C4043 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 3.85e-20
C4044 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 0.538f
C4045 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 0.994f
C4046 VDD96 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.409f
C4047 RST CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.337f
C4048 VDD100 a_47858_n2243# 0.00101f
C4049 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_23030_n8743# 0.0059f
C4050 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 0.0398f
C4051 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_25478_6115# 0.00119f
C4052 a_44357_n10160# m3_20882_n11188# 4.29e-19
C4053 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 6.94e-19
C4054 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.765f
C4055 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00118f
C4056 a_43559_n120# a_43719_n120# 0.186f
C4057 Vdiv96 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 0.00794f
C4058 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_37391_n9984# 0.00964f
C4059 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C4060 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.321f
C4061 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 8.16e-20
C4062 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK 0.00774f
C4063 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 0.127f
C4064 mux_8x1_ibr_0.mux_2x1_ibr_0.I1 mux_8x1_ibr_0.mux_2x1_ibr_0.I0 2.74e-20
C4065 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN 0.316f
C4066 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 5.55e-19
C4067 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.00212f
C4068 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_1.IN2 0.36f
C4069 VDD90 a_29053_5018# 0.00123f
C4070 CLK_div_96_mag_0.JK_FF_mag_2.QB a_26368_n2996# 0.00696f
C4071 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 1.83f
C4072 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 0.00101f
C4073 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.00335f
C4074 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_23589_6159# 4.52e-20
C4075 RST a_47994_n18696# 1.23e-20
C4076 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB a_28016_n8779# 0.00392f
C4077 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 1.76f
C4078 VDD93 a_28580_n8735# 3.14e-19
C4079 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 0.00114f
C4080 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 6.82e-19
C4081 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 0.0512f
C4082 F1 a_37168_6821# 0.00731f
C4083 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 1.6e-19
C4084 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 a_36202_6265# 0.00216f
C4085 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00183f
C4086 a_44407_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.46e-19
C4087 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 m3_20882_n11188# 8.64e-19
C4088 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 6.62e-20
C4089 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 0.00975f
C4090 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0443f
C4091 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_48888_n15585# 0.00118f
C4092 a_42083_n15712# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 0.132f
C4093 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 0.0646f
C4094 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0899f
C4095 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.362f
C4096 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT a_50923_n10161# 9.1e-19
C4097 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 2.81e-20
C4098 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.338f
C4099 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_43947_n9019# 2.96e-19
C4100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_44734_2768# 0.0733f
C4101 VDD96 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.651f
C4102 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 8.16e-20
C4103 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.00183f
C4104 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.321f
C4105 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 3.61e-20
C4106 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.121f
C4107 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 3.83f
C4108 CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C4109 VDD93 a_21995_n7106# 3.14e-19
C4110 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 F2 6.25e-19
C4111 CLK dec3x8_ibr_mag_0.and_3_ibr_5.nand3_mag_ibr_0.OUT 0.00254f
C4112 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_43993_n13477# 0.00589f
C4113 VDD108 a_55101_n6818# 3.48e-19
C4114 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0698f
C4115 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.0867f
C4116 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 a_51487_n10161# 1.46e-19
C4117 CLK CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0033f
C4118 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 2.54e-20
C4119 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0343f
C4120 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT 0.00243f
C4121 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 0.0018f
C4122 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0894f
C4123 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_26790_n9831# 0.00372f
C4124 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 2.06e-19
C4125 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 7.08e-20
C4126 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 0.28f
C4127 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.JK_FF_mag_3.QB 1.98f
C4128 CLK_div_96_mag_0.JK_FF_mag_5.QB a_23552_n1789# 2.12e-20
C4129 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00183f
C4130 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 1.17e-19
C4131 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.349f
C4132 VDD93 a_32750_n7675# 0.165f
C4133 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 8.16e-20
C4134 CLK_div_100_mag_0.CLK_div_10_mag_1.CLK a_54663_1671# 0.0101f
C4135 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 a_27170_6159# 0.00372f
C4136 RST a_27334_n16588# 0.00161f
C4137 VDD mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I1 0.422f
C4138 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.107f
C4139 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 3.45e-19
C4140 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 0.0205f
C4141 RST a_53973_n6862# 0.00154f
C4142 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.652f
C4143 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 a_22551_n14504# 0.00369f
C4144 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 0.0775f
C4145 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 1.74e-19
C4146 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 a_50151_n2243# 0.00166f
C4147 RST a_51764_10154# 0.00186f
C4148 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN 0.519f
C4149 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_31291_n17626# 0.00696f
C4150 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_47374_n10160# 0.0733f
C4151 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_53732_n2243# 0.0203f
C4152 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_45541_n18696# 0.069f
C4153 VDD105 a_47453_9057# 3.14e-19
C4154 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.0543f
C4155 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 a_23594_n8743# 0.069f
C4156 a_26814_1919# a_26974_1919# 0.0504f
C4157 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_53375_1671# 0.069f
C4158 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_22839_10099# 0.069f
C4159 RST a_26042_6159# 1.37e-19
C4160 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 9.83e-19
C4161 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_50281_n17599# 0.00119f
C4162 VDD105 a_48380_6284# 3.14e-19
C4163 CLK CLK_div_108_new_mag_0.JK_FF_mag_1.QB 9.53e-20
C4164 VDD105 a_50263_5143# 0.00891f
C4165 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.398f
C4166 RST a_49640_2768# 9.66e-19
C4167 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_46964_n9019# 0.011f
C4168 CLK_div_96_mag_0.JK_FF_mag_0.Q a_25644_n2996# 0.00185f
C4169 VDD105 CLK 1.41f
C4170 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_24512_n18723# 0.0059f
C4171 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.121f
C4172 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 4.23e-20
C4173 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 a_37955_n9984# 0.0157f
C4174 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 0.653f
C4175 a_54509_2768# a_54669_2768# 0.0504f
C4176 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.122f
C4177 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 0.0579f
C4178 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 a_26253_n743# 0.0101f
C4179 VDD93 a_25625_n6010# 2.21e-19
C4180 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_23142_n2930# 8.64e-19
C4181 RST a_45899_7960# 4.48e-19
C4182 VDD96 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_0.OUT 0.762f
C4183 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 0.00114f
C4184 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_50903_n5# 0.069f
C4185 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.00359f
C4186 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.0622f
C4187 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 2.86e-19
C4188 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.343f
C4189 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.458f
C4190 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 a_26250_1919# 1.43e-19
C4191 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 a_31571_n16632# 0.00335f
C4192 VDD108 a_54504_n10161# 0.00888f
C4193 CLK_div_108_new_mag_0.JK_FF_mag_1.Q CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 3.37e-19
C4194 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_47030_n16726# 1.17e-20
C4195 RST a_48534_5187# 9.41e-19
C4196 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 0.0998f
C4197 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0718f
C4198 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_29778_11196# 0.0203f
C4199 RST CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 0.337f
C4200 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00118f
C4201 VDD100 a_50204_2768# 0.00152f
C4202 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.303f
C4203 Vdiv108 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 0.0349f
C4204 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.16f
C4205 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0905f
C4206 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK a_53309_n15631# 2.7e-19
C4207 RST a_27144_10099# 6.26e-19
C4208 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN m3_20882_n11188# 0.00272f
C4209 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK a_53463_n16728# 0.00194f
C4210 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 a_53370_n9020# 0.069f
C4211 CLK_div_90_mag_0.CLK_div_10_mag_0.CLK CLK_div_90_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 1e-19
C4212 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 1.33e-20
C4213 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 a_24491_n7107# 5.1e-19
C4214 VDD110 a_52139_n18696# 3.56e-19
C4215 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K a_50923_n10161# 0.00695f
C4216 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_2.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 2.82e-21
C4217 RST a_53780_n10161# 0.00228f
C4218 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT a_51034_9057# 0.00378f
C4219 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 2.89e-19
C4220 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_51486_1671# 9.32e-19
C4221 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_51393_n6821# 0.069f
C4222 Vdiv110 a_36310_880# 0.00391f
C4223 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 a_47134_n2243# 0.00166f
C4224 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_54597_n15587# 4.52e-20
C4225 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0983f
C4226 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_54751_n16684# 0.00378f
C4227 a_30209_7256# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 1.29e-22
C4228 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0384f
C4229 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.00586f
C4230 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 2.46e-20
C4231 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.998f
C4232 F1 a_37999_280# 2.62e-19
C4233 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 0.783f
C4234 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.391f
C4235 VDD105 VDD110 0.0518f
C4236 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 a_42529_n14305# 1.78e-20
C4237 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 a_32230_5018# 0.0101f
C4238 CLK_div_105_mag_0.CLK_div_10_mag_1.CLK a_54621_10154# 0.00164f
C4239 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.447f
C4240 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 3.48e-19
C4241 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.92f
C4242 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_26932_n2952# 0.00378f
C4243 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.16f
C4244 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 0.977f
C4245 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_39126_n8931# 1.41e-20
C4246 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 Vdiv110 0.0011f
C4247 CLK_div_90_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 a_33204_6159# 2.1e-20
C4248 CLK_div_90_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00943f
C4249 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT a_29341_n16634# 2.88e-20
C4250 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 0.00935f
C4251 VDD90 a_37328_6821# 5.38e-20
C4252 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 a_49098_5187# 0.00372f
C4253 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT 0.0881f
C4254 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN 0.517f
C4255 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT a_51028_n16724# 2.88e-20
C4256 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_44517_n10160# 0.0203f
C4257 Vdiv100 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 0.139f
C4258 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB 0.198f
C4259 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.338f
C4260 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00137f
C4261 Vdiv108 a_53732_n2243# 6.67e-19
C4262 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 4.61f
C4263 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.121f
C4264 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 4.42e-19
C4265 CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 a_29087_8532# 8.64e-19
C4266 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_47030_n16726# 5.83e-19
C4267 CLK_div_108_new_mag_0.JK_FF_mag_1.Q CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.421f
C4268 RST a_45343_n16680# 0.00184f
C4269 CLK CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.298f
C4270 a_44247_n17599# a_44407_n17599# 0.0504f
C4271 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.0063f
C4272 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00166f
C4273 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 0.0655f
C4274 RST a_47134_n2243# 0.00186f
C4275 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_43947_n9019# 0.011f
C4276 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB a_33334_n18723# 0.0112f
C4277 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 0.124f
C4278 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 0.00129f
C4279 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 1f
C4280 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 5.7e-20
C4281 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 a_47914_n16726# 8.64e-19
C4282 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.0635f
C4283 a_51165_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.00696f
C4284 dec3x8_ibr_mag_0.and_3_ibr_5.IN3 a_36042_6821# 0.0079f
C4285 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 a_25055_n7107# 6.14e-21
C4286 a_50111_n5768# CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 1.98e-21
C4287 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00302f
C4288 CLK a_30336_10099# 0.00939f
C4289 Vdiv108 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C4290 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.00125f
C4291 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 a_29862_n9832# 0.00372f
C4292 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00169f
C4293 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 4.02e-20
C4294 a_30244_398# CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 4.52e-20
C4295 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 a_26206_n16632# 0.0101f
C4296 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 2.41f
C4297 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 3.81e-19
C4298 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT 0.00335f
C4299 a_53945_2768# Vdiv110 5.84e-19
C4300 Vdiv96 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 7.46e-19
C4301 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.235f
C4302 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_45969_n2199# 0.0811f
C4303 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 a_29623_6159# 0.069f
C4304 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.121f
C4305 CLK a_32070_5018# 5.65e-19
C4306 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN a_30915_n13291# 0.069f
C4307 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.783f
C4308 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K a_29751_n15493# 3.47e-19
C4309 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT 0.121f
C4310 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB 0.0378f
C4311 a_49789_n9020# CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 4.52e-20
C4312 CLK a_31129_n6271# 0.00479f
C4313 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB a_47863_10154# 0.00696f
C4314 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_44625_n15583# 0.0195f
C4315 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT m3_20882_n11188# 0.00268f
C4316 CLK CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 0.00354f
C4317 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 3.86e-20
C4318 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_28737_n2996# 1.46e-19
C4319 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_45969_n2199# 0.00372f
C4320 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 6.7e-19
C4321 VDD100 a_47698_n2243# 0.00123f
C4322 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 1.33e-20
C4323 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_22466_n8743# 0.0697f
C4324 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.00206f
C4325 a_43793_n10116# m3_20882_n11188# 4.4e-19
C4326 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 a_50353_n9020# 0.069f
C4327 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 0.00975f
C4328 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.24f
C4329 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB 6.38e-19
C4330 CLK_div_96_mag_0.JK_FF_mag_5.QB a_23703_n287# 0.00392f
C4331 F1 Vdiv96 0.0231f
C4332 RST CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.761f
C4333 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.0205f
C4334 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_36827_n10028# 0.00696f
C4335 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 0.515f
C4336 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 a_28623_n15537# 2.79e-20
C4337 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 m3_20882_n11188# 0.0204f
C4338 a_50763_n10161# a_50923_n10161# 0.0504f
C4339 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.0758f
C4340 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 9.55e-20
C4341 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_42529_n14305# 0.0205f
C4342 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 0.407f
C4343 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 8.59e-20
C4344 F1 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.342f
C4345 VDD90 a_28489_5018# 0.00891f
C4346 CLK_div_96_mag_0.JK_FF_mag_2.QB a_26208_n2996# 0.00695f
C4347 CLK CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 5.57e-19
C4348 a_48466_n6273# CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 4.94e-20
C4349 CLK_div_108_new_mag_0.JK_FF_mag_0.QB a_54947_n5721# 0.0114f
C4350 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.019f
C4351 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_23025_6159# 0.0202f
C4352 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 0.0445f
C4353 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 0.116f
C4354 CLK CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 0.0132f
C4355 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 a_36042_6265# 0.00284f
C4356 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.359f
C4357 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0349f
C4358 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 a_28267_n7033# 2.95e-21
C4359 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 1.93f
C4360 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_48324_n15585# 0.011f
C4361 F1 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 0.0863f
C4362 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 3.49e-19
C4363 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 3.97e-19
C4364 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT a_50763_n10161# 2.88e-20
C4365 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_46774_n6273# 1.41e-20
C4366 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_43383_n9019# 0.012f
C4367 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_44170_2768# 0.00378f
C4368 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 0.106f
C4369 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 8.64e-20
C4370 VDD96 CLK 1.89f
C4371 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 9.24e-20
C4372 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN 0.00872f
C4373 VDD93 a_21431_n7106# 3.56e-19
C4374 CLK CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 1.46e-19
C4375 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 3.8e-20
C4376 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 5.85e-19
C4377 VDD108 a_54537_n6818# 3.14e-19
C4378 CLK a_51193_n19793# 2.22e-19
C4379 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 a_44475_n5176# 0.0101f
C4380 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_26226_n9831# 0.069f
C4381 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_26349_n6010# 1.17e-20
C4382 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 0.188f
C4383 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 2.25e-21
C4384 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN 0.0836f
C4385 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 7.34e-20
C4386 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 4.27e-20
C4387 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 4.07e-19
C4388 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_32865_n15491# 4.52e-20
C4389 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_41124_n16098# 0.0111f
C4390 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.121f
C4391 a_47430_n18696# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.0732f
C4392 CLK_div_100_mag_0.CLK_div_10_mag_1.CLK a_54503_1671# 0.00939f
C4393 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C4394 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 a_26606_6159# 0.069f
C4395 RST a_26770_n16588# 0.00192f
C4396 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K a_54658_n9064# 8.64e-19
C4397 a_38966_n8931# a_39126_n8931# 0.0504f
C4398 RST a_53813_n6862# 0.00177f
C4399 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 0.048f
C4400 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 a_25055_n7107# 0.069f
C4401 RST a_51604_10154# 0.00186f
C4402 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 a_49991_n2243# 0.00119f
C4403 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_40972_n9984# 0.0811f
C4404 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_30727_n17626# 0.00964f
C4405 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 1.17e-19
C4406 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_53168_n2243# 1.5e-20
C4407 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_46810_n10116# 0.00378f
C4408 VDD105 a_46889_9057# 3.56e-19
C4409 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 a_29053_5018# 3.6e-22
C4410 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 a_23030_n8743# 1.46e-21
C4411 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 1.98e-19
C4412 RST a_27342_n1855# 0.0019f
C4413 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_52811_1671# 0.00372f
C4414 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.00335f
C4415 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_22275_10099# 0.00372f
C4416 RST a_25478_6115# 7.09e-19
C4417 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT 9.52e-19
C4418 VDD105 a_47816_6284# 3.14e-19
C4419 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB 0.0838f
C4420 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.359f
C4421 a_43963_n1146# a_44123_n1146# 0.0504f
C4422 RST CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.00667f
C4423 VDD105 a_50103_5143# 0.0132f
C4424 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 4.95e-20
C4425 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 0.359f
C4426 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 5.63e-21
C4427 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0228f
C4428 CLK_div_96_mag_0.JK_FF_mag_0.Q a_25484_n2996# 0.00143f
C4429 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 8.59e-20
C4430 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_46400_n9019# 0.00118f
C4431 VDD99 a_27334_n16588# 3.14e-19
C4432 CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0345f
C4433 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 a_37391_n9984# 0.00859f
C4434 CLK_div_108_new_mag_0.JK_FF_mag_1.Q a_53819_n5721# 6.43e-21
C4435 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 7.35e-19
C4436 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 0.00641f
C4437 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT m3_20882_n11188# 4.97e-19
C4438 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.28f
C4439 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 0.0655f
C4440 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 a_26093_n743# 0.0102f
C4441 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 0.124f
C4442 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 2.01e-19
C4443 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 6.69e-19
C4444 VDD90 dec3x8_ibr_mag_0.and_3_ibr_0.nand3_mag_ibr_0.OUT 0.148f
C4445 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_45039_n5176# 0.0036f
C4446 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 0.166f
C4447 CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_90_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 3.34e-19
C4448 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.768f
C4449 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 a_25686_1919# 0.011f
C4450 VDD110 a_51193_n19793# 6e-19
C4451 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 a_28828_1497# 7.48e-20
C4452 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.179f
C4453 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 5.32e-19
C4454 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 8.26e-20
C4455 RST a_45927_6284# 0.00104f
C4456 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 0.0022f
C4457 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0218f
C4458 VDD108 a_53940_n10161# 0.0012f
C4459 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 3.27e-20
C4460 CLK_div_96_mag_0.JK_FF_mag_5.QB CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00999f
C4461 VDD Vdiv100 0.738f
C4462 RST CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.00543f
C4463 a_29801_1733# CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.132f
C4464 RST a_47970_5143# 0.00186f
C4465 Vdiv100 a_43719_n120# 0.0157f
C4466 CLK_div_96_mag_0.JK_FF_mag_2.Q CLK_div_96_mag_0.JK_FF_mag_3.QB 0.307f
C4467 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_29618_11196# 0.0733f
C4468 VDD100 a_49640_2768# 0.00152f
C4469 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_52161_n19793# 0.0084f
C4470 Vdiv108 a_36873_280# 0.00307f
C4471 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0432f
C4472 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 4.42e-19
C4473 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 0.122f
C4474 RST a_26984_10099# 5.13e-19
C4475 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK a_53303_n16728# 0.00194f
C4476 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.911f
C4477 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 a_52806_n9020# 0.00372f
C4478 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.118f
C4479 VDD110 a_51575_n18696# 3.14e-19
C4480 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K a_50763_n10161# 0.00696f
C4481 RST a_53216_n10117# 0.00164f
C4482 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 0.00203f
C4483 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_50922_1671# 3.12e-19
C4484 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.00237f
C4485 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 a_46974_n2243# 0.001f
C4486 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_54033_n15587# 0.0195f
C4487 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 0.122f
C4488 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00157f
C4489 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_54187_n16728# 0.0733f
C4490 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00118f
C4491 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 5.73e-20
C4492 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 a_26036_5018# 3.6e-22
C4493 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 5.51e-20
C4494 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00265f
C4495 VDD90 a_27150_11196# 0.0132f
C4496 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 a_32070_5018# 0.0102f
C4497 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.28f
C4498 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN 0.0405f
C4499 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 5.32e-19
C4500 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_26368_n2996# 0.0733f
C4501 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0385f
C4502 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_26817_n699# 0.0036f
C4503 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_38966_n8931# 1.86e-20
C4504 a_30435_n1855# CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 4.52e-20
C4505 VDD96 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.391f
C4506 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT a_29181_n16634# 9.1e-19
C4507 VDD90 a_37168_6821# 8.75e-20
C4508 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT a_50868_n16724# 9.1e-19
C4509 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 a_48534_5187# 0.069f
C4510 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.0725f
C4511 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_44357_n10160# 0.0733f
C4512 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 a_40254_n8887# 4.9e-20
C4513 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 0.126f
C4514 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.0477f
C4515 a_29241_7256# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 3.38e-20
C4516 Vdiv108 a_53168_n2243# 0.00158f
C4517 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0718f
C4518 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_44061_n15627# 3.43e-19
C4519 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.159f
C4520 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.27f
C4521 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_45907_n16680# 0.0157f
C4522 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 1.96f
C4523 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 a_33744_n17626# 2.58e-20
C4524 CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 7.37e-20
C4525 RST a_44779_n16724# 0.00349f
C4526 RST a_46974_n2243# 0.00186f
C4527 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_43383_n9019# 0.00118f
C4528 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 0.69f
C4529 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 3.09e-19
C4530 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 9.58e-19
C4531 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 a_23510_n15620# 3.17e-19
C4532 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 0.026f
C4533 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 a_51652_2768# 0.001f
C4534 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 a_53216_n10117# 0.0036f
C4535 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 a_24491_n7107# 0.069f
C4536 a_51005_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.00695f
C4537 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_51729_n17599# 0.00378f
C4538 VDD dec3x8_ibr_mag_0.and_3_ibr_3.nand3_mag_ibr_0.OUT 0.719f
C4539 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.0432f
C4540 CLK a_29772_10099# 6.43e-21
C4541 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_34462_n18723# 0.0697f
C4542 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 0.0655f
C4543 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 a_29298_n9832# 0.069f
C4544 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_43831_7266# 9.21e-20
C4545 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.338f
C4546 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 1.57f
C4547 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_21902_n8787# 3.87e-20
C4548 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 a_26046_n16632# 0.0102f
C4549 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.391f
C4550 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00117f
C4551 a_53785_2768# Vdiv110 5.84e-19
C4552 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 1.53e-20
C4553 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_45405_n2199# 0.00964f
C4554 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0836f
C4555 a_36667_n10028# a_36827_n10028# 0.0504f
C4556 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN 0.423f
C4557 CLK a_31506_5018# 0.00134f
C4558 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN a_30210_n13332# 4.43e-21
C4559 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.303f
C4560 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_0.QB 0.00999f
C4561 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 1.17e-19
C4562 CLK a_30165_n6282# 7.37e-19
C4563 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB a_47299_10154# 0.00964f
C4564 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 Vdiv108 0.0488f
C4565 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 8.28e-20
C4566 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0358f
C4567 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB a_26790_n9831# 0.0811f
C4568 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00118f
C4569 CLK_div_96_mag_0.JK_FF_mag_4.Q a_25375_354# 7.32e-19
C4570 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB 0.0615f
C4571 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_45405_n2199# 0.069f
C4572 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.394f
C4573 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_0.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00132f
C4574 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.00113f
C4575 VDD110 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 0.125f
C4576 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK a_44977_n18696# 6.43e-21
C4577 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_24901_n6010# 0.0036f
C4578 CLK_div_105_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 a_55179_7683# 2.44e-20
C4579 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 4.24e-20
C4580 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 0.124f
C4581 Vdiv99 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN 0.0038f
C4582 VDD100 a_47134_n2243# 0.00863f
C4583 VDD96 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 0.31f
C4584 a_43229_n10116# m3_20882_n11188# 4.57e-19
C4585 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 a_49789_n9020# 0.00372f
C4586 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.36f
C4587 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00163f
C4588 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00617f
C4589 a_44846_10154# a_45006_10154# 0.0504f
C4590 CLK_div_96_mag_0.JK_FF_mag_5.QB a_23139_n287# 2.25e-19
C4591 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 1.71e-21
C4592 RST CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.477f
C4593 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_36667_n10028# 0.00695f
C4594 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_3_mag_0.CLK 1e-20
C4595 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 2.57f
C4596 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00122f
C4597 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0854f
C4598 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_0.OUT 0.0622f
C4599 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_51285_n1102# 4.52e-20
C4600 F1 Vdiv108 0.106f
C4601 CLK CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.00156f
C4602 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 2.51e-19
C4603 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 8.58e-20
C4604 CLK_div_105_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT 0.11f
C4605 VDD90 a_28329_5018# 0.0132f
C4606 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT 0.131f
C4607 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.653f
C4608 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 0.431f
C4609 a_45564_9057# a_45724_9057# 0.0504f
C4610 CLK_div_108_new_mag_0.JK_FF_mag_0.QB a_54383_n5721# 2.96e-19
C4611 VDD93 a_27856_n8779# 0.00554f
C4612 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 4.84e-19
C4613 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.122f
C4614 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 8.16e-20
C4615 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 0.175f
C4616 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 a_27324_5062# 0.00372f
C4617 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 1.35e-20
C4618 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB a_46867_7960# 1.45e-20
C4619 F0 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT 0.00112f
C4620 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_47760_n15585# 1.43e-19
C4621 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.875f
C4622 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_45452_1671# 0.00119f
C4623 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.00488f
C4624 RST CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0244f
C4625 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 0.00591f
C4626 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB 0.28f
C4627 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.00822f
C4628 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_46614_n6273# 1.86e-20
C4629 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.JK_FF_mag_0.Q 0.00927f
C4630 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT a_54866_n1102# 1.54e-19
C4631 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 2.57e-20
C4632 Vdiv110 a_55067_297# 0.00125f
C4633 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 CLK_div_105_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00311f
C4634 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.395f
C4635 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 1.98e-19
C4636 CLK CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 0.00345f
C4637 Vdiv96 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 4.46e-19
C4638 CLK_div_96_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 3.34e-19
C4639 RST CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.0042f
C4640 CLK a_31733_n19822# 0.0105f
C4641 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_108_new_mag_0.JK_FF_mag_1.Q 3.16e-21
C4642 Vdiv99 a_36310_n1822# 0.00347f
C4643 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 a_44315_n5176# 0.0102f
C4644 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 a_51492_2768# 1.46e-19
C4645 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 0.339f
C4646 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 9.75e-21
C4647 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 1.53e-19
C4648 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.267f
C4649 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_26189_n6010# 1.5e-20
C4650 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_32301_n15491# 0.0195f
C4651 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_23594_n8743# 0.00118f
C4652 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.28f
C4653 CLK_div_100_mag_0.CLK_div_10_mag_1.CLK a_53939_1671# 6.43e-21
C4654 a_47270_n18696# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.0203f
C4655 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.857f
C4656 RST a_26206_n16632# 0.00341f
C4657 VDD99 Vdiv90 0.114f
C4658 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 0.0703f
C4659 CLK_div_96_mag_0.JK_FF_mag_5.Q CLK_div_96_mag_0.JK_FF_mag_0.Q 0.149f
C4660 RST a_53249_n6862# 0.00251f
C4661 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.00213f
C4662 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 2.21e-19
C4663 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 a_24491_n7107# 0.00372f
C4664 RST a_51040_10154# 0.00169f
C4665 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 a_48986_n2199# 0.0157f
C4666 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_40408_n9984# 0.00964f
C4667 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_30163_n17626# 0.0811f
C4668 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_2.OUT CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT 0.121f
C4669 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_4.QB 0.0387f
C4670 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 8.31e-21
C4671 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN 0.431f
C4672 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_53008_n2243# 1.17e-20
C4673 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C4674 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.397f
C4675 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN 0.00527f
C4676 VDD93 a_37328_6821# 7.02e-19
C4677 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0707f
C4678 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 a_28489_5018# 0.00166f
C4679 RST a_26778_n1855# 0.00101f
C4680 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 9.52e-19
C4681 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C4682 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.768f
C4683 RST a_25318_6115# 0.00109f
C4684 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.00101f
C4685 Vdiv99 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN 0.00397f
C4686 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.0063f
C4687 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.36f
C4688 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 2.19e-20
C4689 VDD105 a_47252_6240# 2.66e-19
C4690 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 0.651f
C4691 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_36178_n16592# 0.00378f
C4692 a_37328_6821# F0 3.14e-19
C4693 VDD105 a_49098_5187# 0.00152f
C4694 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.182f
C4695 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_48466_n6273# 0.012f
C4696 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 4.3e-20
C4697 CLK_div_96_mag_0.JK_FF_mag_0.Q a_24270_n2886# 0.0157f
C4698 VDD99 a_26770_n16588# 3.14e-19
C4699 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT 3.84e-20
C4700 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.IN2 Vdiv99 4.51e-19
C4701 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 a_36827_n10028# 0.0101f
C4702 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 4.25e-20
C4703 a_54498_n9064# a_54658_n9064# 0.0504f
C4704 CLK_div_108_new_mag_0.JK_FF_mag_1.Q a_53255_n5765# 0.00939f
C4705 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_48268_n1102# 4.52e-20
C4706 CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 1.61e-19
C4707 CLK_div_108_new_mag_0.JK_FF_mag_0.QB CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.28f
C4708 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 3.98e-19
C4709 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.0378f
C4710 a_50669_n6865# a_50829_n6865# 0.0504f
C4711 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.0725f
C4712 a_42529_n14305# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN 0.069f
C4713 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_51803_n5724# 0.00118f
C4714 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 4.68e-20
C4715 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 a_25529_n743# 0.00789f
C4716 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 a_53850_6284# 6.43e-21
C4717 VDD93 a_24901_n6010# 3.14e-19
C4718 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.00101f
C4719 RST CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 0.0072f
C4720 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 5.32f
C4721 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.655f
C4722 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 0.198f
C4723 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.055f
C4724 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_44894_2768# 0.00695f
C4725 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 3.86e-20
C4726 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.402f
C4727 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.288f
C4728 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 a_25122_1919# 0.00118f
C4729 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 1.47e-20
C4730 VDD108 a_53780_n10161# 9.82e-19
C4731 RST a_45363_6284# 0.00167f
C4732 CLK CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 0.00542f
C4733 RST a_47810_5143# 0.00169f
C4734 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 1.94f
C4735 CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.IN2 a_51205_n7921# 7.48e-20
C4736 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN 2.86e-19
C4737 Vdiv100 a_43559_n120# 0.203f
C4738 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_29054_11196# 0.00378f
C4739 a_53249_n6862# CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 1.8e-21
C4740 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 0.653f
C4741 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 0.286f
C4742 a_22301_6115# a_22461_6115# 0.0504f
C4743 RST a_26420_10099# 1.8e-19
C4744 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0843f
C4745 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT 0.0763f
C4746 VDD110 a_51011_n18696# 3.14e-19
C4747 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.998f
C4748 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K a_50199_n10117# 0.00964f
C4749 RST a_52652_n10117# 0.00114f
C4750 VDD dec3x8_ibr_mag_0.and_3_ibr_6.IN3 1.05f
C4751 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.0151f
C4752 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K a_31352_6115# 8.64e-19
C4753 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_26420_10099# 0.0697f
C4754 a_48623_n13424# a_48783_n13424# 0.0504f
C4755 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 3.59f
C4756 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_50358_1671# 7.4e-19
C4757 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.122f
C4758 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 a_29213_n7028# 3.11e-21
C4759 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0143f
C4760 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0569f
C4761 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 a_45969_n2199# 0.0157f
C4762 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_53892_n2243# 8.64e-19
C4763 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.00125f
C4764 CLK_div_108_new_mag_0.JK_FF_mag_1.Q CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.235f
C4765 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_28495_6115# 1.41e-20
C4766 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_54027_n16728# 0.0203f
C4767 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.647f
C4768 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB 2.59e-21
C4769 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 a_25472_5018# 0.00166f
C4770 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.0615f
C4771 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_25702_11196# 0.069f
C4772 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.00178f
C4773 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT 0.053f
C4774 VDD90 a_26990_11196# 0.00888f
C4775 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 a_31506_5018# 0.00789f
C4776 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 0.0512f
C4777 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.92f
C4778 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_26208_n2996# 0.0203f
C4779 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 0.359f
C4780 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.28f
C4781 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 0.0709f
C4782 VDD99 dec3x8_ibr_mag_0.and_3_ibr_4.nand3_mag_ibr_0.OUT 8.47e-19
C4783 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 0.58f
C4784 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_47528_n9019# 0.0697f
C4785 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT a_28617_n16634# 0.0731f
C4786 a_45452_1671# a_45612_1671# 0.0504f
C4787 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00178f
C4788 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT a_50304_n16724# 0.0731f
C4789 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_49122_n18696# 9.26e-19
C4790 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_43793_n10116# 0.00378f
C4791 VDD93 a_40972_n9984# 3.14e-19
C4792 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.22f
C4793 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 9.52e-19
C4794 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K a_52839_n5# 0.0027f
C4795 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00166f
C4796 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 4.75f
C4797 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 0.434f
C4798 RST CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00941f
C4799 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0042f
C4800 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT Vdiv110 0.00764f
C4801 Vdiv108 a_53008_n2243# 0.00158f
C4802 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 0.00212f
C4803 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_43901_n15627# 4.47e-19
C4804 CLK_div_100_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_100_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.11f
C4805 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 0.39f
C4806 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.175f
C4807 a_32009_n18723# a_32169_n18723# 0.0504f
C4808 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_45343_n16680# 0.00859f
C4809 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 0.582f
C4810 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 1.17e-19
C4811 RST a_44619_n16724# 0.00207f
C4812 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 6.63e-19
C4813 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 5.98e-20
C4814 RST a_45969_n2199# 9.66e-19
C4815 RST CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0592f
C4816 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.00116f
C4817 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 a_51492_2768# 0.00166f
C4818 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I1 Vdiv100 0.00184f
C4819 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0334f
C4820 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.651f
C4821 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_33898_n18723# 0.0059f
C4822 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_43671_7266# 3.02e-19
C4823 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 a_25482_n16632# 0.0152f
C4824 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.311f
C4825 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.122f
C4826 a_53221_2768# Vdiv110 6.25e-19
C4827 CLK_div_105_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 1.29e-19
C4828 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 6.86e-20
C4829 F1 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 0.00158f
C4830 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 0.447f
C4831 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_44841_n2243# 0.00696f
C4832 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN a_30050_n13332# 3.44e-21
C4833 CLK a_31346_5018# 0.00134f
C4834 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 0.0042f
C4835 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB a_46735_10154# 0.0811f
C4836 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_51397_6284# 4.52e-20
C4837 a_35747_280# Vdiv108 1.13e-20
C4838 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_1.IN2 CLK_div_96_mag_0.JK_FF_mag_0.QB 1.38e-19
C4839 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT 0.768f
C4840 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 0.00118f
C4841 RST CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.0627f
C4842 CLK_div_108_new_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_47528_n9019# 5.01e-20
C4843 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_45343_n16680# 0.00378f
C4844 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB a_26226_n9831# 0.00964f
C4845 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 0.0871f
C4846 VDD90 a_30502_11196# 0.00743f
C4847 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 8.23e-19
C4848 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 m3_20882_n11188# 7.8e-19
C4849 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 0.00115f
C4850 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 0.0151f
C4851 CLK_div_105_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 a_55019_7683# 9.02e-19
C4852 VDD100 a_46974_n2243# 0.0123f
C4853 Vdiv99 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 0.00112f
C4854 CLK CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 4.05e-20
C4855 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 a_44799_n7920# 7.48e-20
C4856 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0592f
C4857 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 0.0844f
C4858 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 5.74e-20
C4859 a_40972_n9984# m3_20882_n11188# 3.71e-19
C4860 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 a_30210_n13332# 0.0121f
C4861 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00531f
C4862 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT 0.00134f
C4863 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT 0.0763f
C4864 CLK_div_96_mag_0.JK_FF_mag_5.QB a_22575_n287# 2.96e-19
C4865 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.745f
C4866 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 8.16e-20
C4867 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_50721_n1102# 0.0202f
C4868 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB 0.198f
C4869 a_44324_1671# Vdiv110 9.95e-20
C4870 Vdiv90 F2 0.00314f
C4871 VDD90 a_27324_5062# 0.00152f
C4872 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.233f
C4873 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 0.777f
C4874 VDD93 a_31128_n7028# 5.19e-19
C4875 CLK_div_108_new_mag_0.JK_FF_mag_0.QB a_53819_n5721# 3.33e-19
C4876 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.251f
C4877 VDD93 dec3x8_ibr_mag_0.and_3_ibr_0.nand3_mag_ibr_0.OUT 0.0233f
C4878 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 1.84e-21
C4879 a_51034_9057# CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 7.43e-22
C4880 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 a_26760_5062# 0.069f
C4881 CLK CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT 0.272f
C4882 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 a_38966_n8931# 0.00149f
C4883 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_44511_n9019# 0.0697f
C4884 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_47196_n15629# 0.00119f
C4885 dec3x8_ibr_mag_0.and_3_ibr_0.nand3_mag_ibr_0.OUT F0 1.04e-19
C4886 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_44888_1671# 1.43e-19
C4887 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_48478_n16682# 0.0036f
C4888 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0905f
C4889 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.977f
C4890 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.28f
C4891 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0281f
C4892 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.523f
C4893 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 0.00164f
C4894 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 3.61e-20
C4895 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 4.89e-20
C4896 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_45449_n6273# 0.0112f
C4897 a_51849_n1102# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 4.52e-20
C4898 RST CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.268f
C4899 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.01f
C4900 CLK_div_96_mag_0.JK_FF_mag_2.Q CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 6.64e-19
C4901 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 1.76e-20
C4902 VDD105 a_51764_10154# 0.0123f
C4903 Vdiv110 a_54907_297# 6.62e-19
C4904 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_44687_n1102# 0.00378f
C4905 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 0.343f
C4906 VDD99 dec3x8_ibr_mag_0.and_3_ibr_5.IN3 0.00762f
C4907 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 0.109f
C4908 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 0.109f
C4909 CLK_div_96_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_29801_1733# 3.25e-19
C4910 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 1.99e-20
C4911 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 a_45189_n15583# 0.0059f
C4912 VDD108 a_53813_n6862# 2.21e-19
C4913 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.159f
C4914 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 a_50199_n10117# 0.0036f
C4915 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 1.28e-20
C4916 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 0.651f
C4917 F2 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 0.00519f
C4918 Vdiv99 a_35747_n1822# 5.8e-19
C4919 VDD mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 0.46f
C4920 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 0.029f
C4921 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 a_43751_n5176# 0.00789f
C4922 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_25625_n6010# 0.0203f
C4923 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 a_21896_n9884# 0.00164f
C4924 RST CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.771f
C4925 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.00183f
C4926 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 0.378f
C4927 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_23030_n8743# 0.011f
C4928 a_47270_n18696# a_47430_n18696# 0.0504f
C4929 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 2.45e-22
C4930 RST a_26046_n16632# 0.0024f
C4931 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 1.86e-19
C4932 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.121f
C4933 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.0147f
C4934 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 2.81e-20
C4935 RST a_53089_n6862# 0.00266f
C4936 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 a_28392_354# 0.00149f
C4937 VDD108 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.742f
C4938 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_48380_6284# 4.52e-20
C4939 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_39844_n10028# 0.00696f
C4940 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 a_48422_n2199# 0.00859f
C4941 RST a_50880_10154# 0.00186f
C4942 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.414f
C4943 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB a_23283_n7106# 1.76e-20
C4944 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 1.83e-19
C4945 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C4946 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C4947 CLK_div_100_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00182f
C4948 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_53469_n15631# 1.19e-20
C4949 VDD105 a_45899_7960# 3.14e-19
C4950 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB a_23748_n9840# 0.0811f
C4951 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 8.16e-20
C4952 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_48558_n18696# 0.0059f
C4953 VDD93 a_37168_6821# 0.00123f
C4954 CLK CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.00461f
C4955 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 a_28329_5018# 0.00119f
C4956 RST a_26214_n1855# 3.73e-19
C4957 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 a_21902_n8787# 2.79e-20
C4958 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 a_28823_n17626# 1.38e-20
C4959 Vdiv105 a_43831_7266# 0.0147f
C4960 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.0675f
C4961 RST a_24153_6159# 0.00168f
C4962 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.0275f
C4963 RST CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.194f
C4964 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 7.24e-19
C4965 a_47492_n5176# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0733f
C4966 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.018f
C4967 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_23589_6159# 0.0059f
C4968 VDD105 a_47092_6240# 3.78e-19
C4969 CLK CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 1.05e-19
C4970 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_35614_n16636# 0.0733f
C4971 a_37168_6821# F0 5.62e-19
C4972 VDD105 a_48534_5187# 0.00152f
C4973 RST a_49276_n17599# 0.00122f
C4974 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_47902_n6273# 2.96e-19
C4975 CLK_div_96_mag_0.JK_FF_mag_0.Q a_23706_n2886# 0.00859f
C4976 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 7.38e-19
C4977 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 a_36667_n10028# 0.0102f
C4978 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.0763f
C4979 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_45724_9057# 0.0203f
C4980 CLK_div_108_new_mag_0.JK_FF_mag_1.Q a_53095_n5765# 0.0101f
C4981 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 m3_20882_n11188# 7.51e-19
C4982 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_47704_n1102# 0.0202f
C4983 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 4.26e-19
C4984 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 a_48888_n15585# 0.00372f
C4985 a_43957_n2243# a_44117_n2243# 0.0504f
C4986 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_51239_n5724# 0.011f
C4987 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 a_25369_n743# 0.00335f
C4988 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 a_53286_6240# 0.00939f
C4989 VDD93 a_24337_n6010# 3.15e-19
C4990 F2 dec3x8_ibr_mag_0.and_3_ibr_4.nand3_mag_ibr_0.OUT 2.94e-19
C4991 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.36f
C4992 a_50922_1671# CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 7.43e-22
C4993 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_44734_2768# 0.00696f
C4994 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K a_25328_n15535# 0.00472f
C4995 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 8.93e-21
C4996 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 4.98e-19
C4997 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN a_45251_n1102# 8.17e-21
C4998 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 5.5e-20
C4999 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 8.16e-20
C5000 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.00183f
C5001 RST a_45131_n17599# 0.00283f
C5002 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK a_39402_n7788# 0.0103f
C5003 a_24778_n9875# a_24938_n9875# 0.0504f
C5004 VDD108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 2.86e-19
C5005 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN a_29708_n8735# 3.59e-20
C5006 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 2.71e-21
C5007 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 4.33e-19
C5008 VDD108 a_53216_n10117# 0.00149f
C5009 RST a_44799_6284# 0.0012f
C5010 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_29618_11196# 8.64e-19
C5011 RST a_47246_5143# 0.00186f
C5012 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN a_45787_574# 0.069f
C5013 CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.IN2 a_50232_n7685# 8.64e-19
C5014 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 4.85e-20
C5015 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 7.06e-19
C5016 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 1.36e-19
C5017 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT a_26099_398# 3.53e-20
C5018 RST CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0765f
C5019 VDD Vdiv 2.79f
C5020 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0169f
C5021 RST a_25856_10099# 0.0011f
C5022 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT a_32076_6159# 5.94e-20
C5023 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 0.00147f
C5024 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_29905_n16590# 0.00378f
C5025 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 a_26820_3016# 1.46e-19
C5026 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 0.0497f
C5027 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.VOUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 2.17e-20
C5028 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K a_49635_n10117# 0.0811f
C5029 RST a_51647_n10161# 0.00218f
C5030 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 2.48e-19
C5031 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_25856_10099# 0.0059f
C5032 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00166f
C5033 VDD90 a_22718_8532# 0.165f
C5034 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.IN1 1.64e-19
C5035 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_49794_1671# 7.4e-19
C5036 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 1.07f
C5037 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 2.59e-21
C5038 CLK_div_108_new_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 3.34e-19
C5039 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 a_45405_n2199# 0.00859f
C5040 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 4.54f
C5041 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 6.41e-20
C5042 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_50447_n18696# 2.79e-20
C5043 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_28335_6115# 1.86e-20
C5044 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_53463_n16728# 1.5e-20
C5045 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_37955_n9984# 0.00372f
C5046 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 a_25312_5018# 0.001f
C5047 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 0.00392f
C5048 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 2f
C5049 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_25138_11196# 0.00372f
C5050 VDD90 a_26426_11196# 0.0012f
C5051 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 0.994f
C5052 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 a_31346_5018# 0.00335f
C5053 CLK a_26349_n6010# 0.00544f
C5054 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 a_51015_7381# 2.48e-19
C5055 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.5e-19
C5056 VDD110 a_46259_n17599# 0.00152f
C5057 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_25644_n2996# 1.5e-20
C5058 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_25375_354# 8.64e-19
C5059 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 4.2e-19
C5060 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_54383_n5721# 4.52e-20
C5061 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT a_28457_n16634# 0.0202f
C5062 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_46964_n9019# 0.0059f
C5063 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.233f
C5064 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 0.0246f
C5065 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00158f
C5066 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT 0.748f
C5067 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT a_50144_n16724# 0.0202f
C5068 VDD93 a_40408_n9984# 3.14e-19
C5069 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.321f
C5070 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 1.96f
C5071 Vdiv108 a_52003_n2199# 7.51e-19
C5072 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K 0.0156f
C5073 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 4.28e-19
C5074 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.338f
C5075 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_24116_n1789# 0.00118f
C5076 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_45603_n5176# 0.00372f
C5077 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_44779_n16724# 0.0101f
C5078 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.211f
C5079 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 3.83e-19
C5080 RST a_44055_n16724# 9.47e-19
C5081 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.346f
C5082 RST a_45405_n2199# 9.41e-19
C5083 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_22559_n7106# 0.0697f
C5084 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.00942f
C5085 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_30502_11196# 0.0202f
C5086 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 a_50928_2768# 3.6e-22
C5087 a_47264_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 2.81e-19
C5088 VDD a_36042_6821# 2.09e-19
C5089 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 8.58e-20
C5090 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN 2.91e-19
C5091 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_29778_11196# 0.00695f
C5092 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 a_30336_10099# 2.79e-20
C5093 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.16f
C5094 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.233f
C5095 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C5096 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.125f
C5097 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 a_25322_n16632# 0.0124f
C5098 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.00488f
C5099 CLK_div_96_mag_0.JK_FF_mag_5.Q CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.235f
C5100 a_52657_2768# Vdiv110 6.45e-19
C5101 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 3.09e-19
C5102 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_44681_n2243# 0.00695f
C5103 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 5.62e-19
C5104 CLK a_30341_5062# 6.21e-19
C5105 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.233f
C5106 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.00761f
C5107 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_50833_6284# 0.0202f
C5108 Vdiv93 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.13f
C5109 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 0.00761f
C5110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_44779_n16724# 0.0733f
C5111 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB a_25662_n9875# 0.00696f
C5112 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT m3_20882_n11188# 8.83e-19
C5113 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.391f
C5114 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 CLK_div_90_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00357f
C5115 VDD90 a_30342_11196# 0.00305f
C5116 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 5.45e-20
C5117 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 a_54597_n15587# 0.00605f
C5118 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 0.321f
C5119 F2 dec3x8_ibr_mag_0.and_3_ibr_5.IN3 0.171f
C5120 VDD100 a_45969_n2199# 0.00152f
C5121 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0622f
C5122 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN 0.519f
C5123 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 6.36e-20
C5124 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 0.00314f
C5125 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.28f
C5126 CLK CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 4.7e-19
C5127 a_40408_n9984# m3_20882_n11188# 3.57e-19
C5128 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 0.129f
C5129 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.122f
C5130 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.655f
C5131 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.0515f
C5132 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 a_30050_n13332# 0.00747f
C5133 a_23703_n287# a_23863_n287# 0.0504f
C5134 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 5.37e-19
C5135 CLK_div_96_mag_0.JK_FF_mag_5.QB a_22011_n287# 0.0114f
C5136 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.00169f
C5137 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 0.69f
C5138 F1 dec3x8_ibr_mag_0.and_3_ibr_6.nand3_mag_ibr_0.OUT 0.0252f
C5139 VDD110 a_44413_n18696# 2.66e-19
C5140 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT Vdiv110 0.00562f
C5141 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 1e-19
C5142 CLK_div_90_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 4.42e-19
C5143 CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 9.83e-19
C5144 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 9.24e-20
C5145 a_43760_1671# Vdiv110 9.95e-20
C5146 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 2.57e-20
C5147 Vdiv90 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT 0.00186f
C5148 VDD90 a_26760_5062# 0.00152f
C5149 Vdiv96 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT 9.23e-19
C5150 CLK_div_108_new_mag_0.JK_FF_mag_0.QB a_53255_n5765# 0.00392f
C5151 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 1.76e-20
C5152 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_45541_n18696# 0.0059f
C5153 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 0.209f
C5154 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_44799_6284# 0.00378f
C5155 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C5156 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 0.283f
C5157 RST CLK_div_96_mag_0.JK_FF_mag_5.QB 0.0683f
C5158 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_28663_n17626# 1.46e-19
C5159 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 8.16e-20
C5160 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 0.0635f
C5161 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00118f
C5162 a_26183_n7107# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 3.42e-20
C5163 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 2.92e-20
C5164 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_43947_n9019# 0.0059f
C5165 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 6.36e-19
C5166 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 0.127f
C5167 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.65f
C5168 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_44324_1671# 0.011f
C5169 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 1.36e-19
C5170 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 a_53780_n10161# 8.64e-19
C5171 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 1.48e-19
C5172 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 0.233f
C5173 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00254f
C5174 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 9.75e-19
C5175 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_22466_n8743# 5e-20
C5176 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_47902_n6273# 0.0059f
C5177 VDD105 a_51604_10154# 0.00863f
C5178 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_44123_n1146# 0.0732f
C5179 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB 0.311f
C5180 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.0915f
C5181 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00156f
C5182 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 2.81e-20
C5183 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.00668f
C5184 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN m3_20882_n11188# 0.00101f
C5185 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB 0.103f
C5186 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 a_44625_n15583# 0.0697f
C5187 a_32295_n16632# a_32455_n16632# 0.0504f
C5188 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.457f
C5189 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 0.359f
C5190 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.103f
C5191 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 m3_20882_n11188# 8.31e-19
C5192 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN a_41124_n16098# 0.069f
C5193 CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 4.44e-20
C5194 CLK_div_108_new_mag_0.JK_FF_mag_1.QB CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C5195 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 9.71e-20
C5196 VDD93 Vdiv96 0.122f
C5197 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_30187_6159# 0.0114f
C5198 Vdiv99 a_35184_n1822# 7.81e-19
C5199 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 0.629f
C5200 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.101f
C5201 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 a_43591_n5176# 0.00335f
C5202 dec3x8_ibr_mag_0.and_3_ibr_4.nand3_mag_ibr_0.OUT dec3x8_ibr_mag_0.and_3_ibr_5.nand3_mag_ibr_0.OUT 6.66e-19
C5203 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT 0.25f
C5204 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.122f
C5205 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_25465_n6010# 0.0733f
C5206 RST CLK_div_96_mag_0.JK_FF_mag_3.Q 0.242f
C5207 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 1.48e-19
C5208 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 a_21736_n9884# 0.00117f
C5209 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 0.321f
C5210 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I1 0.109f
C5211 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 2.08e-19
C5212 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_22466_n8743# 1.43e-19
C5213 a_22275_10099# CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 4.94e-20
C5214 CLK_div_108_new_mag_0.JK_FF_mag_0.QB CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.103f
C5215 RST CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 0.0507f
C5216 RST a_25482_n16632# 0.00139f
C5217 F0 Vdiv96 0.128f
C5218 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.JK_FF_mag_4.QB 1.96f
C5219 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.00656f
C5220 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 0.109f
C5221 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_39690_n8887# 0.00378f
C5222 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 a_47453_9057# 6.06e-21
C5223 RST a_51957_n6821# 0.00203f
C5224 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_47816_6284# 0.0202f
C5225 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 a_47858_n2243# 0.0101f
C5226 RST a_50316_10154# 9.41e-19
C5227 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_39684_n10028# 0.00695f
C5228 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 0.205f
C5229 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_53309_n15631# 1.52e-20
C5230 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB a_23123_n7106# 1.35e-20
C5231 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT 0.345f
C5232 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB a_23184_n9840# 0.00964f
C5233 F0 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 4.45e-19
C5234 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_47994_n18696# 0.0697f
C5235 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 0.209f
C5236 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.749f
C5237 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 a_27324_5062# 0.0157f
C5238 RST a_25650_n1899# 7.66e-19
C5239 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.00586f
C5240 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 a_28663_n17626# 1.09e-20
C5241 Vdiv105 a_43671_7266# 0.2f
C5242 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.103f
C5243 RST a_23589_6159# 0.00105f
C5244 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 2.29e-19
C5245 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K a_53129_n19793# 0.0027f
C5246 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN 0.519f
C5247 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 6.24e-20
C5248 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 0.399f
C5249 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_47430_n18696# 2.79e-20
C5250 a_47332_n5176# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0203f
C5251 VDD105 a_45927_6284# 3.56e-19
C5252 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_23025_6159# 0.0697f
C5253 RST a_48712_n17599# 0.00119f
C5254 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_35454_n16636# 0.0203f
C5255 VDD105 a_47970_5143# 0.00101f
C5256 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_47338_n6273# 1.75e-19
C5257 CLK CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 0.00527f
C5258 CLK_div_96_mag_0.JK_FF_mag_0.Q a_23142_n2930# 0.0101f
C5259 RST CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 0.0768f
C5260 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.00112f
C5261 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 0.408f
C5262 VDD99 a_26046_n16632# 2.21e-19
C5263 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 a_36103_n10028# 0.00789f
C5264 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_45564_9057# 0.0732f
C5265 CLK_div_108_new_mag_0.JK_FF_mag_1.Q a_51803_n5724# 0.069f
C5266 a_53785_2768# a_53945_2768# 0.0504f
C5267 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 2.57e-20
C5268 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C5269 F0 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 0.197f
C5270 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00425f
C5271 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN a_43993_n13477# 2.4e-20
C5272 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 a_48324_n15585# 0.069f
C5273 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.109f
C5274 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_50675_n5724# 1.43e-19
C5275 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 1.34e-19
C5276 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 a_53126_6240# 0.0101f
C5277 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 0.00113f
C5278 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT a_54664_n10161# 1.17e-20
C5279 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_36673_n8887# 0.00378f
C5280 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 0.104f
C5281 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 8.64e-20
C5282 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_44170_2768# 0.00964f
C5283 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 2.98e-19
C5284 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 2.81e-20
C5285 VDD mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.OUT 0.634f
C5286 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 2.89e-20
C5287 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_46974_n2243# 2.81e-19
C5288 RST a_44971_n17599# 0.00283f
C5289 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_23129_n6009# 8.66e-20
C5290 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 1.22f
C5291 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_26368_n2996# 2.88e-20
C5292 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 2.59e-21
C5293 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.011f
C5294 RST a_44235_6240# 9.5e-19
C5295 VDD108 a_52652_n10117# 0.00149f
C5296 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 2.19f
C5297 RST a_47086_5143# 0.00186f
C5298 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.209f
C5299 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.121f
C5300 a_54027_n16728# a_54187_n16728# 0.0504f
C5301 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.977f
C5302 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT a_51652_2768# 1.17e-20
C5303 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK a_50310_n15627# 1.87e-19
C5304 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 5.32e-19
C5305 RST a_25292_10099# 0.00151f
C5306 a_51598_9057# a_51758_9057# 0.0504f
C5307 Vdiv93 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 4.46e-19
C5308 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0698f
C5309 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_29341_n16634# 0.0733f
C5310 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT 3.11e-19
C5311 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 a_32865_n15491# 0.0059f
C5312 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 a_42083_n15712# 0.0177f
C5313 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT m3_20882_n11188# 0.00256f
C5314 CLK_div_96_mag_0.JK_FF_mag_2.QB a_28743_n1899# 1.26e-20
C5315 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 0.0905f
C5316 RST a_51487_n10161# 0.00218f
C5317 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 9.06e-20
C5318 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 a_32175_n17626# 0.00335f
C5319 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 a_44841_n2243# 0.0101f
C5320 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 3.77e-20
C5321 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_30760_n20290# 0.00168f
C5322 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_53303_n16728# 1.17e-20
C5323 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_27170_6159# 0.0114f
C5324 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_37391_n9984# 0.069f
C5325 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K a_50874_n15583# 1.39e-19
C5326 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 a_24307_5062# 0.0157f
C5327 CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 a_40972_n9984# 0.0157f
C5328 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_25465_n6010# 8.64e-19
C5329 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00152f
C5330 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 0.026f
C5331 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 0.0365f
C5332 VDD90 a_26266_11196# 9.82e-19
C5333 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.00656f
C5334 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT 0.00169f
C5335 CLK a_26189_n6010# 0.00539f
C5336 VDD110 a_45695_n17599# 0.00152f
C5337 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_25484_n2996# 1.17e-20
C5338 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_25529_n743# 1.46e-19
C5339 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_53819_n5721# 0.0202f
C5340 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 0.00975f
C5341 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.108f
C5342 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 5.53e-20
C5343 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 7.24e-19
C5344 CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00393f
C5345 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_47994_n18696# 6.43e-21
C5346 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.121f
C5347 Vdiv110 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 5.47e-19
C5348 dec3x8_ibr_mag_0.and_3_ibr_5.IN3 dec3x8_ibr_mag_0.and_3_ibr_5.nand3_mag_ibr_0.OUT 0.117f
C5349 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.0591f
C5350 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB 2e-21
C5351 Vdiv105 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 4.78e-19
C5352 Vdiv108 a_51439_n2199# 7.3e-19
C5353 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_23552_n1789# 0.011f
C5354 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0894f
C5355 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_23948_n18723# 4.52e-20
C5356 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_45039_n5176# 0.069f
C5357 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 1.58e-20
C5358 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_44619_n16724# 0.0102f
C5359 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 0.12f
C5360 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.124f
C5361 RST a_43895_n16724# 8.14e-19
C5362 a_35032_n17626# a_35192_n17626# 0.0504f
C5363 Vdiv110 a_54663_1671# 2.22e-19
C5364 VDD96 Vdiv90 2.48f
C5365 RST a_44841_n2243# 0.00186f
C5366 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 4.52e-20
C5367 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_21995_n7106# 0.0059f
C5368 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00301f
C5369 CLK_div_96_mag_0.JK_FF_mag_3.QB CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.25f
C5370 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0343f
C5371 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.803f
C5372 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 1.35e-20
C5373 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_30342_11196# 0.0731f
C5374 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_29618_11196# 0.00696f
C5375 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 0.273f
C5376 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.257f
C5377 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT a_46867_7960# 0.00138f
C5378 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 8.16e-20
C5379 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0905f
C5380 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 3.61e-21
C5381 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00718f
C5382 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 a_29208_10099# 0.069f
C5383 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 0.00183f
C5384 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 0.00154f
C5385 a_44793_5143# a_44953_5143# 0.0504f
C5386 RST CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 0.105f
C5387 CLK a_29777_5062# 6.02e-19
C5388 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 0.163f
C5389 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0115f
C5390 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN 0.118f
C5391 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_44619_n16724# 0.0203f
C5392 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB a_25502_n9875# 0.00695f
C5393 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_51551_5187# 0.00378f
C5394 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 0.273f
C5395 CLK_div_96_mag_0.JK_FF_mag_0.Q CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 1.48e-20
C5396 VDD90 a_29778_11196# 2.21e-19
C5397 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 a_54033_n15587# 0.0697f
C5398 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_54456_n2199# 0.0036f
C5399 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 0.00183f
C5400 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.00656f
C5401 CLK_div_100_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT 0.11f
C5402 VDD100 a_45405_n2199# 0.00152f
C5403 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 a_54187_n16728# 8.64e-19
C5404 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00118f
C5405 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 0.0432f
C5406 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 a_23709_810# 1.46e-19
C5407 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.00384f
C5408 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN a_23948_n13382# 2.7e-20
C5409 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 3.08e-21
C5410 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_26349_n6010# 0.0202f
C5411 a_39844_n10028# m3_20882_n11188# 3.55e-19
C5412 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 a_25420_n13385# 0.0115f
C5413 CLK_div_105_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 5.13e-19
C5414 VDD96 a_27342_n1855# 6.86e-19
C5415 a_31352_6115# a_31512_6115# 0.0504f
C5416 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0592f
C5417 CLK CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 6.28e-21
C5418 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 4.52e-20
C5419 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.306f
C5420 VDD110 a_44253_n18696# 0.00752f
C5421 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_52161_n19793# 1.45e-20
C5422 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT 0.122f
C5423 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT m3_20882_n11188# 0.00187f
C5424 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K 5.7e-19
C5425 VDD90 a_26196_5018# 0.00101f
C5426 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.43f
C5427 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_44977_n18696# 0.0697f
C5428 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 2.81e-20
C5429 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 a_24391_n20290# 0.0134f
C5430 a_31577_n15535# a_31737_n15535# 0.0504f
C5431 a_29241_7256# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 2.36e-22
C5432 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_44235_6240# 0.0732f
C5433 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.122f
C5434 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 8.58e-20
C5435 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT Vdiv108 0.265f
C5436 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT 0.342f
C5437 RST a_43719_n120# 0.00198f
C5438 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C5439 CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 2.51e-20
C5440 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.231f
C5441 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 2.81e-20
C5442 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.00975f
C5443 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.391f
C5444 CLK CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 0.00547f
C5445 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 a_53216_n10117# 0.069f
C5446 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 0.0435f
C5447 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 0.231f
C5448 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_24391_n20290# 1.4e-19
C5449 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_43760_1671# 0.00118f
C5450 RST CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.00239f
C5451 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.209f
C5452 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_51729_n17599# 0.0036f
C5453 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0501f
C5454 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.994f
C5455 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_44321_n6273# 3.33e-19
C5456 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_1.IN2 0.109f
C5457 CLK CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 7.03e-21
C5458 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 Vdiv105 0.269f
C5459 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 1.03e-19
C5460 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_47338_n6273# 0.0697f
C5461 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 9.73e-19
C5462 VDD105 a_51040_10154# 0.00123f
C5463 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 8.94e-19
C5464 a_35747_n1222# Vdiv99 1.87e-19
C5465 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_43963_n1146# 0.0203f
C5466 RST CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 1.55e-19
C5467 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 0.108f
C5468 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_2.OUT CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_0.OUT 0.00183f
C5469 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 8.2e-19
C5470 RST a_33583_n16588# 0.00106f
C5471 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 3.42e-19
C5472 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 0.0327f
C5473 VDD99 CLK_div_96_mag_0.JK_FF_mag_5.QB 7.46e-19
C5474 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00544f
C5475 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.16f
C5476 VDD108 a_53089_n6862# 0.00108f
C5477 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00335f
C5478 VDD100 a_46755_574# 3.14e-19
C5479 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_29623_6159# 2.96e-19
C5480 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 a_50204_2768# 0.0036f
C5481 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_0.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.49e-19
C5482 dec3x8_ibr_mag_0.and_3_ibr_4.nand3_mag_ibr_0.OUT a_37328_6265# 3.58e-20
C5483 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_24901_n6010# 0.00378f
C5484 RST a_26974_1919# 0.00173f
C5485 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.00145f
C5486 CLK CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.29e-19
C5487 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT 0.998f
C5488 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 7.08e-20
C5489 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.0718f
C5490 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN a_32750_n7675# 4.15e-20
C5491 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT 1.69e-19
C5492 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_21902_n8787# 0.00119f
C5493 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 0.0655f
C5494 VDD108 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.657f
C5495 RST a_25322_n16632# 0.00125f
C5496 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT 0.649f
C5497 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 1.65f
C5498 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB 9.12e-20
C5499 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.00975f
C5500 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 5.98e-20
C5501 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.051f
C5502 RST CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.205f
C5503 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_39126_n8931# 0.0732f
C5504 RST a_51393_n6821# 0.00137f
C5505 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 a_46889_9057# 9.45e-19
C5506 RST a_49752_10154# 9.66e-19
C5507 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 a_47698_n2243# 0.0102f
C5508 CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 1.53e-19
C5509 F0 Vdiv108 3.98e-19
C5510 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 a_23948_n13382# 0.0202f
C5511 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 mux_8x1_ibr_0.mux_2x1_ibr_0.I0 0.0073f
C5512 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_52002_n15583# 0.0114f
C5513 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN 0.0181f
C5514 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB a_22620_n9884# 0.00696f
C5515 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_51285_n1102# 0.0059f
C5516 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 1.89e-19
C5517 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.00447f
C5518 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 a_26760_5062# 0.00859f
C5519 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 0.249f
C5520 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 2.56e-19
C5521 RST a_25490_n1899# 9.2e-19
C5522 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.653f
C5523 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB 7.08e-20
C5524 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.348f
C5525 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN a_40818_n8887# 4.94e-20
C5526 RST a_23025_6159# 7.59e-20
C5527 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 0.12f
C5528 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT 0.0951f
C5529 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 2.86f
C5530 a_47332_n5176# a_47492_n5176# 0.0504f
C5531 a_46768_n5176# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 1.5e-20
C5532 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 0.0014f
C5533 VDD105 a_45363_6284# 3.14e-19
C5534 VDD99 CLK_div_96_mag_0.JK_FF_mag_3.Q 0.00133f
C5535 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_34890_n16636# 1.5e-20
C5536 CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 1.52e-20
C5537 VDD105 a_47810_5143# 0.00123f
C5538 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.0063f
C5539 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 6.96e-19
C5540 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB 3.21e-19
C5541 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN 1e-19
C5542 CLK_div_96_mag_0.JK_FF_mag_0.Q a_22982_n2930# 0.0102f
C5543 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.0485f
C5544 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 a_55357_n20487# 0.019f
C5545 VDD110 a_42521_n13474# 0.165f
C5546 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 a_35943_n10028# 0.00335f
C5547 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_45000_9057# 0.00378f
C5548 CLK_div_108_new_mag_0.JK_FF_mag_1.Q a_51239_n5724# 3.74e-21
C5549 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 1.47e-20
C5550 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.338f
C5551 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 3e-20
C5552 CLK a_21995_n7106# 3.7e-19
C5553 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 0.977f
C5554 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_50111_n5768# 0.00119f
C5555 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 a_51961_6284# 9.45e-19
C5556 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT a_54504_n10161# 1.5e-20
C5557 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 a_53280_5143# 0.00164f
C5558 a_50675_n5724# CLK_div_108_new_mag_0.CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 1.46e-22
C5559 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_36109_n8931# 0.0732f
C5560 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB 0.25f
C5561 RST CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 6.71e-19
C5562 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_43606_2768# 0.0811f
C5563 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN 2.86e-19
C5564 CLK_div_105_mag_0.CLK_div_10_mag_1.CLK CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 4.19e-19
C5565 RST a_44407_n17599# 0.0037f
C5566 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_26208_n2996# 9.1e-19
C5567 a_23703_n287# CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 3.23e-20
C5568 VDD108 a_51647_n10161# 0.00743f
C5569 RST a_44075_6240# 8.88e-19
C5570 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.195f
C5571 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT m3_20882_n11188# 0.00379f
C5572 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 a_29801_1733# 0.0134f
C5573 a_52156_n16680# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 4.81e-20
C5574 RST a_46081_5187# 9.66e-19
C5575 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_45753_n15583# 0.00118f
C5576 RST CLK_div_96_mag_0.JK_FF_mag_2.Q 0.324f
C5577 VDD99 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 0.00101f
C5578 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT 0.664f
C5579 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 2.11e-19
C5580 CLK CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 0.00862f
C5581 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.179f
C5582 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 a_50763_n10161# 8.64e-19
C5583 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.00441f
C5584 CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 3.64e-20
C5585 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT a_51492_2768# 1.5e-20
C5586 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 0.00213f
C5587 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 5.13e-19
C5588 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 8.94e-19
C5589 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 0.0138f
C5590 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK a_50150_n15627# 2.69e-19
C5591 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN 0.112f
C5592 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_55357_n20487# 3.02e-19
C5593 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 7.97e-19
C5594 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_29181_n16634# 0.0203f
C5595 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 a_32301_n15491# 0.0697f
C5596 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_23594_n8743# 0.00372f
C5597 CLK_div_96_mag_0.JK_FF_mag_2.QB a_28583_n1899# 1.62e-20
C5598 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.192f
C5599 RST a_50923_n10161# 0.00212f
C5600 Vdiv99 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN 0.0109f
C5601 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.0215f
C5602 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 a_32015_n17626# 0.00789f
C5603 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 a_44681_n2243# 0.0102f
C5604 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.IN2 a_35747_n1222# 0.00372f
C5605 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.467f
C5606 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C5607 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 CLK_div_99_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 8.04e-19
C5608 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_26606_6159# 2.96e-19
C5609 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 0.321f
C5610 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.792f
C5611 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 a_23743_5062# 0.00859f
C5612 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K a_50310_n15627# 8.21e-19
C5613 CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 a_40408_n9984# 0.00859f
C5614 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 0.0435f
C5615 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.121f
C5616 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0622f
C5617 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 a_23948_n13382# 0.0186f
C5618 VDD90 a_25702_11196# 0.00149f
C5619 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_50987_5143# 2.88e-20
C5620 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.109f
C5621 CLK a_25625_n6010# 0.00148f
C5622 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C5623 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_24153_6159# 0.00118f
C5624 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 1.15f
C5625 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.109f
C5626 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 0.0129f
C5627 VDD96 dec3x8_ibr_mag_0.and_3_ibr_5.IN3 0.00104f
C5628 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 2.36e-20
C5629 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT a_52839_n5# 3.92e-20
C5630 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 2.81e-20
C5631 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.121f
C5632 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 dec3x8_ibr_mag_0.and_3_ibr_4.nand3_mag_ibr_0.OUT 5.81e-20
C5633 VDD93 a_39684_n10028# 2.21e-19
C5634 RST CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT 0.107f
C5635 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00183f
C5636 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_48268_n1102# 0.0059f
C5637 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.0592f
C5638 Vdiv110 a_36873_280# 2.66e-19
C5639 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 6.02e-20
C5640 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.28f
C5641 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 3.6e-19
C5642 a_23019_5018# a_23179_5018# 0.0504f
C5643 CLK a_35186_n18723# 0.0101f
C5644 a_27381_n699# CLK_div_96_mag_0.JK_FF_mag_2.QB 5.3e-20
C5645 Vdiv108 a_50875_n2243# 6.67e-19
C5646 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.175f
C5647 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 0.233f
C5648 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_48888_n15585# 0.069f
C5649 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_22988_n1789# 1.43e-19
C5650 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.08f
C5651 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 9.24e-20
C5652 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_50304_n16724# 4.66e-19
C5653 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_44055_n16724# 0.0152f
C5654 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 4.28e-19
C5655 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.768f
C5656 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_50310_n15627# 1.16e-20
C5657 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0717f
C5658 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00119f
C5659 Vdiv110 a_54503_1671# 1.8e-19
C5660 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 0.517f
C5661 VDD96 a_33405_7558# 0.00829f
C5662 RST a_44681_n2243# 8.64e-19
C5663 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.00118f
C5664 a_22711_n14504# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT 0.0732f
C5665 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_29778_11196# 9.1e-19
C5666 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.36f
C5667 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.00157f
C5668 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_29054_11196# 0.00964f
C5669 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT a_51647_n10161# 1.17e-20
C5670 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB 3.49e-19
C5671 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT a_43831_7266# 0.0294f
C5672 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT 0.748f
C5673 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.187f
C5674 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 a_28644_10099# 0.00372f
C5675 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.00584f
C5676 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0622f
C5677 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.519f
C5678 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_47858_n2243# 2.88e-20
C5679 a_35943_n10028# a_36103_n10028# 0.0504f
C5680 CLK a_29213_5018# 5.65e-19
C5681 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.768f
C5682 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB 0.911f
C5683 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 1.36e-20
C5684 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.IN2 0.0655f
C5685 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.121f
C5686 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_44055_n16724# 1.5e-20
C5687 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_50987_5143# 0.0733f
C5688 CLK CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 0.00347f
C5689 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.121f
C5690 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 a_29680_398# 4.9e-20
C5691 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 3.4e-19
C5692 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 CLK_div_96_mag_0.JK_FF_mag_4.QB 0.199f
C5693 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT 0.053f
C5694 VDD100 a_44841_n2243# 0.00101f
C5695 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_23142_n2930# 2.88e-20
C5696 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 8.59e-20
C5697 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_26189_n6010# 0.0731f
C5698 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN 0.0549f
C5699 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_26778_n1855# 1.71e-20
C5700 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 7.08e-20
C5701 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN 7e-19
C5702 a_39684_n10028# m3_20882_n11188# 3.55e-19
C5703 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 0.359f
C5704 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0118f
C5705 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 4.52e-20
C5706 VDD96 a_26778_n1855# 3.14e-19
C5707 VDD93 Vdiv93 2.97f
C5708 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 0.413f
C5709 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 0.327f
C5710 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 0.109f
C5711 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.401f
C5712 Vdiv108 CLK_div_108_new_mag_0.JK_FF_mag_1.Q 0.158f
C5713 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_40818_n8887# 0.012f
C5714 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 0.144f
C5715 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_47528_n9019# 0.0202f
C5716 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C5717 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_0.OUT a_26214_n1855# 0.00378f
C5718 F0 Vdiv93 0.111f
C5719 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.399f
C5720 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.235f
C5721 VDD90 a_26036_5018# 0.00123f
C5722 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 2e-19
C5723 CLK_div_96_mag_0.JK_FF_mag_4.QB CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.0113f
C5724 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K Vdiv110 0.0121f
C5725 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 1.98e-19
C5726 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_44075_6240# 0.0203f
C5727 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 6.33e-20
C5728 RST a_43559_n120# 0.00189f
C5729 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.00602f
C5730 Vdiv Vdiv100 2.62e-19
C5731 Vdiv110 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 0.0013f
C5732 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.0496f
C5733 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 a_52652_n10117# 0.00372f
C5734 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 7.49e-20
C5735 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 a_50316_10154# 0.069f
C5736 CLK_div_96_mag_0.JK_FF_mag_5.Q CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 0.0254f
C5737 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_96_mag_0.JK_FF_mag_2.Q 2.14e-19
C5738 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT 2.81e-20
C5739 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_47190_n16726# 1.46e-19
C5740 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.0432f
C5741 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 1.18f
C5742 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.0635f
C5743 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 1.05e-20
C5744 RST CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K 0.447f
C5745 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN 0.299f
C5746 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.648f
C5747 F0 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 0.378f
C5748 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_24922_n17626# 8.64e-19
C5749 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.0622f
C5750 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.318f
C5751 VDD105 a_50880_10154# 0.00101f
C5752 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 3.26e-20
C5753 dec3x8_ibr_mag_0.and_3_ibr_6.nand3_mag_ibr_0.OUT dec3x8_ibr_mag_0.and_3_ibr_7.nand3_mag_ibr_0.OUT 6.66e-19
C5754 RST a_33019_n16588# 0.00129f
C5755 CLK_div_105_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00943f
C5756 VDD VDD99 0.331f
C5757 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT 0.00335f
C5758 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 a_30209_7256# 0.0112f
C5759 CLK_div_96_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 8.04e-19
C5760 CLK_div_108_new_mag_0.JK_FF_mag_1.QB CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0383f
C5761 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.0979f
C5762 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 2.29e-20
C5763 dec3x8_ibr_mag_0.and_3_ibr_5.IN3 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 0.0986f
C5764 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_51397_6284# 0.0059f
C5765 VDD108 a_51957_n6821# 3.14e-19
C5766 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB 0.0378f
C5767 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT 0.121f
C5768 F1 Vdiv110 0.117f
C5769 VDD VDD100 0.401f
C5770 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 a_23289_n6009# 0.00144f
C5771 VDD100 a_43719_n120# 0.234f
C5772 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_29059_6159# 3.25e-19
C5773 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0889f
C5774 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 a_46614_n6273# 0.00149f
C5775 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 1.08e-20
C5776 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_55161_n15587# 0.00118f
C5777 dec3x8_ibr_mag_0.and_3_ibr_4.nand3_mag_ibr_0.OUT a_37168_6265# 6.08e-20
C5778 RST a_26814_1919# 0.0013f
C5779 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.322f
C5780 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 6.23e-20
C5781 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.519f
C5782 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.748f
C5783 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN 0.0116f
C5784 RST a_54658_n9064# 7.78e-19
C5785 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 3.87f
C5786 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_38966_n8931# 0.0203f
C5787 RST a_50829_n6865# 0.00206f
C5788 F1 a_37436_n1822# 0.0144f
C5789 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_54663_1671# 0.0203f
C5790 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 5.7e-20
C5791 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 a_47134_n2243# 0.00789f
C5792 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_24127_10099# 0.0203f
C5793 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_48534_5187# 0.00378f
C5794 VDD99 a_33583_n16588# 3.14e-19
C5795 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_51438_n15583# 2.96e-19
C5796 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB a_22460_n9884# 0.00695f
C5797 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 8.58e-20
C5798 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00107f
C5799 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.00125f
C5800 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 3.38e-19
C5801 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_52156_n16680# 0.0811f
C5802 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_50721_n1102# 0.0697f
C5803 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 a_26196_5018# 0.0101f
C5804 RST a_24116_n1789# 9.81e-19
C5805 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.16f
C5806 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.00434f
C5807 a_46608_n5176# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 1.17e-20
C5808 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.783f
C5809 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.038f
C5810 VDD105 a_44799_6284# 3.14e-19
C5811 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT 0.159f
C5812 CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.338f
C5813 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_34730_n16636# 1.17e-20
C5814 VDD105 a_47246_5143# 0.00863f
C5815 CLK_div_96_mag_0.JK_FF_mag_0.QB CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.25f
C5816 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 0.0718f
C5817 CLK_div_96_mag_0.JK_FF_mag_0.Q a_22418_n2930# 0.00789f
C5818 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_28823_n17626# 1.17e-20
C5819 VDD99 a_25322_n16632# 2.21e-19
C5820 dec3x8_ibr_mag_0.and_3_ibr_3.nand3_mag_ibr_0.OUT Vdiv 5.94e-20
C5821 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 2.73e-21
C5822 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.652f
C5823 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.124f
C5824 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_44511_n9019# 0.0202f
C5825 CLK a_21431_n7106# 3.7e-19
C5826 a_26208_n2996# a_26368_n2996# 0.0504f
C5827 F1 dec3x8_ibr_mag_0.and_3_ibr_1.nand3_mag_ibr_0.OUT 0.217f
C5828 a_49945_n6865# a_50105_n6865# 0.0504f
C5829 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT 0.267f
C5830 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_44888_1671# 0.0202f
C5831 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.122f
C5832 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 a_51397_6284# 6.06e-21
C5833 RST CLK_div_105_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 0.00649f
C5834 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.00586f
C5835 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT a_53940_n10161# 0.0203f
C5836 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.198f
C5837 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.397f
C5838 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 a_36202_6821# 0.00418f
C5839 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 0.11f
C5840 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 a_53120_5143# 0.00117f
C5841 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_35949_n8931# 0.0203f
C5842 RST CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0042f
C5843 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.0792f
C5844 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0622f
C5845 RST a_32169_n18723# 7.78e-19
C5846 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 8.58e-20
C5847 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_30435_n1855# 0.00118f
C5848 RST CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.178f
C5849 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB a_23030_n8743# 5e-20
C5850 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 1.35e-19
C5851 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN a_46867_7960# 0.069f
C5852 RST a_44247_n17599# 0.00334f
C5853 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_25806_n17626# 0.0202f
C5854 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.403f
C5855 RST CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0235f
C5856 CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 8.16e-19
C5857 CLK_div_96_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 2.34e-19
C5858 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 0.00574f
C5859 F1 a_37436_880# 0.0145f
C5860 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_25644_n2996# 0.0731f
C5861 VDD108 a_51487_n10161# 0.00305f
C5862 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 0.36f
C5863 a_53309_n15631# a_53469_n15631# 0.0504f
C5864 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 0.0129f
C5865 CLK CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 5.57e-19
C5866 RST a_45517_5187# 9.41e-19
C5867 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 0.0145f
C5868 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_0.OUT CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00137f
C5869 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_45189_n15583# 0.011f
C5870 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 a_50232_n7685# 0.0134f
C5871 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.802f
C5872 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 0.21f
C5873 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 0.124f
C5874 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.398f
C5875 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00233f
C5876 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 1.15f
C5877 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 m3_20882_n11188# 0.00199f
C5878 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT a_50928_2768# 0.0203f
C5879 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 2.47e-19
C5880 CLK a_43671_7266# 4.82e-19
C5881 RST CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 0.696f
C5882 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB a_25625_n6010# 0.00695f
C5883 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT 0.00154f
C5884 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN 0.00525f
C5885 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_55197_n20487# 9.21e-20
C5886 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_28617_n16634# 1.5e-20
C5887 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK a_50304_n16724# 0.00192f
C5888 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 a_25532_3016# 0.0036f
C5889 CLK_div_96_mag_0.JK_FF_mag_2.QB CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.0592f
C5890 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.161f
C5891 RST a_32076_6159# 2.78e-19
C5892 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0871f
C5893 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_23030_n8743# 0.069f
C5894 Vdiv99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 3.98e-19
C5895 RST a_50763_n10161# 0.00203f
C5896 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.4f
C5897 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 9.82e-21
C5898 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.103f
C5899 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 a_31451_n17626# 0.0102f
C5900 RST CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00516f
C5901 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 1.36e-19
C5902 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_48380_6284# 0.0059f
C5903 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 a_44117_n2243# 0.00789f
C5904 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 9.71e-20
C5905 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C5906 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT a_54187_n16728# 2.88e-20
C5907 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_26042_6159# 3.25e-19
C5908 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.0378f
C5909 CLK CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.00131f
C5910 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K a_50150_n15627# 0.00598f
C5911 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 a_23179_5018# 0.0101f
C5912 CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 a_39844_n10028# 0.0101f
C5913 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.261f
C5914 a_52002_n15583# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 4.52e-20
C5915 VDD90 a_25138_11196# 0.00149f
C5916 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 2.48e-20
C5917 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT 0.572f
C5918 CLK a_25465_n6010# 0.00145f
C5919 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_50827_5143# 9.1e-19
C5920 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.913f
C5921 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 a_30398_n699# 0.0157f
C5922 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_23589_6159# 0.011f
C5923 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.108f
C5924 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 2.27e-20
C5925 CLK_div_96_mag_0.JK_FF_mag_2.Q CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.235f
C5926 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT 0.647f
C5927 CLK CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 1.29e-19
C5928 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 a_35614_n16636# 8.64e-19
C5929 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 1.98e-19
C5930 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 6.88e-21
C5931 VDD93 a_39120_n10028# 0.00305f
C5932 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_47704_n1102# 0.0697f
C5933 dec3x8_ibr_mag_0.and_3_ibr_5.IN3 a_37168_6265# 0.00657f
C5934 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 1.89e-20
C5935 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.769f
C5936 CLK a_35026_n18723# 0.00939f
C5937 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 0.00488f
C5938 Vdiv108 a_50715_n2243# 6.67e-19
C5939 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.235f
C5940 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 1.9e-20
C5941 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 4.1e-21
C5942 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_22424_n1833# 0.00119f
C5943 RST CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.285f
C5944 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C5945 CLK_div_90_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN Vdiv90 0.00226f
C5946 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 a_52951_7381# 0.01f
C5947 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_50144_n16724# 6.02e-19
C5948 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 3.78e-20
C5949 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_43895_n16724# 0.0124f
C5950 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT m3_20882_n11188# 0.00155f
C5951 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 8.64e-20
C5952 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 3.09e-19
C5953 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 0.342f
C5954 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_50150_n15627# 1.49e-20
C5955 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_23289_n6009# 1.17e-20
C5956 Vdiv110 a_53939_1671# 4.73e-20
C5957 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_47264_n17599# 1.04e-19
C5958 VDD96 a_33245_7558# 0.00428f
C5959 RST CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 0.0547f
C5960 CLK_div_100_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 a_43719_n120# 9.02e-19
C5961 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 a_52139_n18696# 0.00372f
C5962 F1 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT 1.54e-19
C5963 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 6.7e-19
C5964 a_22551_n14504# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT 0.0202f
C5965 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_29618_11196# 2.88e-20
C5966 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 0.0638f
C5967 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 8.16e-20
C5968 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 3.94e-19
C5969 CLK CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 1.29e-19
C5970 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_28490_11196# 0.0811f
C5971 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 a_28644_10099# 0.069f
C5972 F1 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT 0.00305f
C5973 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT a_51487_n10161# 1.5e-20
C5974 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 4.2e-20
C5975 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT a_43671_7266# 0.00894f
C5976 CLK_div_100_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 4.25e-20
C5977 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0636f
C5978 RST CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.264f
C5979 CLK_div_105_mag_0.CLK_div_10_mag_1.CLK a_55179_7683# 0.198f
C5980 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 0.0154f
C5981 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 1.83f
C5982 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_47698_n2243# 9.1e-19
C5983 CLK a_29053_5018# 5.65e-19
C5984 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_33429_n15491# 0.00118f
C5985 VDD93 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 3.57e-19
C5986 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.338f
C5987 a_51871_n5# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 1.45e-20
C5988 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 2.57e-19
C5989 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_50827_5143# 0.0203f
C5990 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 2.37f
C5991 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_43895_n16724# 1.17e-20
C5992 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 0.205f
C5993 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.397f
C5994 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 a_36873_n1222# 0.00372f
C5995 VDD90 a_29054_11196# 3.14e-19
C5996 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT 3.09e-19
C5997 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.0622f
C5998 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0759f
C5999 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT 0.121f
C6000 VDD F2 4.51f
C6001 VDD100 a_44681_n2243# 0.00123f
C6002 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 2.57e-19
C6003 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.00627f
C6004 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_43826_n7684# 0.00263f
C6005 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 5.05e-20
C6006 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_22982_n2930# 9.1e-19
C6007 CLK_div_100_mag_0.CLK_div_10_mag_1.CLK CLK_div_100_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 2.16e-19
C6008 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_25625_n6010# 9.1e-19
C6009 CLK CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 0.126f
C6010 a_39120_n10028# m3_20882_n11188# 8.45e-19
C6011 VDD96 a_26214_n1855# 3.14e-19
C6012 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.651f
C6013 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB a_47534_n10160# 0.00695f
C6014 VDD VDD108 0.62f
C6015 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_1.IN2 1.48e-20
C6016 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_0.QB 1.4e-19
C6017 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_26778_n1855# 0.0059f
C6018 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_40254_n8887# 2.96e-19
C6019 a_54907_297# a_55067_297# 0.186f
C6020 Vdiv100 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.OUT 0.00282f
C6021 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_46964_n9019# 4.52e-20
C6022 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.768f
C6023 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.00118f
C6024 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_54537_n6818# 0.0036f
C6025 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 4.75e-20
C6026 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 7.16e-20
C6027 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00118f
C6028 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_0.OUT a_25650_n1899# 0.0732f
C6029 VDD90 a_25472_5018# 0.00863f
C6030 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.348f
C6031 CLK CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.00668f
C6032 a_54182_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0733f
C6033 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN 0.128f
C6034 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 1.1e-19
C6035 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_29213_5018# 2.88e-20
C6036 RST a_23863_n287# 9.45e-19
C6037 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB m3_20882_n11188# 0.00467f
C6038 CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN a_29087_8532# 0.132f
C6039 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_50447_n18696# 9.32e-19
C6040 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 0.00477f
C6041 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_27375_n17626# 0.0036f
C6042 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.313f
C6043 CLK CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 1.17e-20
C6044 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 a_49752_10154# 0.00372f
C6045 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.101f
C6046 CLK_div_96_mag_0.JK_FF_mag_5.Q CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_1.IN2 0.109f
C6047 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_2.OUT CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_0.OUT 0.00183f
C6048 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0343f
C6049 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C6050 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 6.01e-19
C6051 CLK_div_108_new_mag_0.JK_FF_mag_1.QB a_51957_n6821# 0.0811f
C6052 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 a_51764_10154# 0.001f
C6053 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 0.283f
C6054 RST a_37801_n8887# 7.24e-19
C6055 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C6056 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0636f
C6057 RST CLK_div_96_mag_0.JK_FF_mag_3.QB 0.119f
C6058 VDD105 a_50316_10154# 0.00152f
C6059 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 2.89e-20
C6060 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 a_29213_n7028# 0.00952f
C6061 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 0.00205f
C6062 dec3x8_ibr_mag_0.and_3_ibr_6.nand3_mag_ibr_0.OUT a_39580_6265# 3.58e-20
C6063 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 1.53e-19
C6064 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 0.412f
C6065 VDD96 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 1.37f
C6066 RST a_32455_n16632# 0.00222f
C6067 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.768f
C6068 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.00118f
C6069 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 a_29241_7256# 0.00929f
C6070 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C6071 CLK_div_96_mag_0.JK_FF_mag_0.Q CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C6072 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_53129_n19793# 0.01f
C6073 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_50833_6284# 0.0697f
C6074 VDD108 a_51393_n6821# 3.14e-19
C6075 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.289f
C6076 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 a_23129_n6009# 0.00169f
C6077 VDD100 a_43559_n120# 0.0407f
C6078 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 a_44779_n16724# 8.64e-19
C6079 CLK CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 0.00325f
C6080 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 9.96e-20
C6081 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 0.0659f
C6082 a_51015_7381# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 3.38e-20
C6083 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_28495_6115# 0.00392f
C6084 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0316f
C6085 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 0.636f
C6086 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 a_45449_n6273# 0.069f
C6087 Vdiv105 Vdiv96 0.00192f
C6088 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_54597_n15587# 0.011f
C6089 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT 0.122f
C6090 RST a_26250_1919# 3.52e-19
C6091 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT a_26343_n7107# 0.0203f
C6092 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.27f
C6093 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_54751_n16684# 0.0036f
C6094 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.122f
C6095 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 2.59e-21
C6096 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 3.23f
C6097 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0592f
C6098 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.122f
C6099 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K a_51481_n9064# 0.00392f
C6100 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 8.46e-19
C6101 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.24f
C6102 RST a_54498_n9064# 6.43e-19
C6103 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 a_45899_7960# 0.01f
C6104 F0 dec3x8_ibr_mag_0.and_3_ibr_6.nand3_mag_ibr_0.OUT 0.332f
C6105 RST a_50669_n6865# 0.00103f
C6106 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_54503_1671# 0.0732f
C6107 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00103f
C6108 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 a_46974_n2243# 0.00335f
C6109 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_23967_10099# 0.0732f
C6110 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 0.23f
C6111 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_4.IN2 CLK_div_96_mag_0.JK_FF_mag_5.QB 0.199f
C6112 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_50874_n15583# 3.08e-19
C6113 VDD99 a_33019_n16588# 3.14e-19
C6114 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_47970_5143# 0.0733f
C6115 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB Vdiv110 0.0101f
C6116 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_51592_n16680# 0.00964f
C6117 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK m3_20882_n11188# 4.97e-20
C6118 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_48252_n9063# 0.0203f
C6119 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 4.84e-19
C6120 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 a_26036_5018# 0.0102f
C6121 RST a_23552_n1789# 0.00163f
C6122 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.25f
C6123 VDD105 a_44235_6240# 2.66e-19
C6124 CLK CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 0.00791f
C6125 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.198f
C6126 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 m3_20882_n11188# 0.00141f
C6127 VDD105 a_47086_5143# 0.0123f
C6128 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 0.25f
C6129 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 6.63e-19
C6130 CLK_div_96_mag_0.JK_FF_mag_0.Q a_22258_n2930# 0.00335f
C6131 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_28663_n17626# 1.5e-20
C6132 CLK_div_108_new_mag_0.JK_FF_mag_1.Q a_50111_n5768# 2.79e-20
C6133 VDD93 a_40818_n8887# 3.56e-19
C6134 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_43947_n9019# 4.52e-20
C6135 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 4.31e-20
C6136 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 2.8e-19
C6137 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 5.52e-20
C6138 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 1.32e-21
C6139 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_44324_1671# 4.52e-20
C6140 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00137f
C6141 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.748f
C6142 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT a_53780_n10161# 0.0733f
C6143 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.00163f
C6144 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 a_49488_n13383# 0.00476f
C6145 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 a_52293_n17599# 0.00372f
C6146 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 a_36042_6821# 0.00284f
C6147 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 0.118f
C6148 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.471f
C6149 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_29871_n1855# 0.011f
C6150 RST a_32009_n18723# 6.43e-19
C6151 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 2.11e-21
C6152 RST a_35192_n17626# 5.2e-19
C6153 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_25646_n17626# 0.0731f
C6154 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_21841_n6009# 0.0036f
C6155 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_25484_n2996# 0.0202f
C6156 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 0.0529f
C6157 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00118f
C6158 VDD108 a_50923_n10161# 2.21e-19
C6159 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.00154f
C6160 CLK a_32175_n17626# 0.00117f
C6161 RST a_44953_5143# 0.00186f
C6162 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 0.198f
C6163 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_96_mag_0.JK_FF_mag_0.Q 3.42e-20
C6164 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_44625_n15583# 1.43e-19
C6165 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 a_54498_n9064# 0.00119f
C6166 VDD93 a_26790_n9831# 3.15e-19
C6167 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.0105f
C6168 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 0.00975f
C6169 a_53129_n19793# CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 2.94e-20
C6170 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.0654f
C6171 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 m3_20882_n11188# 7.32e-19
C6172 VDD110 a_41124_n14596# 2.21e-19
C6173 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_40408_n9984# 0.00378f
C6174 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT a_50768_2768# 0.0733f
C6175 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 0.0388f
C6176 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.0175f
C6177 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.397f
C6178 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 a_22711_n14504# 6.63e-20
C6179 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB a_25465_n6010# 0.00696f
C6180 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_28457_n16634# 1.17e-20
C6181 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 8.16e-20
C6182 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK a_50144_n16724# 0.00192f
C6183 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 a_48017_9057# 0.0697f
C6184 RST a_50199_n10117# 0.00121f
C6185 CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 CLK_div_105_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00357f
C6186 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 9.87e-20
C6187 VDD100 CLK_div_105_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 0.0024f
C6188 VDD99 a_32169_n18723# 2.21e-19
C6189 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN 0.519f
C6190 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 0.36f
C6191 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 a_31291_n17626# 0.0101f
C6192 RST Vdiv100 0.00629f
C6193 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 a_43957_n2243# 0.00335f
C6194 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_47816_6284# 0.0697f
C6195 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT a_54027_n16728# 9.1e-19
C6196 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 2.8e-19
C6197 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0301f
C6198 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_25478_6115# 0.00392f
C6199 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_51849_n1102# 0.00118f
C6200 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT 0.739f
C6201 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K a_48888_n15585# 8.11e-19
C6202 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 a_23019_5018# 0.0102f
C6203 CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 a_39684_n10028# 0.0102f
C6204 Vdiv108 CLK_div_108_new_mag_0.JK_FF_mag_0.QB 1.95f
C6205 RST CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.0172f
C6206 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.768f
C6207 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 a_30469_n16590# 0.00372f
C6208 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 0.124f
C6209 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_50263_5143# 0.0731f
C6210 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.199f
C6211 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 a_52156_n16680# 0.00372f
C6212 CLK a_24901_n6010# 0.00178f
C6213 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_23025_6159# 1.43e-19
C6214 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 a_29834_n699# 0.00859f
C6215 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0622f
C6216 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.012f
C6217 CLK CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00433f
C6218 a_36042_6821# a_36202_6821# 0.0504f
C6219 CLK CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT 0.3f
C6220 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 0.102f
C6221 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 3.92e-20
C6222 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN a_49488_n13383# 0.069f
C6223 VDD93 a_38960_n10028# 0.00743f
C6224 CLK CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_2.OUT 0.236f
C6225 VDD96 CLK_div_96_mag_0.JK_FF_mag_5.QB 0.914f
C6226 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.0576f
C6227 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_45235_n9063# 0.0203f
C6228 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0399f
C6229 VDD dec3x8_ibr_mag_0.and_3_ibr_5.nand3_mag_ibr_0.OUT 0.671f
C6230 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.159f
C6231 CLK a_34462_n18723# 6.43e-21
C6232 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.209f
C6233 a_48469_1671# a_48629_1671# 0.0504f
C6234 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_45612_1671# 0.00111f
C6235 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 2.86f
C6236 Vdiv108 a_50151_n2243# 0.00158f
C6237 RST CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.266f
C6238 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 0.0659f
C6239 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_96_mag_0.JK_FF_mag_3.QB 2.06e-19
C6240 RST a_47492_n5176# 0.00156f
C6241 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.121f
C6242 CLK_div_90_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_33405_7558# 5.39e-20
C6243 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT 0.00296f
C6244 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_49042_n16682# 0.0157f
C6245 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 3.07e-20
C6246 a_26790_n9831# m3_20882_n11188# 2.96e-19
C6247 RST CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 0.002f
C6248 CLK CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 5.96e-19
C6249 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_48888_n15585# 0.0114f
C6250 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 5.24e-20
C6251 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 0.191f
C6252 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_23129_n6009# 1.5e-20
C6253 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 1f
C6254 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 a_51575_n18696# 0.069f
C6255 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 1.99e-19
C6256 CLK_div_96_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_28828_1497# 0.069f
C6257 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_108_new_mag_0.JK_FF_mag_1.Q 0.107f
C6258 a_44321_n6273# CLK_div_108_new_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 5.01e-20
C6259 CLK_div_100_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 a_43559_n120# 2.44e-20
C6260 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 3.67e-20
C6261 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.019f
C6262 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 Vdiv 0.111f
C6263 a_22551_n14504# a_22711_n14504# 0.0504f
C6264 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 1.99e-19
C6265 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.00452f
C6266 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.198f
C6267 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 2.61e-19
C6268 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00158f
C6269 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN m3_20882_n11188# 0.00101f
C6270 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT a_50923_n10161# 0.0203f
C6271 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN 0.00253f
C6272 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.768f
C6273 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 RST 0.169f
C6274 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 1.82e-19
C6275 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 0.108f
C6276 CLK_div_105_mag_0.CLK_div_10_mag_1.CLK a_55019_7683# 0.0133f
C6277 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 1.36e-19
C6278 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 a_29341_n16634# 8.64e-19
C6279 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 a_22466_n8743# 6.43e-21
C6280 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_47134_n2243# 0.0731f
C6281 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 2.81e-20
C6282 CLK a_28489_5018# 0.00134f
C6283 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.00481f
C6284 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_32865_n15491# 0.011f
C6285 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 0.0334f
C6286 VDD96 CLK_div_96_mag_0.JK_FF_mag_3.Q 4f
C6287 CLK_div_90_mag_0.CLK_div_10_mag_0.CLK CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 0.149f
C6288 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_4.QB 0.25f
C6289 Vdiv93 CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 0.009f
C6290 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C6291 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.00871f
C6292 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_50263_5143# 1.5e-20
C6293 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 2.59e-21
C6294 CLK CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.00461f
C6295 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 a_51481_n9064# 0.00119f
C6296 VDD90 a_28490_11196# 3.14e-19
C6297 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_53168_n2243# 1.46e-19
C6298 VDD VDD105 0.475f
C6299 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_30187_6159# 7.4e-19
C6300 VDD100 a_44117_n2243# 0.00892f
C6301 VDD mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT 0.659f
C6302 a_48475_2768# a_48635_2768# 0.0504f
C6303 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 a_22421_810# 0.0036f
C6304 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 9.24e-20
C6305 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_22418_n2930# 0.0731f
C6306 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_25465_n6010# 2.88e-20
C6307 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.447f
C6308 a_38960_n10028# m3_20882_n11188# 8.45e-19
C6309 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT Vdiv110 2.57e-21
C6310 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT 0.121f
C6311 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB a_47374_n10160# 0.00696f
C6312 CLK_div_90_mag_0.CLK_div_10_mag_0.CLK a_22455_5018# 0.00164f
C6313 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 1.99e-19
C6314 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_26214_n1855# 0.0697f
C6315 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_39690_n8887# 1.75e-19
C6316 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 0.0591f
C6317 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN 0.517f
C6318 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 3.84e-20
C6319 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 2.49e-20
C6320 CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0263f
C6321 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_0.OUT a_25490_n1899# 0.0203f
C6322 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 0.00998f
C6323 F1 Vdiv99 9.46e-19
C6324 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 2.19e-20
C6325 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 7.98e-20
C6326 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_48832_n1102# 0.00118f
C6327 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00156f
C6328 VDD90 a_25312_5018# 0.0123f
C6329 VDD96 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 1.24f
C6330 a_54022_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0203f
C6331 VDD90 dec3x8_ibr_mag_0.and_3_ibr_1.nand3_mag_ibr_0.OUT 0.0267f
C6332 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_29053_5018# 9.1e-19
C6333 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 0.0172f
C6334 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K a_31177_7256# 0.0027f
C6335 RST a_23703_n287# 0.00102f
C6336 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K 2.32f
C6337 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0622f
C6338 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 0.065f
C6339 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_50287_n18696# 0.00111f
C6340 RST CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.0239f
C6341 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.792f
C6342 a_48023_n7840# CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 0.00263f
C6343 CLK CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 1.29e-19
C6344 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 4.07e-19
C6345 a_25529_n743# CLK_div_96_mag_0.JK_FF_mag_0.Q 3.87e-20
C6346 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 0.00761f
C6347 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 8.26e-20
C6348 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB 1.97f
C6349 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 6.87e-20
C6350 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_45131_n17599# 0.0101f
C6351 CLK_div_108_new_mag_0.JK_FF_mag_1.QB a_51393_n6821# 0.00964f
C6352 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 a_51604_10154# 0.00166f
C6353 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_55357_n20487# 5.39e-20
C6354 RST CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 4.25e-20
C6355 a_53813_n6862# CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 1.8e-21
C6356 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 0.209f
C6357 RST a_37237_n8887# 8.63e-19
C6358 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.00488f
C6359 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.507f
C6360 VDD105 a_49752_10154# 0.00152f
C6361 dec3x8_ibr_mag_0.and_3_ibr_6.nand3_mag_ibr_0.OUT a_39420_6265# 6.08e-20
C6362 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 3.28e-19
C6363 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.12f
C6364 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 3.34e-21
C6365 RST a_32295_n16632# 0.00206f
C6366 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 3.79e-20
C6367 dec3x8_ibr_mag_0.and_3_ibr_1.nand3_mag_ibr_0.OUT a_38454_6821# 3.58e-20
C6368 VDD108 a_54658_n9064# 6.01e-19
C6369 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 2.11e-19
C6370 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.0838f
C6371 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 0.25f
C6372 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.233f
C6373 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_96_mag_0.JK_FF_mag_2.Q 7.24e-19
C6374 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.00975f
C6375 a_31571_n16632# a_31731_n16632# 0.0504f
C6376 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_28623_n15537# 1.24e-20
C6377 CLK a_25364_n19822# 2.29e-19
C6378 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 a_37999_n1222# 0.00372f
C6379 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 0.0871f
C6380 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_54033_n15587# 1.43e-19
C6381 CLK CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 1.22e-19
C6382 RST a_25686_1919# 5.97e-19
C6383 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT a_26183_n7107# 0.0732f
C6384 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.0675f
C6385 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 0.0151f
C6386 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K a_50917_n9020# 1.75e-19
C6387 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_22718_8532# 1.4e-19
C6388 CLK a_31128_n7028# 2.43e-19
C6389 RST CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.VOUT 0.0494f
C6390 RST a_53934_n9020# 2.23e-19
C6391 F0 a_38454_6265# 8.64e-19
C6392 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_53939_1671# 0.00378f
C6393 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 0.00761f
C6394 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_23403_10099# 0.00378f
C6395 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 0.0598f
C6396 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_50310_n15627# 0.00392f
C6397 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_47810_5143# 0.0203f
C6398 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT 0.00183f
C6399 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_51028_n16724# 0.00696f
C6400 CLK_div_96_mag_0.JK_FF_mag_3.QB CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.103f
C6401 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_48092_n9063# 0.0732f
C6402 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.225f
C6403 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 0.0022f
C6404 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 a_25472_5018# 0.00789f
C6405 RST a_22988_n1789# 0.0013f
C6406 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 a_45927_6284# 8.17e-21
C6407 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 6.22e-20
C6408 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.311f
C6409 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_27381_n699# 0.0811f
C6410 a_45131_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.00696f
C6411 VDD105 a_44075_6240# 0.00752f
C6412 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 1.87e-19
C6413 VDD105 a_46081_5187# 0.00152f
C6414 CLK CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 0.00249f
C6415 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C6416 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0622f
C6417 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 1.41e-20
C6418 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.109f
C6419 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0635f
C6420 VDD108 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.391f
C6421 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_28099_n17626# 0.0203f
C6422 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.00942f
C6423 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 0.23f
C6424 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB 7.08e-20
C6425 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 0.0501f
C6426 VDD93 a_40254_n8887# 3.14e-19
C6427 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 0.00118f
C6428 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 0.768f
C6429 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.0635f
C6430 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 a_51729_n17599# 0.069f
C6431 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT a_53216_n10117# 0.00378f
C6432 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 a_48783_n13424# 0.00107f
C6433 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.652f
C6434 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 a_31128_n7028# 0.00347f
C6435 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.00488f
C6436 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_29307_n1855# 1.43e-19
C6437 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.26f
C6438 RST a_31445_n18723# 3.71e-19
C6439 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 5.73e-20
C6440 a_30164_n7017# CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.069f
C6441 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_25082_n17626# 9.1e-19
C6442 RST a_35032_n17626# 5.2e-19
C6443 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 0.878f
C6444 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_47338_n6273# 0.00378f
C6445 a_22011_n287# CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 2.73e-19
C6446 a_26820_3016# a_26980_3016# 0.0504f
C6447 Vdiv105 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT 8.87e-20
C6448 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.00205f
C6449 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.322f
C6450 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 a_30435_n1855# 1.63e-20
C6451 CLK a_32015_n17626# 0.00164f
C6452 RST CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.00543f
C6453 a_22264_n1833# a_22424_n1833# 0.0504f
C6454 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.0635f
C6455 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 9.69e-19
C6456 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 1.05e-19
C6457 RST a_44793_5143# 8.64e-19
C6458 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 8.28e-20
C6459 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_51961_6284# 0.00118f
C6460 VDD108 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.399f
C6461 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_44061_n15627# 0.00119f
C6462 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 0.69f
C6463 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 a_53934_n9020# 1.43e-19
C6464 VDD93 a_26226_n9831# 3.14e-19
C6465 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.365f
C6466 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.211f
C6467 a_53303_n16728# a_53463_n16728# 0.0504f
C6468 CLK CLK_div_99_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.102f
C6469 CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 8.07e-21
C6470 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN 0.108f
C6471 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_39844_n10028# 0.0733f
C6472 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT a_50204_2768# 0.00378f
C6473 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00943f
C6474 a_50829_n6865# CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 8.31e-21
C6475 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB a_24901_n6010# 0.00964f
C6476 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 1.58e-20
C6477 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 a_22551_n14504# 4.15e-19
C6478 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 1.48e-19
C6479 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 0.655f
C6480 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 9.62e-20
C6481 VDD mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.46f
C6482 Vdiv99 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.IN1 0.0241f
C6483 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 a_47453_9057# 0.0059f
C6484 RST a_49635_n10117# 0.00114f
C6485 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 1.84e-19
C6486 RST CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.101f
C6487 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_39844_n10028# 2.88e-20
C6488 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.0592f
C6489 VDD99 a_35192_n17626# 0.0132f
C6490 RST CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.0834f
C6491 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.258f
C6492 Vdiv90 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT 0.243f
C6493 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 a_30727_n17626# 0.00859f
C6494 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 6.91e-20
C6495 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_26990_11196# 1.46e-19
C6496 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN a_25488_n15535# 1.03e-20
C6497 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT a_53463_n16728# 0.0731f
C6498 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_51285_n1102# 0.011f
C6499 CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 3.15e-20
C6500 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K a_48324_n15585# 3.47e-19
C6501 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0702f
C6502 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 1.18f
C6503 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 2.62e-19
C6504 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 a_22455_5018# 0.00789f
C6505 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 0.0404f
C6506 CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 a_39120_n10028# 0.00789f
C6507 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K a_50144_n16724# 8.64e-19
C6508 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 a_29905_n16590# 0.069f
C6509 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00183f
C6510 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.107f
C6511 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.16f
C6512 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 a_51592_n16680# 0.069f
C6513 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_50103_5143# 0.0202f
C6514 a_46768_n5176# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.46e-19
C6515 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.0215f
C6516 CLK a_24337_n6010# 0.00178f
C6517 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 a_29270_n743# 0.0101f
C6518 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 8.4e-19
C6519 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_22461_6115# 0.00119f
C6520 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.996f
C6521 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN 0.107f
C6522 a_29708_n8735# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 4.52e-20
C6523 VDD VDD96 0.487f
C6524 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN a_48783_n13424# 4.43e-21
C6525 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 6.18e-19
C6526 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 1.08f
C6527 VDD93 a_37955_n9984# 0.00149f
C6528 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.642f
C6529 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_45075_n9063# 0.0732f
C6530 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.225f
C6531 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.338f
C6532 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_45452_1671# 0.00486f
C6533 CLK a_33898_n18723# 6.06e-21
C6534 VDD mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I1 0.423f
C6535 Vdiv108 a_49991_n2243# 0.00158f
C6536 VDD100 Vdiv100 0.126f
C6537 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_47196_n15629# 2.79e-20
C6538 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 0.392f
C6539 RST a_47332_n5176# 0.00172f
C6540 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_47492_n5176# 2.88e-20
C6541 CLK_div_90_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_33245_7558# 9.16e-20
C6542 a_26226_n9831# m3_20882_n11188# 2.84e-19
C6543 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_48478_n16682# 0.00859f
C6544 CLK CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 5.57e-19
C6545 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_48324_n15585# 2.96e-19
C6546 a_34308_n17626# a_34468_n17626# 0.0504f
C6547 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_22565_n6009# 0.0203f
C6548 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 7.24e-19
C6549 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.1f
C6550 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.00668f
C6551 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 0.00975f
C6552 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 2.59e-21
C6553 RST CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.261f
C6554 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 1.66f
C6555 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.00157f
C6556 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 m3_20882_n11188# 0.00156f
C6557 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 a_45753_n15583# 0.00372f
C6558 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 2.87e-19
C6559 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT a_50763_n10161# 0.0733f
C6560 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.JK_FF_mag_0.QB 2.26e-19
C6561 a_44069_5143# a_44229_5143# 0.0504f
C6562 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 a_48741_9057# 0.0101f
C6563 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 a_21902_n8787# 0.00939f
C6564 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_46974_n2243# 0.0202f
C6565 CLK a_28329_5018# 0.00134f
C6566 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_32301_n15491# 1.43e-19
C6567 VDD96 a_26974_1919# 0.00533f
C6568 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0683f
C6569 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT 0.32f
C6570 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 1f
C6571 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_50103_5143# 1.17e-20
C6572 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_48944_6284# 0.00118f
C6573 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 a_50917_n9020# 1.43e-19
C6574 VDD100 a_43957_n2243# 0.0132f
C6575 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 8.16e-20
C6576 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_29623_6159# 7.4e-19
C6577 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN 0.012f
C6578 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 0.0881f
C6579 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_22258_n2930# 0.0202f
C6580 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.122f
C6581 a_37955_n9984# m3_20882_n11188# 3.71e-19
C6582 VDD96 a_25490_n1899# 0.00533f
C6583 CLK_div_96_mag_0.JK_FF_mag_5.Q CLK_div_96_mag_0.JK_FF_mag_0.QB 0.308f
C6584 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.00975f
C6585 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB a_46810_n10116# 0.00964f
C6586 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.122f
C6587 CLK_div_90_mag_0.CLK_div_10_mag_0.CLK a_22295_5018# 0.00117f
C6588 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_24153_6159# 0.00372f
C6589 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 0.397f
C6590 CLK_div_108_new_mag_0.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K 5.25e-20
C6591 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_36178_n16592# 0.0036f
C6592 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_39126_n8931# 0.00392f
C6593 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB a_45612_1671# 1.86e-20
C6594 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT 0.233f
C6595 a_48098_n10160# a_48258_n10160# 0.0504f
C6596 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 a_51165_n17599# 3.66e-20
C6597 VDD mux_8x1_ibr_0.mux_2x1_ibr_0.I0 1.44f
C6598 mux_8x1_ibr_0.mux_2x1_ibr_0.I1 Vdiv108 0.00509f
C6599 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00164f
C6600 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.233f
C6601 VDD90 a_24307_5062# 0.00152f
C6602 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_48268_n1102# 0.011f
C6603 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 1.32e-19
C6604 a_53458_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 1.5e-20
C6605 a_54022_n17599# a_54182_n17599# 0.0504f
C6606 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 2.34e-19
C6607 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0135f
C6608 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.0591f
C6609 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.121f
C6610 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_28489_5018# 0.0731f
C6611 RST a_48635_2768# 0.00186f
C6612 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 1.96f
C6613 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 0.16f
C6614 RST a_23139_n287# 0.00248f
C6615 VDD100 dec3x8_ibr_mag_0.and_3_ibr_3.nand3_mag_ibr_0.OUT 0.0367f
C6616 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.398f
C6617 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_49122_n18696# 7.4e-19
C6618 VDD100 a_51871_n5# 3.14e-19
C6619 CLK_div_96_mag_0.JK_FF_mag_0.QB a_24270_n2886# 0.0811f
C6620 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.16f
C6621 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0225f
C6622 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 0.397f
C6623 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0048f
C6624 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0635f
C6625 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.305f
C6626 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.36f
C6627 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT 0.664f
C6628 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.304f
C6629 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 4.52e-20
C6630 Vdiv105 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 1.08e-19
C6631 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_44971_n17599# 0.0102f
C6632 CLK_div_108_new_mag_0.JK_FF_mag_1.QB a_50829_n6865# 0.00696f
C6633 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 a_51040_10154# 3.6e-22
C6634 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_55197_n20487# 9.16e-20
C6635 RST a_36673_n8887# 2.23e-19
C6636 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT 1.19f
C6637 VDD96 CLK_div_96_mag_0.JK_FF_mag_2.Q 2.13f
C6638 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK a_50105_n6865# 0.00233f
C6639 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0706f
C6640 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_96_mag_0.JK_FF_mag_2.QB 6.48e-19
C6641 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 6.43e-20
C6642 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 9.46e-19
C6643 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 a_29213_n7028# 0.00347f
C6644 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 0.00265f
C6645 RST a_31731_n16632# 0.00273f
C6646 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00639f
C6647 dec3x8_ibr_mag_0.and_3_ibr_1.nand3_mag_ibr_0.OUT a_38294_6821# 6.08e-20
C6648 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.16f
C6649 VDD108 a_54498_n9064# 2.65e-19
C6650 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 0.395f
C6651 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 a_28268_n6266# 0.00665f
C6652 a_28267_n7033# CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.069f
C6653 VDD dec3x8_ibr_mag_0.and_3_ibr_3.IN1 1.73f
C6654 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.121f
C6655 VDD108 a_50669_n6865# 2.21e-19
C6656 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.0758f
C6657 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_28463_n15537# 1.59e-20
C6658 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C6659 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_50987_5143# 8.64e-19
C6660 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00156f
C6661 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C6662 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.399f
C6663 F1 a_37999_n1222# 2.62e-19
C6664 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.314f
C6665 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.16f
C6666 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_53469_n15631# 0.00119f
C6667 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT 0.298f
C6668 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.338f
C6669 RST a_25122_1919# 5.97e-19
C6670 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT a_25619_n7107# 0.00378f
C6671 Vdiv110 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT 0.00876f
C6672 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 F1 3.02e-20
C6673 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K a_50353_n9020# 2.96e-19
C6674 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 0.00975f
C6675 RST a_53370_n9020# 0.00121f
C6676 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 5.32e-19
C6677 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_5.QB 0.248f
C6678 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0201f
C6679 F0 a_38294_6265# 0.00181f
C6680 Vdiv108 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0343f
C6681 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 0.00586f
C6682 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.103f
C6683 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 0.00975f
C6684 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_47246_5143# 1.5e-20
C6685 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 0.399f
C6686 VDD99 a_32295_n16632# 2.77e-19
C6687 a_33359_11196# a_33519_11196# 0.0504f
C6688 RST CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.00738f
C6689 CLK_div_108_new_mag_0.JK_FF_mag_1.QB CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.198f
C6690 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_50868_n16724# 0.00695f
C6691 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_47528_n9019# 0.00378f
C6692 CLK_div_90_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 3.87e-19
C6693 RST a_26980_3016# 0.00195f
C6694 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 0.329f
C6695 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 a_25312_5018# 0.00335f
C6696 RST a_22424_n1833# 9.48e-19
C6697 Vdiv100 CLK_div_100_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 0.0289f
C6698 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.647f
C6699 CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 a_40818_n8887# 0.069f
C6700 RST CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.193f
C6701 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C6702 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_26817_n699# 0.00964f
C6703 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 0.122f
C6704 RST a_51034_9057# 1.23e-20
C6705 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_45695_n17599# 0.00378f
C6706 a_44971_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.00695f
C6707 a_46608_n5176# a_46768_n5176# 0.0504f
C6708 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN 0.125f
C6709 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT a_50874_n15583# 0.00378f
C6710 VDD105 a_45517_5187# 0.00152f
C6711 a_26253_n743# CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 3.87e-20
C6712 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 a_51652_2768# 0.00335f
C6713 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_27939_n17626# 0.0733f
C6714 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 3.28e-19
C6715 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 8.04e-19
C6716 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.00111f
C6717 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 0.119f
C6718 VDD93 a_39690_n8887# 3.14e-19
C6719 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 a_50903_n5# 0.00929f
C6720 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.25f
C6721 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0501f
C6722 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 a_48623_n13424# 0.00271f
C6723 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.397f
C6724 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 0.0437f
C6725 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.289f
C6726 RST a_30881_n18723# 3.96e-19
C6727 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_28743_n1899# 0.00119f
C6728 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 0.00935f
C6729 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0622f
C6730 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 0.00188f
C6731 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_24922_n17626# 2.88e-20
C6732 RST a_34468_n17626# 0.00108f
C6733 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.652f
C6734 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.652f
C6735 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.0854f
C6736 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.321f
C6737 F2 Vdiv100 0.00618f
C6738 CLK_div_105_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 4.42e-19
C6739 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0622f
C6740 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB 0.311f
C6741 F0 Vdiv110 0.534f
C6742 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 7.98e-19
C6743 a_29801_1733# CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.00168f
C6744 VDD108 a_50199_n10117# 3.14e-19
C6745 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN 4.36e-20
C6746 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_51397_6284# 0.011f
C6747 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB 0.103f
C6748 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 a_53370_n9020# 0.011f
C6749 VDD108 Vdiv100 0.11f
C6750 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 0.0224f
C6751 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_25420_n13385# 0.0131f
C6752 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_45343_n16680# 0.0036f
C6753 CLK a_24391_n20290# 0.00132f
C6754 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 8.16e-20
C6755 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN a_30244_398# 4.94e-20
C6756 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT a_37436_880# 9.43e-19
C6757 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_39684_n10028# 0.0203f
C6758 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK a_47196_n15629# 1.88e-19
C6759 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 a_55161_n15587# 0.00372f
C6760 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.231f
C6761 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB a_24337_n6010# 0.0811f
C6762 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN a_47723_574# 0.069f
C6763 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.103f
C6764 a_23956_n14213# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 3.01e-20
C6765 RST a_48258_n10160# 0.00218f
C6766 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00637f
C6767 VDD99 a_31445_n18723# 3.14e-19
C6768 Vdiv93 CLK_div_93_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 1.39e-19
C6769 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_39684_n10028# 9.1e-19
C6770 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0018f
C6771 VDD99 a_35032_n17626# 0.00888f
C6772 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 a_30163_n17626# 0.0157f
C6773 RST a_54182_n17599# 0.00154f
C6774 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 1.36e-19
C6775 VDD99 a_36588_n15495# 3.56e-19
C6776 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.11f
C6777 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 1.08f
C6778 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN a_25328_n15535# 1.29e-20
C6779 a_55156_n18696# CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 1.54e-19
C6780 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT a_53303_n16728# 0.0202f
C6781 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.00157f
C6782 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_50721_n1102# 1.43e-19
C6783 a_28386_n743# CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 9.14e-19
C6784 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 a_22295_5018# 0.00335f
C6785 CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 a_38960_n10028# 0.00335f
C6786 VDD93 dec3x8_ibr_mag_0.and_3_ibr_1.nand3_mag_ibr_0.OUT 6.58e-19
C6787 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 0.00975f
C6788 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.24f
C6789 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 a_29110_n743# 0.0102f
C6790 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.343f
C6791 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.283f
C6792 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 1.54e-21
C6793 CLK_div_108_new_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 3.34e-19
C6794 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB 0.28f
C6795 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.0635f
C6796 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_42529_n14305# 0.00379f
C6797 Vdiv110 m3_20882_n11188# 0.0163f
C6798 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 8.58e-20
C6799 dec3x8_ibr_mag_0.and_3_ibr_1.nand3_mag_ibr_0.OUT F0 0.00225f
C6800 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN a_48623_n13424# 3.44e-21
C6801 VDD99 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.99e-19
C6802 VDD93 a_37391_n9984# 0.00149f
C6803 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.802f
C6804 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_44511_n9019# 0.00378f
C6805 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 0.00178f
C6806 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 0.231f
C6807 VDD a_37168_6265# 2.21e-19
C6808 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0622f
C6809 a_22295_5018# a_22455_5018# 0.0504f
C6810 CLK a_33334_n18723# 9.45e-19
C6811 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_44888_1671# 3.25e-19
C6812 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.0784f
C6813 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 8.39e-21
C6814 Vdiv108 a_48986_n2199# 7.51e-19
C6815 RST a_46768_n5176# 0.00345f
C6816 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_47332_n5176# 9.1e-19
C6817 VDD mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_1.IN2 0.456f
C6818 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 0.122f
C6819 CLK a_30502_11196# 0.00117f
C6820 a_25662_n9875# m3_20882_n11188# 2.88e-19
C6821 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_47914_n16726# 0.0101f
C6822 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.0228f
C6823 CLK_div_105_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.144f
C6824 RST CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0677f
C6825 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 0.00158f
C6826 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_51393_n6821# 0.00378f
C6827 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_47760_n15585# 3.12e-19
C6828 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 1.09e-20
C6829 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.0718f
C6830 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 7.08e-20
C6831 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_22405_n6009# 0.0733f
C6832 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0352f
C6833 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_49042_n16682# 0.0811f
C6834 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 0.00335f
C6835 a_25646_n17626# a_25806_n17626# 0.0504f
C6836 F2 dec3x8_ibr_mag_0.and_3_ibr_3.nand3_mag_ibr_0.OUT 0.111f
C6837 VDD110 a_55310_n17599# 3.14e-19
C6838 VDD99 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 0.161f
C6839 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT 0.233f
C6840 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 0.116f
C6841 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 a_45189_n15583# 0.069f
C6842 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 0.122f
C6843 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 0.215f
C6844 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 4.36e-20
C6845 a_29110_n743# a_29270_n743# 0.0504f
C6846 VDD108 dec3x8_ibr_mag_0.and_3_ibr_3.nand3_mag_ibr_0.OUT 0.154f
C6847 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT a_50199_n10117# 0.00378f
C6848 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 2.71e-21
C6849 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 0.397f
C6850 Vdiv99 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.245f
C6851 CLK_div_96_mag_0.JK_FF_mag_2.QB CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 2.53e-20
C6852 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C6853 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB a_50928_2768# 0.00695f
C6854 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 2.51e-19
C6855 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 a_48581_9057# 0.00939f
C6856 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_53973_n6862# 2.88e-20
C6857 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 a_21742_n8787# 0.0101f
C6858 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 0.0128f
C6859 CLK a_27324_5062# 6.21e-19
C6860 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I1 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.11f
C6861 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_31737_n15535# 0.00119f
C6862 a_23709_810# a_23869_810# 0.0504f
C6863 VDD110 a_51165_n17599# 0.00101f
C6864 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0569f
C6865 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 1.17e-19
C6866 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_48380_6284# 0.011f
C6867 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 a_50353_n9020# 0.011f
C6868 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.311f
C6869 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.235f
C6870 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C6871 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB a_23594_n8743# 0.0114f
C6872 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_29059_6159# 3.12e-19
C6873 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.0615f
C6874 CLK CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.00118f
C6875 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT a_33652_n13270# 8.09e-22
C6876 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB 0.144f
C6877 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_96_mag_0.JK_FF_mag_0.Q 0.107f
C6878 a_37391_n9984# m3_20882_n11188# 3.57e-19
C6879 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.121f
C6880 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 1.49e-21
C6881 VDD96 a_24116_n1789# 3.76e-19
C6882 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB a_46246_n10116# 0.0811f
C6883 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.359f
C6884 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_23589_6159# 0.069f
C6885 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.391f
C6886 CLK CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT 0.235f
C6887 RST CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN 0.0411f
C6888 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB a_45452_1671# 1.41e-20
C6889 RST CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.0495f
C6890 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0343f
C6891 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_53249_n6862# 1.46e-19
C6892 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 4.46e-20
C6893 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 a_21995_n7106# 0.069f
C6894 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 9.38e-20
C6895 VDD90 a_23743_5062# 0.00152f
C6896 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_47704_n1102# 1.43e-19
C6897 a_53298_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 1.17e-20
C6898 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_28329_5018# 0.0202f
C6899 RST a_48475_2768# 0.00186f
C6900 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT a_54664_n10161# 0.0202f
C6901 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 CLK_div_99_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 8.04e-19
C6902 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_31661_10099# 4.52e-20
C6903 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.0854f
C6904 RST a_22575_n287# 0.001f
C6905 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 0.029f
C6906 RST CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0175f
C6907 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_48558_n18696# 7.4e-19
C6908 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.0592f
C6909 CLK_div_96_mag_0.JK_FF_mag_0.QB a_23706_n2886# 0.00964f
C6910 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 8.33e-20
C6911 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 6.04e-20
C6912 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 9.89e-20
C6913 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 3.61e-20
C6914 F0 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT 2.41e-19
C6915 VDD100 a_48629_1671# 0.00746f
C6916 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_53129_n19793# 0.0096f
C6917 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 3.67e-20
C6918 RST CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 0.166f
C6919 F0 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT 5.24e-19
C6920 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 0.116f
C6921 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.104f
C6922 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.179f
C6923 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_44407_n17599# 0.00789f
C6924 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 3.56e-19
C6925 CLK_div_108_new_mag_0.JK_FF_mag_1.QB a_50669_n6865# 0.00695f
C6926 a_35949_n8931# a_36109_n8931# 0.0504f
C6927 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK a_49945_n6865# 0.00211f
C6928 RST a_36109_n8931# 6.43e-19
C6929 CLK CLK_div_100_mag_0.CLK_div_10_mag_1.CLK 1.22e-19
C6930 CLK_div_100_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 1.29e-19
C6931 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.00139f
C6932 RST CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.193f
C6933 RST a_31571_n16632# 0.00273f
C6934 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_2.Q 0.00335f
C6935 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_29905_n16590# 0.0036f
C6936 CLK_div_96_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.00384f
C6937 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 0.0165f
C6938 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 a_33429_n15491# 0.00372f
C6939 VDD108 a_53934_n9020# 3.16e-19
C6940 VDD100 a_48635_2768# 0.0132f
C6941 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 0.00178f
C6942 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 2.48e-19
C6943 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_27180_n15491# 0.0114f
C6944 a_52161_n19793# CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.00138f
C6945 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 7.38e-19
C6946 VDD105 a_51758_9057# 3.78e-19
C6947 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN 1.54e-19
C6948 F1 a_36873_n1222# 2.15e-19
C6949 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.0854f
C6950 a_54621_10154# a_54781_10154# 0.0504f
C6951 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 a_30164_n7017# 0.0193f
C6952 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 5.26e-19
C6953 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT 0.00168f
C6954 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 1.45e-19
C6955 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_53463_n16728# 1.46e-19
C6956 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.046f
C6957 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K a_49789_n9020# 0.012f
C6958 RST a_52806_n9020# 0.00154f
C6959 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 1.18f
C6960 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 8.59e-20
C6961 RST CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 0.118f
C6962 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 3.67e-20
C6963 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_47086_5143# 1.17e-20
C6964 RST a_30164_n7017# 2.96e-19
C6965 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 1.86e-19
C6966 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.121f
C6967 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB 0.0384f
C6968 RST a_26820_3016# 0.00195f
C6969 RST a_22264_n1833# 8.86e-19
C6970 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 0.053f
C6971 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 0.0854f
C6972 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB 0.915f
C6973 CLK CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00147f
C6974 a_44436_9057# CLK_div_105_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 5.94e-20
C6975 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_26253_n743# 0.00696f
C6976 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K a_45899_7960# 0.0027f
C6977 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT a_50310_n15627# 0.0732f
C6978 VDD105 a_44953_5143# 0.00101f
C6979 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.92f
C6980 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_27375_n17626# 0.00378f
C6981 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 a_51492_2768# 0.00789f
C6982 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 2.33e-19
C6983 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.00174f
C6984 CLK_div_100_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.144f
C6985 a_25484_n2996# a_25644_n2996# 0.0504f
C6986 CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 0.149f
C6987 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 0.231f
C6988 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 a_48944_6284# 9.26e-19
C6989 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.395f
C6990 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0228f
C6991 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 4.54f
C6992 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 1.06e-19
C6993 VDD99 a_26980_3016# 0.00244f
C6994 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 4.33e-20
C6995 a_53973_n6862# CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT 1.8e-21
C6996 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 0.25f
C6997 RST a_30317_n18723# 3.96e-19
C6998 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 1.61e-19
C6999 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.36f
C7000 RST a_34308_n17626# 0.00173f
C7001 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_50447_n18696# 0.00119f
C7002 RST a_35460_n15495# 2.67e-19
C7003 CLK Vdiv108 0.00437f
C7004 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 3.23e-20
C7005 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT Vdiv100 0.244f
C7006 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 8.93e-21
C7007 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 8.36e-19
C7008 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00183f
C7009 VDD108 a_49635_n10117# 3.14e-19
C7010 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 a_23289_n6009# 0.0122f
C7011 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB 0.0381f
C7012 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.121f
C7013 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 9.52e-19
C7014 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C7015 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.768f
C7016 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN 0.00126f
C7017 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_50833_6284# 1.43e-19
C7018 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 a_52806_n9020# 0.00118f
C7019 VDD93 a_25502_n9875# 2.21e-19
C7020 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_24358_n17626# 0.069f
C7021 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT a_36873_880# 0.00949f
C7022 a_51015_7381# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 2.36e-22
C7023 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_39120_n10028# 1.5e-20
C7024 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK a_47036_n15629# 2.69e-19
C7025 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 a_54597_n15587# 0.069f
C7026 a_53732_n2243# a_53892_n2243# 0.0504f
C7027 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB 0.198f
C7028 F2 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 0.443f
C7029 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 4.1e-21
C7030 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0894f
C7031 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0231f
C7032 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.429f
C7033 RST a_48098_n10160# 0.00218f
C7034 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.321f
C7035 VDD99 a_30881_n18723# 3.14e-19
C7036 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_39120_n10028# 0.0731f
C7037 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.402f
C7038 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB m3_20882_n11188# 0.00361f
C7039 dec3x8_ibr_mag_0.and_3_ibr_2.nand3_mag_ibr_0.OUT dec3x8_ibr_mag_0.and_3_ibr_6.nand3_mag_ibr_0.OUT 0.00141f
C7040 RST a_54022_n17599# 0.00195f
C7041 VDD99 a_34468_n17626# 0.0012f
C7042 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.321f
C7043 VDD99 a_36024_n15495# 3.14e-19
C7044 RST CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 0.117f
C7045 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 a_31352_6115# 6.36e-19
C7046 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 1.79e-19
C7047 a_51961_6284# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 4.52e-20
C7048 CLK_div_96_mag_0.JK_FF_mag_5.Q CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 9.24e-19
C7049 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_47970_5143# 8.64e-19
C7050 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_50157_n1146# 0.00119f
C7051 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00101f
C7052 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K 1.22e-23
C7053 CLK_div_105_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 3.38e-19
C7054 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 9.73e-19
C7055 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 0.00216f
C7056 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 a_25640_n18723# 2.79e-20
C7057 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_30398_n699# 0.0811f
C7058 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.69f
C7059 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.28f
C7060 VDD108 a_47332_n5176# 2.21e-19
C7061 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 a_28546_n743# 0.00707f
C7062 Vdiv110 m1_42708_4265# 0.00151f
C7063 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0622f
C7064 VDD96 a_23863_n287# 0.00536f
C7065 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 0.026f
C7066 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_25640_n18723# 0.00119f
C7067 a_45603_n5176# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.0811f
C7068 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.00157f
C7069 VDD93 a_36827_n10028# 9.82e-19
C7070 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 9.9e-19
C7071 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 3.98e-20
C7072 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 6.69e-19
C7073 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_44324_1671# 2.96e-19
C7074 VDD110 Vdiv108 0.779f
C7075 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 6.88e-21
C7076 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 a_52839_n5# 0.0096f
C7077 Vdiv108 a_48422_n2199# 7.3e-19
C7078 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 0.0034f
C7079 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 7.81e-19
C7080 RST a_46608_n5176# 0.00345f
C7081 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_46768_n5176# 0.0731f
C7082 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0343f
C7083 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_47754_n16726# 0.0102f
C7084 CLK a_30342_11196# 0.00164f
C7085 a_25502_n9875# m3_20882_n11188# 2.88e-19
C7086 F1 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 0.00223f
C7087 CLK_div_96_mag_0.JK_FF_mag_4.QB CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_0.OUT 0.343f
C7088 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_50829_n6865# 0.0733f
C7089 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 6.36e-20
C7090 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_47196_n15629# 0.00392f
C7091 CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 a_54866_n1102# 0.069f
C7092 VDD100 Vdiv 0.192f
C7093 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_21841_n6009# 0.00378f
C7094 VDD105 dec3x8_ibr_mag_0.and_3_ibr_3.nand3_mag_ibr_0.OUT 7.15e-19
C7095 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.487f
C7096 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_48478_n16682# 0.00964f
C7097 VDD96 CLK_div_96_mag_0.JK_FF_mag_3.QB 0.902f
C7098 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.0515f
C7099 F2 a_36202_6821# 3.45e-20
C7100 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0636f
C7101 VDD110 a_54746_n17599# 3.14e-19
C7102 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_30496_10099# 0.0203f
C7103 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.00131f
C7104 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.363f
C7105 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.877f
C7106 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 0.0591f
C7107 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 1.08f
C7108 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.00166f
C7109 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB a_50768_2768# 0.00696f
C7110 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 5.7f
C7111 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB 1.22e-19
C7112 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 0.28f
C7113 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.321f
C7114 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.00335f
C7115 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 a_48017_9057# 1.25e-20
C7116 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_53813_n6862# 9.1e-19
C7117 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.649f
C7118 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C7119 CLK a_26760_5062# 6.02e-19
C7120 a_26250_1919# CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 3.53e-20
C7121 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 1.01f
C7122 VDD96 a_26250_1919# 3.14e-19
C7123 VDD110 a_51005_n17599# 0.00123f
C7124 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.00396f
C7125 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT a_51015_7381# 7.43e-22
C7126 Vdiv90 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT 2.68e-19
C7127 CLK_div_96_mag_0.JK_FF_mag_4.Q a_23869_810# 0.0022f
C7128 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_47816_6284# 1.43e-19
C7129 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_32635_11196# 8.64e-19
C7130 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_27150_11196# 1.17e-20
C7131 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 a_49789_n9020# 0.00118f
C7132 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 a_24491_n7107# 4.52e-20
C7133 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.089f
C7134 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 a_26636_n8734# 0.069f
C7135 VDD96 CLK_div_90_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 0.00215f
C7136 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.00518f
C7137 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB a_23030_n8743# 2.96e-19
C7138 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK 2.14e-20
C7139 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_28495_6115# 9.32e-19
C7140 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.338f
C7141 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 a_51849_n1102# 0.00372f
C7142 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00229f
C7143 RST a_47905_1671# 1.23e-20
C7144 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT a_30915_n13291# 2.05e-19
C7145 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB 0.0312f
C7146 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00183f
C7147 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.122f
C7148 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.159f
C7149 a_36827_n10028# m3_20882_n11188# 3.55e-19
C7150 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_4.Q 0.00358f
C7151 VDD96 a_23552_n1789# 3.19e-19
C7152 RST CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 0.158f
C7153 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 1.93e-20
C7154 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0894f
C7155 RST a_26636_n8734# 0.00126f
C7156 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT 0.0693f
C7157 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 6.63e-19
C7158 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_48148_n17599# 0.0101f
C7159 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT a_31177_7256# 3.92e-20
C7160 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 a_21431_n7106# 0.00372f
C7161 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 1.96f
C7162 VDD90 a_23179_5018# 0.00101f
C7163 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_47140_n1146# 0.00119f
C7164 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 0.11f
C7165 CLK_div_96_mag_0.JK_FF_mag_5.Q a_23869_810# 0.00335f
C7166 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 0.21f
C7167 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT a_54504_n10161# 0.0731f
C7168 RST a_47911_2768# 0.00169f
C7169 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN a_52951_7381# 0.069f
C7170 RST CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.177f
C7171 RST a_22011_n287# 4.11e-19
C7172 Vdiv110 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.119f
C7173 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB a_51758_9057# 1.86e-20
C7174 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 9.52e-19
C7175 RST a_28734_n9876# 0.00147f
C7176 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_47994_n18696# 3.12e-19
C7177 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB m3_20882_n11188# 0.00346f
C7178 CLK_div_96_mag_0.JK_FF_mag_0.QB a_23142_n2930# 0.00696f
C7179 RST CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 0.33f
C7180 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 7.43e-20
C7181 CLK_div_108_new_mag_0.JK_FF_mag_1.Q CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.267f
C7182 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 5.32e-21
C7183 CLK CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 1.8e-19
C7184 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.IN1 1.2e-19
C7185 VDD100 a_48469_1671# 2.66e-19
C7186 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.0206f
C7187 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT 0.163f
C7188 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 2.39e-19
C7189 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.392f
C7190 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB 0.92f
C7191 VDD99 a_22551_n14504# 2.21e-19
C7192 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB 0.106f
C7193 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.233f
C7194 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 1.22f
C7195 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_45251_n1102# 4.52e-20
C7196 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_44247_n17599# 0.00335f
C7197 VDD99 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 1.08e-20
C7198 CLK CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00511f
C7199 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 0.205f
C7200 CLK_div_108_new_mag_0.CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN a_51205_n7921# 0.069f
C7201 CLK CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 7.15e-19
C7202 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00118f
C7203 a_24153_6159# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 4.52e-20
C7204 RST a_35949_n8931# 7.78e-19
C7205 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.298f
C7206 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 a_40375_n7552# 6.83e-19
C7207 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 4.52e-20
C7208 CLK_div_90_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_32640_6159# 5.94e-20
C7209 RST a_30469_n16590# 0.00137f
C7210 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.013f
C7211 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.0432f
C7212 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 a_32865_n15491# 0.069f
C7213 RST CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.207f
C7214 VDD100 a_48475_2768# 0.00891f
C7215 VDD108 a_53370_n9020# 3.16e-19
C7216 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB 0.0838f
C7217 F2 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 0.366f
C7218 VDD108 a_49945_n6865# 0.00108f
C7219 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_29461_n2996# 8.64e-19
C7220 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_26616_n15491# 2.96e-19
C7221 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00148f
C7222 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 7.33e-20
C7223 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_5.Q 0.00383f
C7224 VDD105 a_51598_9057# 2.66e-19
C7225 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 6.32e-22
C7226 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_33519_11196# 0.0202f
C7227 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN 0.519f
C7228 CLK CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00131f
C7229 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_110_mag_0.CLK_div_10_mag_0.CLK 0.0212f
C7230 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_47430_n18696# 0.00119f
C7231 Vdiv108 a_55101_n6818# 0.0157f
C7232 VDD93 Vdiv99 0.634f
C7233 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.911f
C7234 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 5.37e-19
C7235 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K a_48252_n9063# 1.01e-20
C7236 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K 0.00102f
C7237 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN 0.0103f
C7238 RST a_51641_n9064# 0.00214f
C7239 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 0.104f
C7240 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.0175f
C7241 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT 0.00183f
C7242 VDD99 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 1.08e-20
C7243 VDD99 a_31571_n16632# 2.21e-19
C7244 F0 Vdiv99 0.229f
C7245 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.514f
C7246 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 5.18e-19
C7247 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 0.00488f
C7248 CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.11f
C7249 RST a_26256_3016# 0.00173f
C7250 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN 9.25e-19
C7251 RST a_54866_n1102# 6.14e-19
C7252 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 4.41e-20
C7253 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_25478_6115# 1.41e-20
C7254 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00118f
C7255 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 a_48832_n1102# 0.00372f
C7256 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 dec3x8_ibr_mag_0.and_3_ibr_5.nand3_mag_ibr_0.OUT 0.0184f
C7257 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_26093_n743# 0.00695f
C7258 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 2.62e-20
C7259 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT a_50150_n15627# 0.0203f
C7260 VDD105 a_44793_5143# 0.00123f
C7261 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 3.38e-19
C7262 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.352f
C7263 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.517f
C7264 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 a_50928_2768# 0.0102f
C7265 RST CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 0.161f
C7266 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT 3.11e-19
C7267 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.121f
C7268 VDD93 a_38966_n8931# 2.27e-19
C7269 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.744f
C7270 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 1.72e-19
C7271 Vdiv105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 8.11e-20
C7272 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 a_36742_n16592# 0.0157f
C7273 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 a_32175_n17626# 5.98e-19
C7274 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 1.85e-19
C7275 VDD99 a_26820_3016# 0.00244f
C7276 Vdiv93 a_43826_n7684# 7.8e-19
C7277 CLK CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 0.165f
C7278 VDD110 Vdiv93 0.26f
C7279 RST a_33744_n17626# 0.00108f
C7280 RST a_34896_n15539# 7.84e-19
C7281 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN m3_20882_n11188# 0.00101f
C7282 a_22460_n9884# a_22620_n9884# 0.0504f
C7283 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 0.0365f
C7284 mux_8x1_ibr_0.mux_2x1_ibr_0.I1 a_38561_880# 0.00372f
C7285 VDD108 a_48258_n10160# 0.0132f
C7286 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 a_23129_n6009# 0.0151f
C7287 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 a_27150_11196# 1.38e-20
C7288 Vdiv99 m3_20882_n11188# 0.295f
C7289 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 1.5f
C7290 CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 0.124f
C7291 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_50269_6240# 0.00119f
C7292 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0377f
C7293 F2 Vdiv 0.0198f
C7294 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 1.26f
C7295 RST CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.00104f
C7296 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.189f
C7297 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_51551_5187# 0.0036f
C7298 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_23794_n17626# 0.00372f
C7299 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 Vdiv110 0.00436f
C7300 CLK CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 3.48e-19
C7301 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 1.1e-19
C7302 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.00586f
C7303 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 1.98e-19
C7304 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_38960_n10028# 1.17e-20
C7305 VDD105 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 0.00791f
C7306 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.359f
C7307 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.109f
C7308 VDD108 Vdiv 0.235f
C7309 CLK CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT 1.46e-19
C7310 Vdiv100 mux_8x1_ibr_0.mux_2x1_ibr_0.I0 0.062f
C7311 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.261f
C7312 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN a_29862_n9832# 5.06e-20
C7313 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.209f
C7314 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.113f
C7315 RST a_47534_n10160# 0.00187f
C7316 F0 a_36310_n1822# 0.0151f
C7317 CLK_div_108_new_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN a_44799_n7920# 0.069f
C7318 VDD99 a_30317_n18723# 3.56e-19
C7319 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_38960_n10028# 0.0202f
C7320 VDD99 a_34308_n17626# 9.82e-19
C7321 RST a_53458_n17599# 0.00247f
C7322 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.652f
C7323 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0502f
C7324 VDD99 a_35460_n15495# 3.14e-19
C7325 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 0.00216f
C7326 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_25702_11196# 0.0036f
C7327 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.0795f
C7328 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.IN2 9.24e-19
C7329 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN 0.516f
C7330 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 0.0127f
C7331 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_29834_n699# 0.00964f
C7332 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.321f
C7333 VDD108 a_46768_n5176# 0.00305f
C7334 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 0.026f
C7335 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 0.101f
C7336 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.00252f
C7337 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 5.6e-19
C7338 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.0725f
C7339 Vdiv110 a_55357_n20487# 0.198f
C7340 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0894f
C7341 VDD93 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.IN2 2.57e-19
C7342 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.359f
C7343 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_28099_n17626# 0.00695f
C7344 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 4.78e-20
C7345 Vdiv96 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 2.42e-19
C7346 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.0477f
C7347 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 0.0204f
C7348 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_25076_n18723# 1.43e-19
C7349 VDD93 a_36667_n10028# 0.0012f
C7350 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0134f
C7351 a_45039_n5176# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.00964f
C7352 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_23706_n2886# 0.00378f
C7353 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT 0.352f
C7354 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT 0.0334f
C7355 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB 0.0378f
C7356 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 0.121f
C7357 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_24391_n20290# 0.00168f
C7358 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 0.00101f
C7359 a_53464_n18696# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0732f
C7360 RST a_32795_11196# 8.64e-19
C7361 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_43760_1671# 0.0114f
C7362 Vdiv108 a_47858_n2243# 6.67e-19
C7363 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 1.18f
C7364 F0 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.IN2 0.162f
C7365 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 0.0635f
C7366 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.14f
C7367 RST CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.103f
C7368 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 a_47492_n5176# 0.0101f
C7369 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_46608_n5176# 0.0202f
C7370 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.103f
C7371 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 0.00182f
C7372 a_24938_n9875# m3_20882_n11188# 6.85e-19
C7373 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_47190_n16726# 0.00789f
C7374 F0 a_36310_880# 0.0151f
C7375 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN a_42521_n13474# 2.7e-20
C7376 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_50669_n6865# 0.0203f
C7377 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 2.82f
C7378 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.0445f
C7379 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_47914_n16726# 0.00696f
C7380 VDD96 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 2.39e-20
C7381 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_43993_n13477# 0.0115f
C7382 F2 a_36042_6821# 5.87e-20
C7383 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN 1.75e-19
C7384 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_30336_10099# 0.0732f
C7385 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN a_30209_7256# 0.069f
C7386 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 1.12e-19
C7387 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 a_51961_6284# 0.00372f
C7388 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 0.23f
C7389 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 a_53934_n9020# 0.0697f
C7390 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB a_48741_9057# 1.86e-20
C7391 Vdiv110 CLK_div_108_new_mag_0.JK_FF_mag_0.QB 0.00103f
C7392 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 1.48e-20
C7393 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_39844_n10028# 8.64e-19
C7394 RST CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.2f
C7395 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB a_50204_2768# 0.00964f
C7396 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 4.25e-20
C7397 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK a_37801_n8887# 9.45e-19
C7398 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 a_22718_8532# 0.0134f
C7399 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 2.96e-19
C7400 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_53249_n6862# 0.0731f
C7401 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00183f
C7402 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 1.22f
C7403 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 3.28e-19
C7404 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 0.434f
C7405 RST CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN 0.00861f
C7406 CLK a_26196_5018# 5.65e-19
C7407 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 2.86e-19
C7408 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 4.8e-20
C7409 VDD96 a_25686_1919# 3.14e-19
C7410 VDD110 a_50441_n17599# 0.00891f
C7411 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT 1.01e-19
C7412 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00354f
C7413 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 a_30760_n20290# 0.0134f
C7414 CLK_div_96_mag_0.JK_FF_mag_4.Q a_23709_810# 0.00239f
C7415 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 9.14e-19
C7416 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_47252_6240# 0.00119f
C7417 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_26990_11196# 1.5e-20
C7418 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.00544f
C7419 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.189f
C7420 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 a_26072_n8734# 6.03e-21
C7421 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB a_22466_n8743# 3.33e-19
C7422 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_28335_6115# 0.00111f
C7423 CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 7.51e-20
C7424 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 a_51285_n1102# 0.069f
C7425 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT a_30210_n13332# 0.0731f
C7426 a_47751_2768# a_47911_2768# 0.0504f
C7427 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 0.026f
C7428 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 0.00494f
C7429 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.28f
C7430 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.401f
C7431 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 a_50922_1671# 0.0697f
C7432 a_36667_n10028# m3_20882_n11188# 3.55e-19
C7433 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 1.54e-19
C7434 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB 0.28f
C7435 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 0.798f
C7436 VDD96 a_22988_n1789# 3.19e-19
C7437 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.12f
C7438 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.08f
C7439 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_44413_n18696# 0.00119f
C7440 a_28574_n9876# a_28734_n9876# 0.0504f
C7441 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_34890_n16636# 1.46e-19
C7442 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 6.82e-19
C7443 RST a_26072_n8734# 0.00126f
C7444 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB 2.46e-21
C7445 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_45363_6284# 4.52e-20
C7446 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_47988_n17599# 0.0102f
C7447 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 a_48023_n7840# 6.83e-19
C7448 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 0.652f
C7449 RST CLK_div_108_new_mag_0.JK_FF_mag_1.CLK 0.0108f
C7450 VDD90 a_23019_5018# 0.00123f
C7451 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 2.34f
C7452 CLK_div_96_mag_0.JK_FF_mag_5.Q a_23709_810# 0.00789f
C7453 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.0795f
C7454 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT a_53940_n10161# 9.1e-19
C7455 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0871f
C7456 RST a_47751_2768# 0.00186f
C7457 CLK CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB 0.363f
C7458 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 a_51604_10154# 1.46e-19
C7459 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.IN1 a_22985_810# 8.64e-19
C7460 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 dec3x8_ibr_mag_0.and_3_ibr_3.nand3_mag_ibr_0.OUT 0.338f
C7461 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB a_51598_9057# 1.41e-20
C7462 RST a_28574_n9876# 0.0017f
C7463 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 0.515f
C7464 CLK_div_96_mag_0.JK_FF_mag_0.QB a_22982_n2930# 0.00695f
C7465 VDD100 a_47905_1671# 3.14e-19
C7466 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB a_22565_n6009# 0.00695f
C7467 CLK_div_108_new_mag_0.JK_FF_mag_1.Q a_51205_n7921# 2.99e-19
C7468 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00154f
C7469 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 1.76e-20
C7470 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0122f
C7471 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 5.05f
C7472 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_44687_n1102# 0.0202f
C7473 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 m3_20882_n11188# 0.00177f
C7474 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 0.25f
C7475 a_44324_1671# CLK_div_100_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 5.94e-20
C7476 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 a_42521_n13474# 0.0202f
C7477 CLK_div_108_new_mag_0.CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN a_50232_n7685# 3.25e-19
C7478 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.118f
C7479 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.45e-19
C7480 RST CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.104f
C7481 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_27529_n18723# 0.069f
C7482 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.121f
C7483 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_105_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00154f
C7484 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 9.73e-19
C7485 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.VOUT CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 5.03e-20
C7486 RST a_29905_n16590# 0.00136f
C7487 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN 0.207f
C7488 VDD99 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 1.08e-20
C7489 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_25420_n13385# 8.64e-19
C7490 VDD108 a_52806_n9020# 3.57e-19
C7491 VDD100 a_47911_2768# 0.00123f
C7492 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00434f
C7493 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 1.08f
C7494 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.122f
C7495 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_28552_354# 1.41e-20
C7496 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_26052_n15491# 3.33e-19
C7497 CLK CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.00324f
C7498 a_27227_398# CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 4.52e-20
C7499 VDD105 a_51034_9057# 3.14e-19
C7500 VDD96 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.28f
C7501 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 a_48944_6284# 0.00372f
C7502 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_33359_11196# 0.0731f
C7503 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 a_50917_n9020# 0.0697f
C7504 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 0.0529f
C7505 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 2.52f
C7506 Vdiv108 a_54537_n6818# 0.00859f
C7507 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_40254_n8887# 4.52e-20
C7508 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 1.02f
C7509 a_54503_1671# a_54663_1671# 0.0504f
C7510 a_23967_10099# a_24127_10099# 0.0504f
C7511 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT 1.74e-19
C7512 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 2.12e-19
C7513 CLK_div_100_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 6.89e-19
C7514 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0894f
C7515 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K a_48092_n9063# 6.09e-21
C7516 RST a_51481_n9064# 0.00154f
C7517 VDD99 RST 7.25f
C7518 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.CLK 1.61f
C7519 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 0.493f
C7520 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_45006_10154# 0.00695f
C7521 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.321f
C7522 VDD100 RST 2.83f
C7523 VDD99 a_30469_n16590# 3.14e-19
C7524 CLK CLK_div_110_mag_0.CLK_div_10_mag_0.CLK 0.0624f
C7525 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.108f
C7526 RST CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.0901f
C7527 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K a_25322_n16632# 8.64e-19
C7528 VDD96 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 0.246f
C7529 RST a_26096_3016# 0.00189f
C7530 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_45724_9057# 0.00111f
C7531 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.195f
C7532 dec3x8_ibr_mag_0.and_3_ibr_0.nand3_mag_ibr_0.OUT dec3x8_ibr_mag_0.and_3_ibr_4.nand3_mag_ibr_0.OUT 0.00141f
C7533 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 a_25650_n1899# 2.37e-20
C7534 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00118f
C7535 RST a_54302_n1102# 6.14e-19
C7536 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.768f
C7537 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.00118f
C7538 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 a_48268_n1102# 0.069f
C7539 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_25318_6115# 1.86e-20
C7540 CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 a_39126_n8931# 2.79e-20
C7541 a_53458_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.46e-19
C7542 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 3.43e-19
C7543 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 a_37328_6265# 0.00103f
C7544 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0016f
C7545 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.0172f
C7546 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 0.768f
C7547 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT 0.0894f
C7548 VDD105 a_44229_5143# 0.00892f
C7549 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT a_47835_7960# 3.38e-20
C7550 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 a_50768_2768# 0.0101f
C7551 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 4.46e-20
C7552 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.233f
C7553 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 0.00975f
C7554 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_37237_n8887# 4.52e-20
C7555 a_51481_n9064# a_51641_n9064# 0.0504f
C7556 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.0894f
C7557 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_52923_9057# 4.52e-20
C7558 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB 0.00585f
C7559 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_25508_n8734# 0.00378f
C7560 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_45131_n17599# 2.88e-20
C7561 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.00975f
C7562 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 m3_20882_n11188# 0.0325f
C7563 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 1.84e-20
C7564 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 0.126f
C7565 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 1.82e-19
C7566 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 a_47816_6284# 6.43e-21
C7567 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 0.0165f
C7568 VDD96 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.994f
C7569 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 a_36178_n16592# 0.00859f
C7570 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 a_32015_n17626# 5.98e-19
C7571 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.00761f
C7572 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 9.88e-20
C7573 VDD99 a_26256_3016# 0.0012f
C7574 Vdiv105 Vdiv110 0.316f
C7575 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.00143f
C7576 CLK dec3x8_ibr_mag_0.and_3_ibr_6.nand3_mag_ibr_0.OUT 0.00229f
C7577 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB 2.59e-21
C7578 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 3.18e-19
C7579 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 1.38e-19
C7580 RST a_33180_n17626# 0.00214f
C7581 CLK_div_108_new_mag_0.JK_FF_mag_1.Q CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.IN2 0.00549f
C7582 VDD100 a_54866_n1102# 3.56e-19
C7583 RST a_34736_n15539# 9.41e-19
C7584 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_42521_n13474# 0.0186f
C7585 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 m3_20882_n11188# 0.00673f
C7586 mux_8x1_ibr_0.mux_2x1_ibr_0.I1 a_37999_880# 0.069f
C7587 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN 1.4e-21
C7588 a_26096_3016# a_26256_3016# 0.0504f
C7589 VDD108 a_48098_n10160# 0.00888f
C7590 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 a_22565_n6009# 0.0102f
C7591 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 2.37f
C7592 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.233f
C7593 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C7594 Vdiv96 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 0.00544f
C7595 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 a_26990_11196# 1.09e-20
C7596 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 a_28583_n1899# 1.01e-20
C7597 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 6.68e-19
C7598 VDD105 Vdiv 0.251f
C7599 VDD mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT 0.659f
C7600 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 2.34e-19
C7601 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.0838f
C7602 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00157f
C7603 RST a_43757_n6273# 5.78e-20
C7604 VDD93 a_24778_n9875# 0.00108f
C7605 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00279f
C7606 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00118f
C7607 CLK_div_108_new_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 0.00384f
C7608 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_44055_n16724# 8.66e-20
C7609 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C7610 a_51652_2768# Vdiv110 0.00138f
C7611 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 F0 7.46e-21
C7612 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 0.00103f
C7613 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 9.73e-19
C7614 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK a_47190_n16726# 0.00193f
C7615 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN a_29298_n9832# 1.76e-20
C7616 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK 4.24f
C7617 RST a_47374_n10160# 0.00228f
C7618 F0 a_35747_n1822# 9.5e-19
C7619 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 0.0591f
C7620 VDD99 a_33744_n17626# 0.00149f
C7621 RST a_53298_n17599# 0.00247f
C7622 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 3.84e-20
C7623 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 6.89e-19
C7624 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.103f
C7625 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT a_32455_n16632# 2.88e-20
C7626 F1 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 0.16f
C7627 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT 0.117f
C7628 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 a_52115_5187# 0.00372f
C7629 CLK a_50281_n17599# 3.76e-20
C7630 CLK_div_105_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.00154f
C7631 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 0.0153f
C7632 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 2.81e-20
C7633 CLK CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 5.14e-20
C7634 RST CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.0545f
C7635 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.122f
C7636 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_29270_n743# 0.00696f
C7637 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.654f
C7638 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_45695_n17599# 0.0036f
C7639 VDD108 a_46608_n5176# 0.00743f
C7640 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB a_48092_n9063# 0.00392f
C7641 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.00584f
C7642 Vdiv110 a_55197_n20487# 0.0132f
C7643 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_53464_n18696# 0.00119f
C7644 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_27939_n17626# 0.00696f
C7645 VDD96 a_23139_n287# 3.18e-19
C7646 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C7647 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 0.0814f
C7648 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_24512_n18723# 0.011f
C7649 VDD93 a_36103_n10028# 0.00888f
C7650 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_23142_n2930# 0.0733f
C7651 VDD110 dec3x8_ibr_mag_0.and_3_ibr_6.nand3_mag_ibr_0.OUT 0.00134f
C7652 CLK_div_108_new_mag_0.JK_FF_mag_0.QB CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.343f
C7653 a_53304_n18696# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0203f
C7654 RST a_32635_11196# 0.00151f
C7655 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.00216f
C7656 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0378f
C7657 Vdiv108 a_47698_n2243# 6.67e-19
C7658 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.00488f
C7659 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.106f
C7660 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 a_47332_n5176# 0.0102f
C7661 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 a_47030_n16726# 0.00335f
C7662 a_24778_n9875# m3_20882_n11188# 6.85e-19
C7663 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 a_30502_11196# 0.00335f
C7664 F0 a_35747_880# 9.5e-19
C7665 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.111f
C7666 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.00154f
C7667 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.122f
C7668 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_50105_n6865# 1.5e-20
C7669 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.352f
C7670 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 3.67e-20
C7671 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.792f
C7672 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 a_40375_n7552# 8.64e-19
C7673 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_47754_n16726# 0.00695f
C7674 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 8.16e-20
C7675 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.0835f
C7676 a_34736_n15539# a_34896_n15539# 0.0504f
C7677 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.122f
C7678 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_29772_10099# 0.00378f
C7679 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00542f
C7680 CLK CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.00289f
C7681 dec3x8_ibr_mag_0.and_3_ibr_5.IN3 dec3x8_ibr_mag_0.and_3_ibr_0.nand3_mag_ibr_0.OUT 0.245f
C7682 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 0.779f
C7683 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 a_51397_6284# 0.069f
C7684 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 a_48986_n2199# 0.00372f
C7685 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 a_53370_n9020# 0.0059f
C7686 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT 0.257f
C7687 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB a_48581_9057# 1.41e-20
C7688 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.125f
C7689 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.0979f
C7690 a_30881_n18723# CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 4.9e-20
C7691 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB a_49640_2768# 0.0811f
C7692 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK a_37237_n8887# 6.06e-21
C7693 VDD100 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.00115f
C7694 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.00118f
C7695 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.765f
C7696 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_53089_n6862# 0.0202f
C7697 CLK a_26036_5018# 5.65e-19
C7698 a_43757_n6273# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0732f
C7699 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 0.286f
C7700 VDD96 a_25122_1919# 3.56e-19
C7701 RST CLK_div_100_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 0.00649f
C7702 VDD110 a_50281_n17599# 0.0132f
C7703 CLK_div_90_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_90_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.11f
C7704 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 2.89e-19
C7705 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 2f
C7706 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN 0.00165f
C7707 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 5.06e-21
C7708 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00137f
C7709 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_26426_11196# 0.0203f
C7710 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 1.4e-20
C7711 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.995f
C7712 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB a_21902_n8787# 0.00392f
C7713 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_48534_5187# 0.0036f
C7714 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00122f
C7715 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 5.08f
C7716 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_27170_6159# 7.4e-19
C7717 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 0.00335f
C7718 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT a_30050_n13332# 0.0202f
C7719 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 a_37999_280# 0.00375f
C7720 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 a_50358_1671# 0.0059f
C7721 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_54947_n5721# 0.00372f
C7722 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 0.0709f
C7723 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 a_29862_n9832# 0.0157f
C7724 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 0.0172f
C7725 a_36103_n10028# m3_20882_n11188# 8.45e-19
C7726 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 1.55e-19
C7727 VDD96 a_26980_3016# 0.00108f
C7728 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 0.109f
C7729 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 1.94e-20
C7730 CLK_div_105_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 3.87e-19
C7731 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 6.89e-19
C7732 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.VOUT CLK_div_93_mag_0.CLK_div_3_mag_0.CLK 0.198f
C7733 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00233f
C7734 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.0592f
C7735 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB 0.25f
C7736 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 a_28010_n9876# 0.00214f
C7737 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 1.89e-21
C7738 a_47374_n10160# a_47534_n10160# 0.0504f
C7739 RST a_25508_n8734# 6.86e-19
C7740 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_44799_6284# 0.0202f
C7741 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 9.62e-20
C7742 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_47424_n17599# 0.00789f
C7743 dec3x8_ibr_mag_0.and_3_ibr_1.nand3_mag_ibr_0.OUT dec3x8_ibr_mag_0.and_3_ibr_2.nand3_mag_ibr_0.OUT 7.01e-19
C7744 VDD90 a_22455_5018# 0.00892f
C7745 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.36f
C7746 a_53298_n17599# a_53458_n17599# 0.0504f
C7747 CLK_div_96_mag_0.JK_FF_mag_5.Q a_23145_810# 0.0102f
C7748 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.122f
C7749 RST a_47187_2768# 9.41e-19
C7750 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT a_53780_n10161# 2.88e-20
C7751 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.313f
C7752 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN a_55019_7683# 2.85e-20
C7753 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 8.24e-19
C7754 Vdiv105 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT 1.33e-19
C7755 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.391f
C7756 CLK_div_108_new_mag_0.JK_FF_mag_1.Q CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 9.71e-20
C7757 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 7.17e-19
C7758 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 a_36202_6821# 8.64e-19
C7759 VDD108 RST 6.77f
C7760 RST a_28010_n9876# 0.00189f
C7761 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.JK_FF_mag_5.Q 0.161f
C7762 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0894f
C7763 Vdiv105 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT 3e-19
C7764 Vdiv90 Vdiv96 1.37f
C7765 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.432f
C7766 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.0343f
C7767 F1 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 0.16f
C7768 RST CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 9.24e-20
C7769 dec3x8_ibr_mag_0.and_3_ibr_5.IN3 a_37168_6821# 0.00657f
C7770 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 9.62e-20
C7771 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB a_22405_n6009# 0.00696f
C7772 VDD100 a_47341_1671# 3.14e-19
C7773 CLK_div_108_new_mag_0.JK_FF_mag_1.Q a_50232_n7685# 0.00263f
C7774 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00545f
C7775 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 0.338f
C7776 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0345f
C7777 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 a_50833_6284# 1.25e-20
C7778 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 a_29214_n6271# 0.00347f
C7779 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0298f
C7780 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 0.15f
C7781 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 a_53738_n1102# 6.43e-21
C7782 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 1.18f
C7783 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 9.52e-19
C7784 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C7785 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.768f
C7786 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT 0.0854f
C7787 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 a_49906_9057# 4.52e-20
C7788 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_26965_n18723# 0.00372f
C7789 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_44475_n5176# 2.88e-20
C7790 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0715f
C7791 CLK_div_108_new_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 3.67e-20
C7792 RST a_29341_n16634# 0.00222f
C7793 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 a_28617_n16634# 1.46e-19
C7794 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 1.12e-19
C7795 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.108f
C7796 VDD108 a_51641_n9064# 2.21e-19
C7797 VDD100 a_47751_2768# 0.00101f
C7798 RST CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 0.105f
C7799 a_30060_9000# CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 1.87e-19
C7800 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.00196f
C7801 a_26183_n7107# a_26343_n7107# 0.0504f
C7802 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT a_35614_n16636# 2.88e-20
C7803 Vdiv110 mux_8x1_ibr_0.mux_2x1_ibr_0.I1 0.00876f
C7804 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 1.64e-20
C7805 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_25488_n15535# 0.00392f
C7806 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_28392_354# 1.86e-20
C7807 Vdiv90 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 0.0537f
C7808 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.321f
C7809 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00917f
C7810 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 0.209f
C7811 VDD105 a_50470_9057# 3.14e-19
C7812 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 a_48380_6284# 0.069f
C7813 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_32795_11196# 9.1e-19
C7814 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 a_50353_n9020# 0.0059f
C7815 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_39690_n8887# 0.0202f
C7816 Vdiv108 a_53973_n6862# 0.0101f
C7817 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 9.9e-19
C7818 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 0.00335f
C7819 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.391f
C7820 Vdiv96 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 0.00292f
C7821 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.00123f
C7822 RST a_50917_n9020# 5.61e-19
C7823 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 0.28f
C7824 CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 2f
C7825 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00976f
C7826 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.0151f
C7827 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_44846_10154# 0.00696f
C7828 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C7829 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.4f
C7830 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 0.198f
C7831 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_53174_n1146# 1.41e-20
C7832 VDD99 a_29905_n16590# 3.14e-19
C7833 a_32635_11196# a_32795_11196# 0.0504f
C7834 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 1f
C7835 CLK CLK_div_96_mag_0.JK_FF_mag_4.QB 0.307f
C7836 Vdiv110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB 9.33e-19
C7837 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.018f
C7838 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_45564_9057# 0.00486f
C7839 RST a_25532_3016# 0.00101f
C7840 RST a_53738_n1102# 2.78e-19
C7841 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB 3.95e-19
C7842 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_24153_6159# 0.0114f
C7843 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 a_37168_6265# 8.19e-19
C7844 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.431f
C7845 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.0622f
C7846 CLK_div_96_mag_0.JK_FF_mag_2.QB CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.198f
C7847 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 0.00116f
C7848 VDD105 a_44069_5143# 0.0132f
C7849 RST CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.00717f
C7850 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.00602f
C7851 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 a_50204_2768# 0.00859f
C7852 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.161f
C7853 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0838f
C7854 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 6.46e-19
C7855 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.925f
C7856 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_36673_n8887# 0.0202f
C7857 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_24944_n8778# 0.0732f
C7858 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_44971_n17599# 9.1e-19
C7859 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 6.11e-19
C7860 RST CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 0.311f
C7861 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 0.285f
C7862 CLK_div_96_mag_0.JK_FF_mag_2.Q CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 1.48e-20
C7863 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 1.12e-19
C7864 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 a_51871_n5# 0.0084f
C7865 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 a_47252_6240# 0.00939f
C7866 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.65f
C7867 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0143f
C7868 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 a_35614_n16636# 0.0101f
C7869 VDD99 a_26096_3016# 0.0012f
C7870 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT 0.00982f
C7871 RST a_30496_10099# 7.78e-19
C7872 CLK_div_100_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00943f
C7873 VDD100 a_54302_n1102# 3.14e-19
C7874 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 0.122f
C7875 VDD110 a_55156_n18696# 3.56e-19
C7876 RST CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0732f
C7877 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 4.24e-20
C7878 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN a_28268_n6266# 4.6e-21
C7879 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 a_36873_280# 0.00372f
C7880 VDD108 a_47534_n10160# 0.0012f
C7881 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 a_22405_n6009# 0.0101f
C7882 RST a_32230_5018# 0.00127f
C7883 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 CLK_div_96_mag_0.JK_FF_mag_2.Q 4.57e-20
C7884 RST a_43597_n6273# 7.14e-20
C7885 VDD93 a_23748_n9840# 3.14e-19
C7886 F0 a_36873_n1222# 2.62e-19
C7887 VDD93 a_35184_n1822# 3.39e-19
C7888 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 m3_20882_n11188# 0.00217f
C7889 a_51492_2768# Vdiv110 0.00138f
C7890 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 a_30244_398# 0.069f
C7891 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 0.484f
C7892 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT a_22988_n1789# 3.64e-20
C7893 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 0.167f
C7894 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT 0.00118f
C7895 CLK_div_100_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 3.38e-19
C7896 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK a_47030_n16726# 0.00193f
C7897 a_55161_n15587# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 4.52e-20
C7898 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 2.75e-19
C7899 VDD110 a_52385_n13362# 0.0418f
C7900 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 a_55315_n16684# 0.00372f
C7901 F0 a_35184_n1822# 0.0144f
C7902 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 0.00243f
C7903 RST a_46810_n10116# 0.00164f
C7904 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 5.7e-20
C7905 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB a_45724_9057# 1.86e-20
C7906 Vdiv mux_8x1_ibr_0.mux_2x1_ibr_0.I0 1.49e-19
C7907 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.397f
C7908 VDD99 a_33180_n17626# 0.00149f
C7909 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.00125f
C7910 VDD99 a_34736_n15539# 2.21e-19
C7911 CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K 0.00205f
C7912 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT a_32295_n16632# 9.1e-19
C7913 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 6.11e-19
C7914 F1 a_36873_280# 1.8e-19
C7915 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_41284_n14596# 1.75e-19
C7916 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 a_51551_5187# 0.069f
C7917 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT a_45899_7960# 3.92e-20
C7918 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00367f
C7919 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB 0.103f
C7920 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 0.0622f
C7921 RST CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN 0.00968f
C7922 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.783f
C7923 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 a_23948_n18723# 0.069f
C7924 CLK CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.449f
C7925 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.866f
C7926 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_29110_n743# 0.00695f
C7927 CLK_div_96_mag_0.JK_FF_mag_3.Q a_27227_398# 9.45e-19
C7928 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 0.122f
C7929 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB a_47528_n9019# 3.33e-19
C7930 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 2.81e-20
C7931 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_50157_n1146# 1.41e-20
C7932 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_27375_n17626# 0.00964f
C7933 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 0.124f
C7934 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 2.01e-19
C7935 VDD96 a_22575_n287# 3.18e-19
C7936 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_23948_n18723# 0.00118f
C7937 VDD93 a_35943_n10028# 0.0132f
C7938 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.122f
C7939 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.0836f
C7940 VDD93 a_35184_880# 3.39e-19
C7941 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_22982_n2930# 0.0203f
C7942 a_53304_n18696# a_53464_n18696# 0.0504f
C7943 RST a_32071_11196# 8.68e-19
C7944 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.338f
C7945 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 0.768f
C7946 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 0.00118f
C7947 Vdiv108 a_47134_n2243# 0.00158f
C7948 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0635f
C7949 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT 3.09e-19
C7950 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 a_28617_n16634# 4.52e-19
C7951 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 a_46768_n5176# 0.00789f
C7952 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.11f
C7953 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 2.11e-20
C7954 a_25055_n7107# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB 4.61e-20
C7955 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.657f
C7956 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 a_30342_11196# 0.00789f
C7957 a_23748_n9840# m3_20882_n11188# 3e-19
C7958 F0 a_35184_880# 0.0163f
C7959 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_49945_n6865# 1.17e-20
C7960 CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 a_53174_n1146# 2.79e-20
C7961 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN 1.36e-19
C7962 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 7.06e-19
C7963 CLK_div_96_mag_0.JK_FF_mag_5.QB CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 1.4e-19
C7964 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00352f
C7965 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 8.98e-19
C7966 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.00132f
C7967 a_52806_n9020# CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 4.52e-20
C7968 a_24922_n17626# a_25082_n17626# 0.0504f
C7969 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.00187f
C7970 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 0.359f
C7971 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 0.904f
C7972 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0622f
C7973 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 1.94f
C7974 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB 0.103f
C7975 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.121f
C7976 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 0.0435f
C7977 CLK a_52161_n19793# 2.22e-19
C7978 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 a_48422_n2199# 0.069f
C7979 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_2x1_ibr_0.I1 0.329f
C7980 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 7.24e-19
C7981 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 3.14f
C7982 a_28386_n743# a_28546_n743# 0.0504f
C7983 RST CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.00571f
C7984 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN 0.303f
C7985 F1 a_39580_6821# 0.0103f
C7986 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 0.491f
C7987 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK a_36673_n8887# 6.43e-21
C7988 RST CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 3.79e-19
C7989 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 1.41e-20
C7990 a_22985_810# a_23145_810# 0.0504f
C7991 CLK a_25472_5018# 0.00134f
C7992 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.00103f
C7993 a_43597_n6273# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0203f
C7994 CLK_div_96_mag_0.JK_FF_mag_0.QB CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.199f
C7995 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 CLK_div_90_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 8.04e-19
C7996 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 4.39e-19
C7997 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN 0.00956f
C7998 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 8.16e-20
C7999 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.321f
C8000 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 0.321f
C8001 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_55161_n15587# 0.0114f
C8002 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.122f
C8003 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_26266_11196# 0.0733f
C8004 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_55315_n16684# 0.0811f
C8005 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 a_46889_9057# 4.52e-20
C8006 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 4.2e-19
C8007 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 1.93f
C8008 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 a_24944_n8778# 2.79e-20
C8009 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB 2.42e-21
C8010 VDD108 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK 1.42f
C8011 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_26606_6159# 7.4e-19
C8012 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.101f
C8013 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_54383_n5721# 0.069f
C8014 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 0.0209f
C8015 a_35943_n10028# m3_20882_n11188# 8.45e-19
C8016 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 a_29298_n9832# 0.00859f
C8017 RST a_48747_10154# 0.00186f
C8018 F1 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 0.00224f
C8019 VDD96 a_22264_n1833# 0.00534f
C8020 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.0435f
C8021 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.198f
C8022 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 a_30341_5062# 0.00372f
C8023 RST CLK_div_108_new_mag_0.JK_FF_mag_1.QB 0.168f
C8024 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 a_27850_n9876# 0.00182f
C8025 RST a_24944_n8778# 0.00229f
C8026 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.352f
C8027 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.122f
C8028 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_54866_n1102# 0.0114f
C8029 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_47264_n17599# 0.00335f
C8030 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 0.249f
C8031 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_22275_10099# 4.52e-20
C8032 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0894f
C8033 VDD105 RST 2.84f
C8034 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 8.02e-20
C8035 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT 4.36e-19
C8036 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 5.11e-19
C8037 VDD90 a_22295_5018# 0.0132f
C8038 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 0.399f
C8039 CLK_div_96_mag_0.JK_FF_mag_5.Q a_22985_810# 0.0101f
C8040 RST a_46623_2768# 9.66e-19
C8041 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT 0.0121f
C8042 F0 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 0.136f
C8043 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0175f
C8044 RST a_27850_n9876# 0.00189f
C8045 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.74f
C8046 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 0.00335f
C8047 VDD110 a_52161_n19793# 3.14e-19
C8048 CLK_div_105_mag_0.CLK_div_10_mag_1.CLK CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 3.1e-22
C8049 VDD100 a_46777_1671# 3.56e-19
C8050 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB a_21841_n6009# 0.00964f
C8051 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB a_53940_n10161# 0.00695f
C8052 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K 0.0484f
C8053 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 a_50269_6240# 0.00939f
C8054 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 3.38e-19
C8055 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 2.86e-19
C8056 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 5.18e-20
C8057 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 a_53174_n1146# 0.00939f
C8058 VDD99 F2 0.296f
C8059 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 1.82e-19
C8060 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_44315_n5176# 9.1e-19
C8061 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_40408_n9984# 0.0036f
C8062 CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 8.98e-19
C8063 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 0.0285f
C8064 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 8.16e-20
C8065 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.0343f
C8066 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 0.0592f
C8067 VDD100 F2 0.0978f
C8068 RST a_29181_n16634# 0.00206f
C8069 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_53286_6240# 1.41e-20
C8070 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 1f
C8071 VDD90 a_30060_9000# 5.92e-19
C8072 CLK CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.471f
C8073 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 a_51758_9057# 0.0101f
C8074 VDD100 a_47187_2768# 0.00152f
C8075 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0622f
C8076 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT a_35454_n16636# 9.1e-19
C8077 CLK CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 1.48e-20
C8078 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.523f
C8079 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.349f
C8080 VDD100 VDD108 0.748f
C8081 VDD105 a_49906_9057# 3.56e-19
C8082 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_32635_11196# 2.88e-20
C8083 a_53897_10154# a_54057_10154# 0.0504f
C8084 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0205f
C8085 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 1.16f
C8086 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.0622f
C8087 Vdiv108 a_53813_n6862# 0.0102f
C8088 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK 5.6e-20
C8089 CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 1.99e-19
C8090 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C8091 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT a_23139_n287# 0.0202f
C8092 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.231f
C8093 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.00975f
C8094 RST a_50353_n9020# 5.02e-19
C8095 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 0.0398f
C8096 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00531f
C8097 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_44282_10154# 0.00964f
C8098 VDD90 a_24127_10099# 2.21e-19
C8099 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_0.OUT 0.0888f
C8100 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_4.IN2 a_22011_n287# 4.52e-20
C8101 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 3.71e-20
C8102 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_53014_n1146# 1.86e-20
C8103 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 Vdiv108 0.0335f
C8104 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 2.47e-19
C8105 a_23973_11196# a_24133_11196# 0.0504f
C8106 VDD99 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 1.08e-20
C8107 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_45000_9057# 3.25e-19
C8108 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.394f
C8109 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C8110 RST a_24968_3016# 0.00101f
C8111 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 3.43e-19
C8112 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_23589_6159# 2.96e-19
C8113 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 0.39f
C8114 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 0.215f
C8115 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN 0.00617f
C8116 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN 0.107f
C8117 RST CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.055f
C8118 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT a_51764_10154# 1.17e-20
C8119 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0622f
C8120 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 0.0655f
C8121 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.431f
C8122 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 0.0205f
C8123 RST CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_4.IN2 0.00125f
C8124 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 4.75e-20
C8125 a_52293_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.0811f
C8126 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 a_49640_2768# 0.0157f
C8127 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_2.OUT CLK_div_96_mag_0.JK_FF_mag_5.QB 0.103f
C8128 CLK CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.0215f
C8129 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_24784_n8778# 0.0203f
C8130 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_44407_n17599# 0.0731f
C8131 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.00205f
C8132 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 8.97e-19
C8133 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 7.49e-20
C8134 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 1f
C8135 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 a_47092_6240# 0.0101f
C8136 VDD108 a_43757_n6273# 2.65e-19
C8137 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_45251_n1102# 0.0059f
C8138 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 8.59e-20
C8139 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 a_35454_n16636# 0.0102f
C8140 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB 6.46e-19
C8141 VDD99 a_25532_3016# 0.00146f
C8142 RST a_30336_10099# 6.43e-19
C8143 CLK_div_105_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 a_43831_7266# 9.02e-19
C8144 VDD100 a_53738_n1102# 3.14e-19
C8145 VDD110 a_54592_n18696# 3.14e-19
C8146 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 6.82e-19
C8147 VDD108 a_47374_n10160# 9.82e-19
C8148 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.29f
C8149 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 a_21841_n6009# 0.00859f
C8150 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 3.38e-19
C8151 RST CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.0798f
C8152 CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 3.27e-19
C8153 RST a_32070_5018# 0.00169f
C8154 mux_8x1_ibr_0.mux_2x1_ibr_0.I0 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.OUT 0.419f
C8155 a_50903_n5# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 3.38e-20
C8156 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 8.04e-19
C8157 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 a_53732_n2243# 3.6e-22
C8158 RST a_31129_n6271# 6.53e-20
C8159 VDD93 a_23184_n9840# 3.14e-19
C8160 F0 a_35747_n1222# 6.89e-19
C8161 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00136f
C8162 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_50263_5143# 1.46e-19
C8163 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT F2 4.43e-19
C8164 CLK CLK_div_99_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.00338f
C8165 a_50928_2768# Vdiv110 5.84e-19
C8166 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00166f
C8167 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.27f
C8168 CLK CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00118f
C8169 a_53008_n2243# a_53168_n2243# 0.0504f
C8170 VDD110 a_52225_n13362# 0.235f
C8171 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_2.OUT 3.81e-20
C8172 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 a_54751_n16684# 0.069f
C8173 a_48148_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0733f
C8174 RST a_46246_n10116# 0.00114f
C8175 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_50269_6240# 1.41e-20
C8176 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.742f
C8177 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_2.OUT CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 0.00118f
C8178 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 0.0635f
C8179 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT 0.768f
C8180 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB a_45564_9057# 1.41e-20
C8181 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT 0.00296f
C8182 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.652f
C8183 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.0343f
C8184 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT a_31731_n16632# 0.0731f
C8185 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.00205f
C8186 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K F1 3.36e-20
C8187 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 0.191f
C8188 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_41124_n14596# 0.00369f
C8189 CLK_div_100_mag_0.CLK_div_10_mag_1.CLK CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.122f
C8190 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.233f
C8191 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 a_46755_574# 1.29e-22
C8192 a_39420_6821# a_39580_6821# 0.0504f
C8193 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 9.45e-20
C8194 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.122f
C8195 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 1.22e-19
C8196 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_24133_11196# 0.0202f
C8197 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 4.64e-20
C8198 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 a_43826_n7684# 8.64e-19
C8199 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 8.19e-19
C8200 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.122f
C8201 RST CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 0.0625f
C8202 CLK_div_96_mag_0.JK_FF_mag_3.Q a_26663_398# 6.06e-21
C8203 CLK Vdiv110 1.88f
C8204 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.121f
C8205 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.346f
C8206 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_32225_10099# 0.069f
C8207 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_49997_n1146# 1.86e-20
C8208 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 5.76e-20
C8209 CLK a_44687_n1102# 6.43e-21
C8210 CLK_div_108_new_mag_0.JK_FF_mag_0.QB CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.0378f
C8211 VDD96 a_22011_n287# 3.6e-19
C8212 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_26811_n17626# 0.0811f
C8213 CLK_div_105_mag_0.CLK_div_10_mag_1.CLK CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.122f
C8214 RST CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 0.213f
C8215 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.16f
C8216 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 a_51764_10154# 0.00335f
C8217 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00229f
C8218 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_22418_n2930# 1.5e-20
C8219 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00118f
C8220 RST a_31507_11196# 0.00192f
C8221 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.088f
C8222 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_50675_n5724# 0.00378f
C8223 Vdiv108 a_46974_n2243# 0.00158f
C8224 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K a_53304_n18696# 8.64e-19
C8225 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 a_28457_n16634# 5.83e-19
C8226 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 5.11e-19
C8227 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 a_46608_n5176# 0.00335f
C8228 a_23184_n9840# m3_20882_n11188# 2.88e-19
C8229 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 a_29778_11196# 0.0102f
C8230 a_52923_9057# CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 2.05e-19
C8231 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN 0.111f
C8232 RST CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.313f
C8233 VDD96 RST 3.16f
C8234 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.654f
C8235 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 a_45603_n5176# 0.0157f
C8236 CLK a_30760_n20290# 0.00132f
C8237 VDD mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT 0.663f
C8238 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.28f
C8239 Vdiv90 Vdiv93 7.8e-19
C8240 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.0495f
C8241 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 Vdiv108 1.36e-19
C8242 F1 a_39420_6821# 0.00741f
C8243 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK a_36109_n8931# 0.00939f
C8244 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 4.31e-19
C8245 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 0.122f
C8246 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.109f
C8247 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK CLK_div_108_new_mag_0.JK_FF_mag_1.QB 0.307f
C8248 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB 0.144f
C8249 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN 0.514f
C8250 CLK a_25312_5018# 0.00134f
C8251 a_43597_n6273# a_43757_n6273# 0.0504f
C8252 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_54978_6284# 0.0114f
C8253 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_22718_8532# 0.00168f
C8254 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_54597_n15587# 2.96e-19
C8255 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 8.58e-20
C8256 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.653f
C8257 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 0.313f
C8258 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.792f
C8259 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_25702_11196# 0.00378f
C8260 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_54751_n16684# 0.00964f
C8261 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.27f
C8262 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 0.0854f
C8263 VDD110 Vdiv110 0.544f
C8264 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_26042_6159# 3.12e-19
C8265 a_51983_7381# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 1.29e-22
C8266 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 0.231f
C8267 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB 0.915f
C8268 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 a_47453_9057# 0.069f
C8269 VDD99 dec3x8_ibr_mag_0.and_3_ibr_5.nand3_mag_ibr_0.OUT 0.158f
C8270 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB 1.14e-19
C8271 RST a_48587_10154# 0.00186f
C8272 VDD96 a_26256_3016# 2.21e-19
C8273 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 a_28734_n9876# 0.0101f
C8274 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 0.29f
C8275 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 m3_20882_n11188# 0.0326f
C8276 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_46259_n17599# 0.00372f
C8277 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 1.65f
C8278 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 8.16e-20
C8279 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.398f
C8280 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.507f
C8281 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 3.72e-19
C8282 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 1.85e-19
C8283 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 a_29777_5062# 0.069f
C8284 RST a_24784_n8778# 0.003f
C8285 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_54302_n1102# 2.96e-19
C8286 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.122f
C8287 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN m3_20882_n11188# 2.88e-19
C8288 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_25076_n18723# 0.0202f
C8289 a_30209_7256# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 1.45e-20
C8290 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.00488f
C8291 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.338f
C8292 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT a_35460_n15495# 0.00378f
C8293 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB 0.103f
C8294 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB 0.0835f
C8295 CLK_div_96_mag_0.JK_FF_mag_5.Q a_22421_810# 0.00859f
C8296 RST CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 1.1f
C8297 Vdiv100 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT 1.7e-19
C8298 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_22685_11196# 0.069f
C8299 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 a_50316_10154# 0.0036f
C8300 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 0.00528f
C8301 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.398f
C8302 CLK_div_96_mag_0.JK_FF_mag_3.QB CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.0592f
C8303 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.0275f
C8304 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 0.0275f
C8305 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 2.39e-21
C8306 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.0979f
C8307 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.125f
C8308 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT 0.269f
C8309 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.0228f
C8310 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB a_21277_n6009# 0.0811f
C8311 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_29777_5062# 0.00378f
C8312 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB a_53780_n10161# 0.00696f
C8313 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.994f
C8314 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.00975f
C8315 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN m3_20882_n11188# 0.00101f
C8316 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 a_50109_6240# 0.0101f
C8317 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.0529f
C8318 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00952f
C8319 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT a_53934_n9020# 0.0202f
C8320 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 3.38e-19
C8321 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 a_53014_n1146# 0.0101f
C8322 VDD105 VDD99 0.0582f
C8323 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.103f
C8324 RST CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 0.0958f
C8325 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 0.016f
C8326 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT 0.0173f
C8327 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_43751_n5176# 0.0731f
C8328 VDD105 VDD100 1.1f
C8329 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_53126_6240# 1.86e-20
C8330 RST a_28617_n16634# 0.00273f
C8331 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 0.4f
C8332 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT 0.0238f
C8333 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB m3_20882_n11188# 0.00326f
C8334 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 3.37e-21
C8335 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 a_51598_9057# 0.00939f
C8336 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.00164f
C8337 VDD100 a_46623_2768# 0.00152f
C8338 VDD108 a_50917_n9020# 3.14e-19
C8339 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT a_34890_n16636# 0.0731f
C8340 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 0.00125f
C8341 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0024f
C8342 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.395f
C8343 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.0495f
C8344 Vdiv108 a_53249_n6862# 0.00789f
C8345 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 2.77e-19
C8346 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.VOUT CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 4e-20
C8347 CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 3.39e-20
C8348 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K 0.487f
C8349 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 0.0592f
C8350 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.0718f
C8351 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0352f
C8352 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 3.92e-19
C8353 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0346f
C8354 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT a_22575_n287# 4.52e-20
C8355 RST a_49789_n9020# 5.02e-19
C8356 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB 0.25f
C8357 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_43718_10154# 0.0811f
C8358 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.318f
C8359 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.392f
C8360 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_51849_n1102# 0.0114f
C8361 VDD99 a_29181_n16634# 2.21e-19
C8362 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_45363_6284# 0.0059f
C8363 CLK_div_100_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_55067_297# 5.39e-20
C8364 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_44436_9057# 2.96e-19
C8365 VDD90 a_24133_11196# 0.00743f
C8366 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 0.226f
C8367 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 0.497f
C8368 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.391f
C8369 CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C8370 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 0.995f
C8371 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 8.58e-20
C8372 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_23025_6159# 3.33e-19
C8373 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 1.49e-19
C8374 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.211f
C8375 RST CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.00219f
C8376 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT a_51604_10154# 1.5e-20
C8377 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 9.66e-19
C8378 VDD93 a_28267_n7033# 3.14e-19
C8379 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT 0.345f
C8380 a_51729_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.00964f
C8381 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.74f
C8382 Vdiv108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 1.8e-21
C8383 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 9.05e-22
C8384 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB 1.99f
C8385 RST CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.335f
C8386 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00131f
C8387 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.178f
C8388 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.0948f
C8389 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_44247_n17599# 0.0202f
C8390 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 a_25806_n17626# 0.00335f
C8391 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.649f
C8392 CLK_div_96_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 6.11e-19
C8393 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_48466_n6273# 0.00372f
C8394 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 a_45927_6284# 0.069f
C8395 VDD108 a_43597_n6273# 5.99e-19
C8396 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_44687_n1102# 0.0697f
C8397 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 a_30165_n6282# 9.22e-21
C8398 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0385f
C8399 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 a_34890_n16636# 0.00789f
C8400 CLK CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 1.2e-19
C8401 VDD99 a_24968_3016# 0.00149f
C8402 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 a_51983_7381# 0.0084f
C8403 RST a_29772_10099# 3.71e-19
C8404 CLK CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 1.31f
C8405 CLK_div_105_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 a_43671_7266# 2.44e-20
C8406 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1.21e-19
C8407 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.741f
C8408 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00118f
C8409 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.394f
C8410 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 0.409f
C8411 CLK_div_108_new_mag_0.JK_FF_mag_1.Q CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 0.00335f
C8412 VDD110 a_54028_n18696# 3.14e-19
C8413 a_21736_n9884# a_21896_n9884# 0.0504f
C8414 a_28583_n1899# a_28743_n1899# 0.0504f
C8415 VDD108 a_46810_n10116# 0.00149f
C8416 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 a_43559_n120# 0.019f
C8417 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 a_21277_n6009# 0.0157f
C8418 RST a_31506_5018# 0.00186f
C8419 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.395f
C8420 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 a_53168_n2243# 1.86e-20
C8421 RST CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN 0.0163f
C8422 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 4.11e-19
C8423 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 1.65e-21
C8424 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0995f
C8425 VDD110 a_55161_n15587# 3.56e-19
C8426 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.122f
C8427 a_50768_2768# Vdiv110 5.84e-19
C8428 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 0.128f
C8429 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K m3_20882_n11188# 0.00466f
C8430 VDD110 a_55315_n16684# 3.14e-19
C8431 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.647f
C8432 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT a_50917_n9020# 0.0202f
C8433 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_40972_n9984# 0.00372f
C8434 Vdiv90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 3.1e-22
C8435 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_40254_n8887# 0.0059f
C8436 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 0.294f
C8437 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 1.83e-19
C8438 VDD110 a_49488_n13383# 3.14e-19
C8439 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 5.11e-19
C8440 a_47988_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0203f
C8441 RST a_45241_n10160# 0.00218f
C8442 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_50109_6240# 1.86e-20
C8443 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.27f
C8444 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 a_30187_6159# 9.45e-19
C8445 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 0.026f
C8446 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT a_31571_n16632# 0.0202f
C8447 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 9.73e-19
C8448 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 0.0011f
C8449 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.311f
C8450 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 2.64e-19
C8451 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 0.994f
C8452 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_23973_11196# 0.0731f
C8453 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB 0.0384f
C8454 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.121f
C8455 RST CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.265f
C8456 VDD mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 0.402f
C8457 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 0.00394f
C8458 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_36742_n16592# 0.0811f
C8459 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 0.492f
C8460 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00118f
C8461 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.00158f
C8462 CLK_div_96_mag_0.JK_FF_mag_3.Q a_26099_398# 6.43e-21
C8463 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB a_46400_n9019# 0.0112f
C8464 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT 0.122f
C8465 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.654f
C8466 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_31661_10099# 0.00372f
C8467 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 0.00602f
C8468 CLK a_44123_n1146# 0.00939f
C8469 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 3.08e-20
C8470 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_48832_n1102# 0.0114f
C8471 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT 2.81e-20
C8472 VDD90 F1 0.141f
C8473 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT 0.00543f
C8474 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 0.109f
C8475 F2 dec3x8_ibr_mag_0.and_3_ibr_5.nand3_mag_ibr_0.OUT 9.78e-19
C8476 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_37237_n8887# 0.0059f
C8477 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 a_51604_10154# 0.00789f
C8478 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_51239_n5724# 0.0059f
C8479 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.0622f
C8480 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 m3_20882_n11188# 0.00118f
C8481 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_22258_n2930# 1.17e-20
C8482 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.0592f
C8483 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 0.25f
C8484 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K 6.19e-20
C8485 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 5.32e-19
C8486 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_50111_n5768# 0.0732f
C8487 Vdiv90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 9e-19
C8488 Vdiv108 a_45969_n2199# 7.51e-19
C8489 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.338f
C8490 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.313f
C8491 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN 0.00279f
C8492 a_22620_n9884# m3_20882_n11188# 2.92e-19
C8493 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 a_29618_11196# 0.0101f
C8494 CLK CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 1.05e-19
C8495 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 0.0655f
C8496 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.00169f
C8497 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0454f
C8498 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB 7.08e-20
C8499 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 a_45039_n5176# 0.00859f
C8500 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.338f
C8501 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_29116_398# 0.00378f
C8502 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C8503 RST CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 0.237f
C8504 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 1.44e-19
C8505 VDD dec3x8_ibr_mag_0.and_3_ibr_0.nand3_mag_ibr_0.OUT 0.712f
C8506 RST CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.196f
C8507 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00118f
C8508 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 a_30915_n13291# 0.015f
C8509 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 0.395f
C8510 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.0725f
C8511 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 0.0635f
C8512 CLK CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.00254f
C8513 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 CLK_div_93_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.305f
C8514 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK a_35949_n8931# 0.0101f
C8515 RST CLK_div_93_mag_0.CLK_div_3_mag_0.CLK 0.0535f
C8516 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.648f
C8517 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.00975f
C8518 CLK a_24307_5062# 6.21e-19
C8519 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.019f
C8520 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 0.122f
C8521 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 7.1e-22
C8522 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_54414_6284# 2.96e-19
C8523 VDD105 F2 0.323f
C8524 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_54033_n15587# 3.33e-19
C8525 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_55132_5187# 0.0811f
C8526 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.649f
C8527 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_54187_n16728# 0.00696f
C8528 VDD108 CLK_div_108_new_mag_0.JK_FF_mag_1.QB 0.916f
C8529 VDD96 VDD99 0.665f
C8530 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 1.29e-19
C8531 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_47246_5143# 1.46e-19
C8532 RST CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN 0.022f
C8533 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.23f
C8534 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_25478_6115# 9.32e-19
C8535 VDD105 VDD108 0.0011f
C8536 RST a_51011_n18696# 1.23e-20
C8537 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 2.81e-20
C8538 VDD99 a_37328_6265# 0.0011f
C8539 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 a_46889_9057# 0.00372f
C8540 VDD96 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.751f
C8541 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 a_28574_n9876# 0.0102f
C8542 RST a_48023_10154# 0.00169f
C8543 a_53126_6240# a_53286_6240# 0.0504f
C8544 CLK_div_100_mag_0.CLK_div_10_mag_1.CLK CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.42f
C8545 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.321f
C8546 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_47196_n15629# 1.24e-20
C8547 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 0.321f
C8548 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.768f
C8549 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_45695_n17599# 0.069f
C8550 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT a_23283_n7106# 0.0203f
C8551 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 4.93e-20
C8552 a_27850_n9876# a_28010_n9876# 0.0504f
C8553 a_53844_5143# a_54004_5143# 0.0504f
C8554 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_53738_n1102# 3.25e-19
C8555 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.11f
C8556 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_33353_10099# 0.00119f
C8557 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.00164f
C8558 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_45517_5187# 0.00378f
C8559 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_24512_n18723# 4.52e-20
C8560 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK 0.209f
C8561 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT a_34896_n15539# 0.0732f
C8562 CLK_div_96_mag_0.JK_FF_mag_5.Q a_21857_810# 0.0157f
C8563 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.253f
C8564 RST a_23283_n7106# 0.00264f
C8565 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.00118f
C8566 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 5.7e-19
C8567 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_22121_11196# 0.00372f
C8568 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.28f
C8569 a_54866_n1102# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 4.52e-20
C8570 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.748f
C8571 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_22988_n1789# 0.00378f
C8572 CLK a_42083_n15712# 0.0012f
C8573 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 4.33e-19
C8574 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_53221_2768# 0.069f
C8575 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 a_31177_7256# 0.0096f
C8576 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.122f
C8577 VDD a_37168_6821# 2.21e-19
C8578 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0707f
C8579 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0854f
C8580 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 6.11e-19
C8581 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_29213_5018# 0.0733f
C8582 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB a_53216_n10117# 0.00964f
C8583 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 m3_20882_n11188# 1.85e-19
C8584 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0854f
C8585 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 9.98e-19
C8586 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 a_48944_6284# 0.069f
C8587 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.11f
C8588 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 a_50827_5143# 3.6e-22
C8589 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN 7.87e-19
C8590 RST CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 4.25e-20
C8591 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT a_53370_n9020# 4.52e-20
C8592 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.321f
C8593 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 a_51849_n1102# 9.45e-19
C8594 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 2.45e-22
C8595 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_43591_n5176# 0.0202f
C8596 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.338f
C8597 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 1.57f
C8598 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 0.0147f
C8599 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.121f
C8600 RST a_28457_n16634# 0.00273f
C8601 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_51961_6284# 0.0114f
C8602 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 m3_20882_n11188# 8.75e-19
C8603 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.187f
C8604 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 a_51034_9057# 6.43e-21
C8605 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT 0.159f
C8606 VDD108 a_50353_n9020# 3.14e-19
C8607 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 9.9e-19
C8608 a_29181_n16634# a_29341_n16634# 0.0504f
C8609 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C8610 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT a_34730_n16636# 0.0202f
C8611 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 9.64e-19
C8612 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 0.0124f
C8613 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 0.00542f
C8614 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 6.88e-21
C8615 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 9.14e-19
C8616 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 5.48e-20
C8617 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_26426_11196# 0.00695f
C8618 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 2.42f
C8619 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.0496f
C8620 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN 0.112f
C8621 Vdiv108 a_53089_n6862# 0.00335f
C8622 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 0.0409f
C8623 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 4.31e-19
C8624 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_53458_n17599# 0.00164f
C8625 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 0.338f
C8626 F1 dec3x8_ibr_mag_0.and_3_ibr_7.nand3_mag_ibr_0.OUT 0.272f
C8627 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.273f
C8628 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 CLK_div_105_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 0.00442f
C8629 RST a_48252_n9063# 7.78e-19
C8630 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 0.36f
C8631 VDD90 a_23403_10099# 3.14e-19
C8632 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_51285_n1102# 2.96e-19
C8633 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 2.11e-19
C8634 RST CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 0.00215f
C8635 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT 0.00147f
C8636 VDD99 a_28617_n16634# 7.34e-19
C8637 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 7.07e-19
C8638 CLK a_48783_n13424# 0.00487f
C8639 CLK_div_100_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_54907_297# 9.16e-20
C8640 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT m3_20882_n11188# 0.00187f
C8641 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_44799_6284# 0.0697f
C8642 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0885f
C8643 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT 0.0948f
C8644 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_43872_9057# 0.0114f
C8645 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 1.14e-20
C8646 VDD90 a_23973_11196# 0.00305f
C8647 VDD110 a_42083_n15712# 0.173f
C8648 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 9.71f
C8649 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 a_23510_n15620# 0.0178f
C8650 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.0108f
C8651 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_22461_6115# 0.00392f
C8652 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 1.32e-21
C8653 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 1.01f
C8654 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_43993_n13477# 0.0131f
C8655 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C8656 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C8657 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 0.0224f
C8658 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0894f
C8659 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 1.81e-19
C8660 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 0.00182f
C8661 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN a_52839_n5# 5.1e-20
C8662 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 8.59e-20
C8663 RST CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT 0.376f
C8664 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 3.98e-20
C8665 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.00539f
C8666 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT a_51040_10154# 0.0203f
C8667 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 6.57e-19
C8668 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.105f
C8669 VDD93 a_26343_n7107# 0.00503f
C8670 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.395f
C8671 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB 1.96f
C8672 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 3.28e-19
C8673 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.442f
C8674 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 1.5e-20
C8675 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 Vdiv110 0.00131f
C8676 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0209f
C8677 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00391f
C8678 VDD99 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 0.0448f
C8679 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 a_25646_n17626# 0.00789f
C8680 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_47902_n6273# 0.069f
C8681 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 a_45363_6284# 6.06e-21
C8682 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 a_29214_n6271# 0.00943f
C8683 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 a_34730_n16636# 0.00335f
C8684 VDD100 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 0.0983f
C8685 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 0.321f
C8686 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 a_47810_5143# 3.6e-22
C8687 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT a_54658_n9064# 0.0203f
C8688 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.121f
C8689 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.298f
C8690 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 a_51015_7381# 0.0105f
C8691 RST a_29208_10099# 3.96e-19
C8692 CLK CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.471f
C8693 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 7.36e-21
C8694 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.121f
C8695 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.0435f
C8696 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT 0.0622f
C8697 VDD99 a_23948_n13382# 0.165f
C8698 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.0685f
C8699 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 1.16f
C8700 VDD100 a_53014_n1146# 2.21e-19
C8701 CLK_div_108_new_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 6.02e-20
C8702 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_25646_n17626# 1.46e-19
C8703 VDD108 a_46246_n10116# 0.00149f
C8704 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_43793_n10116# 0.069f
C8705 a_26814_1919# CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 3.13e-20
C8706 a_50150_n15627# a_50310_n15627# 0.0504f
C8707 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_26760_5062# 0.00378f
C8708 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 2.97e-20
C8709 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.647f
C8710 RST a_31346_5018# 0.00186f
C8711 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 6.64e-19
C8712 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 a_53008_n2243# 2.55e-20
C8713 VDD93 a_22460_n9884# 2.21e-19
C8714 VDD110 a_54597_n15587# 3.14e-19
C8715 a_50868_n16724# a_51028_n16724# 0.0504f
C8716 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.122f
C8717 a_50204_2768# Vdiv110 6.25e-19
C8718 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 a_28552_354# 2.79e-20
C8719 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 1.17e-19
C8720 VDD110 a_54751_n16684# 3.14e-19
C8721 F2 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.00117f
C8722 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT a_50353_n9020# 4.52e-20
C8723 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_40408_n9984# 0.069f
C8724 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 a_32070_5018# 3.6e-22
C8725 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_39690_n8887# 0.0697f
C8726 CLK_div_105_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_105_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.11f
C8727 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.529f
C8728 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT 0.0343f
C8729 Vdiv93 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 3.8e-19
C8730 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT 0.338f
C8731 a_47424_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 1.5e-20
C8732 a_47988_n17599# a_48148_n17599# 0.0504f
C8733 CLK a_51205_n7921# 0.0103f
C8734 RST a_45081_n10160# 0.00218f
C8735 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_48944_6284# 0.0114f
C8736 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.0917f
C8737 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 0.394f
C8738 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 2.57f
C8739 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 0.188f
C8740 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0576f
C8741 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_53464_n18696# 0.00939f
C8742 RST CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0759f
C8743 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 a_29623_6159# 6.06e-21
C8744 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 2.42f
C8745 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 0.654f
C8746 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.0635f
C8747 CLK CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.00364f
C8748 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C8749 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_23409_11196# 9.1e-19
C8750 CLK_div_96_mag_0.JK_FF_mag_2.QB a_27342_n1855# 0.0114f
C8751 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.739f
C8752 CLK_div_96_mag_0.JK_FF_mag_0.QB CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.0592f
C8753 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.274f
C8754 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN 0.00668f
C8755 VDD a_37999_280# 0.00444f
C8756 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT a_36873_280# 0.0964f
C8757 RST CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 0.133f
C8758 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_36178_n16592# 0.00964f
C8759 CLK_div_96_mag_0.JK_FF_mag_3.Q a_25535_354# 0.00939f
C8760 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_33898_n18723# 0.069f
C8761 VDD96 F2 0.221f
C8762 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB a_45235_n9063# 1.86e-20
C8763 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C8764 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 4.39e-19
C8765 CLK a_43963_n1146# 0.0101f
C8766 VDD105 dec3x8_ibr_mag_0.and_3_ibr_5.nand3_mag_ibr_0.OUT 2.54e-21
C8767 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_48268_n1102# 2.96e-19
C8768 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 3.09e-19
C8769 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_36673_n8887# 0.0697f
C8770 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.00975f
C8771 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.233f
C8772 a_35454_n16636# a_35614_n16636# 0.0504f
C8773 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 a_51040_10154# 0.0102f
C8774 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.768f
C8775 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_50675_n5724# 0.0697f
C8776 RST CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT 0.00702f
C8777 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.VOUT 3.56e-19
C8778 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.00384f
C8779 Vdiv105 a_35184_880# 0.00347f
C8780 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_49951_n5768# 0.0203f
C8781 a_33405_7558# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 3.02e-19
C8782 Vdiv108 a_45405_n2199# 7.3e-19
C8783 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_45815_n1102# 0.00118f
C8784 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 a_27496_n2952# 0.00372f
C8785 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 3.4e-19
C8786 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 1.32e-19
C8787 a_30336_10099# a_30496_10099# 0.0504f
C8788 CLK a_29801_1733# 1.99e-19
C8789 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 a_29054_11196# 0.00859f
C8790 a_22460_n9884# m3_20882_n11188# 2.92e-19
C8791 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 0.133f
C8792 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 1.59e-19
C8793 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K a_28463_n15537# 0.00472f
C8794 CLK_div_100_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 4.42e-19
C8795 RST CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0106f
C8796 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 3.49e-19
C8797 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 1.48e-19
C8798 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_28552_354# 0.0732f
C8799 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT 7.24e-19
C8800 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 a_25535_354# 3.13e-20
C8801 CLK_div_108_new_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_48023_n7840# 3.25e-19
C8802 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 0.296f
C8803 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 2.86e-19
C8804 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 a_30210_n13332# 5.19e-20
C8805 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT 0.647f
C8806 VDD105 a_48747_10154# 0.0132f
C8807 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_28817_n18723# 1.09e-20
C8808 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_30469_n16590# 0.0811f
C8809 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT a_51641_n9064# 0.0203f
C8810 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.25f
C8811 a_32070_5018# a_32230_5018# 0.0504f
C8812 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_26183_n7107# 0.00119f
C8813 CLK a_23743_5062# 6.02e-19
C8814 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.159f
C8815 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 0.00718f
C8816 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 1.36e-19
C8817 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_53850_6284# 3.25e-19
C8818 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_53738_n1102# 0.00378f
C8819 F0 a_36873_280# 2.62e-19
C8820 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT 3.84e-20
C8821 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 Vdiv100 3.1e-22
C8822 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_29834_n699# 0.00378f
C8823 VDD110 a_47430_n18696# 2.66e-19
C8824 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_54568_5187# 0.00964f
C8825 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_53469_n15631# 0.00392f
C8826 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0622f
C8827 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_54027_n16728# 0.00695f
C8828 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.00384f
C8829 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 Vdiv110 0.00435f
C8830 RST a_29708_n8735# 6.56e-19
C8831 a_47492_n5176# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.00696f
C8832 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 1.32e-19
C8833 CLK_div_96_mag_0.JK_FF_mag_3.Q a_30589_n2952# 0.0157f
C8834 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_25318_6115# 0.00876f
C8835 a_29270_n743# CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 3.1e-20
C8836 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 0.116f
C8837 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.266f
C8838 CLK CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.IN2 6.62e-20
C8839 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 0.343f
C8840 VDD99 a_37168_6265# 0.00101f
C8841 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 0.0576f
C8842 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 a_28010_n9876# 0.00789f
C8843 RST a_47863_10154# 0.00186f
C8844 VDD96 a_25532_3016# 3.14e-19
C8845 CLK CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 1.48e-20
C8846 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.0072f
C8847 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_47036_n15629# 1.59e-20
C8848 VDD99 a_31733_n19822# 5.92e-19
C8849 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT a_23123_n7106# 0.0732f
C8850 F2 mux_8x1_ibr_0.mux_2x1_ibr_0.I0 4.25e-19
C8851 VDD Vdiv96 0.535f
C8852 CLK_div_105_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 4.39e-19
C8853 CLK_div_96_mag_0.JK_FF_mag_0.Q a_26214_n1855# 6.43e-21
C8854 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_27939_n17626# 8.64e-19
C8855 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 0.0568f
C8856 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_53174_n1146# 0.00486f
C8857 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_32789_10099# 1.43e-19
C8858 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00808f
C8859 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 0.12f
C8860 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_44953_5143# 0.0733f
C8861 VDD mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.461f
C8862 RST CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.107f
C8863 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN a_33812_n13270# 2.31e-19
C8864 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT a_34736_n15539# 0.0203f
C8865 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.391f
C8866 CLK CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 1.05e-19
C8867 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 Vdiv100 0.282f
C8868 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_23552_n1789# 0.0059f
C8869 RST a_46259_n17599# 0.00138f
C8870 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB 0.0378f
C8871 RST a_23123_n7106# 0.00204f
C8872 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 0.121f
C8873 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 1.83e-19
C8874 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.00205f
C8875 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_22424_n1833# 0.0732f
C8876 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_52657_2768# 0.00372f
C8877 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.0995f
C8878 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 1.33f
C8879 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.00739f
C8880 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_29053_5018# 0.0203f
C8881 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB a_52652_n10117# 0.0811f
C8882 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 0.00975f
C8883 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.122f
C8884 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.0835f
C8885 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 a_48380_6284# 6.06e-21
C8886 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 0.0881f
C8887 VDD mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 1.35f
C8888 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 a_50263_5143# 0.00166f
C8889 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 5.25e-20
C8890 F1 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT 0.107f
C8891 a_39580_6821# F0 2.63e-19
C8892 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 a_51285_n1102# 6.06e-21
C8893 CLK CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 0.0132f
C8894 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 3.38e-19
C8895 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 2.71e-21
C8896 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_39120_n10028# 1.46e-19
C8897 F2 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 1.23f
C8898 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_51397_6284# 2.96e-19
C8899 VDD108 a_49789_n9020# 3.56e-19
C8900 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 8.16e-20
C8901 CLK_div_96_mag_0.JK_FF_mag_0.Q CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.41f
C8902 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 0.122f
C8903 VDD108 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 0.165f
C8904 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB 0.199f
C8905 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.441f
C8906 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_26266_11196# 0.00696f
C8907 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 9.12e-19
C8908 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_53298_n17599# 0.00117f
C8909 F0 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 0.136f
C8910 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_26099_398# 0.00378f
C8911 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00252f
C8912 F1 a_39580_6265# 0.0112f
C8913 CLK a_54033_n15587# 6.43e-21
C8914 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_50447_n18696# 0.00939f
C8915 CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 3.81e-19
C8916 RST a_48092_n9063# 6.43e-19
C8917 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.23f
C8918 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00157f
C8919 RST CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN 0.0149f
C8920 VDD90 a_22839_10099# 3.14e-19
C8921 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 2.62e-19
C8922 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_50721_n1102# 3.25e-19
C8923 VDD99 a_28457_n16634# 9.56e-19
C8924 CLK_div_96_mag_0.JK_FF_mag_5.Q a_22418_n2930# 0.00164f
C8925 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN a_44061_n15627# 1.03e-20
C8926 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_28823_n17626# 0.0202f
C8927 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.338f
C8928 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0854f
C8929 VDD93 F1 0.369f
C8930 VDD90 a_23409_11196# 2.21e-19
C8931 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_51438_n15583# 4.52e-20
C8932 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 0.0404f
C8933 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0622f
C8934 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_25640_n18723# 0.00392f
C8935 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.00116f
C8936 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C8937 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.233f
C8938 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.529f
C8939 CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 7.24e-19
C8940 CLK_div_90_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN a_30060_9000# 0.069f
C8941 Vdiv100 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT 0.00186f
C8942 RST a_44413_n18696# 7.81e-19
C8943 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT a_50880_10154# 0.0733f
C8944 F1 F0 3.15f
C8945 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C8946 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT 0.338f
C8947 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.346f
C8948 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 5.98e-20
C8949 a_40375_n7552# CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.132f
C8950 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 0.01f
C8951 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 a_25082_n17626# 0.0102f
C8952 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 6.69e-19
C8953 RST CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.183f
C8954 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 a_47246_5143# 0.00166f
C8955 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT a_54498_n9064# 0.0732f
C8956 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_54182_n17599# 2.88e-20
C8957 CLK CLK_div_96_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0023f
C8958 RST a_28644_10099# 3.96e-19
C8959 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_0.OUT 0.122f
C8960 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_50105_n6865# 9.44e-21
C8961 RST CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 0.00103f
C8962 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0286f
C8963 VDD100 a_51849_n1102# 3.56e-19
C8964 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 5.32e-19
C8965 a_47723_574# CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 2.48e-19
C8966 CLK_div_93_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 0.124f
C8967 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 2.34e-19
C8968 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 7.24e-19
C8969 VDD96 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.746f
C8970 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_43229_n10116# 0.00372f
C8971 VDD108 a_45241_n10160# 0.00743f
C8972 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 0.878f
C8973 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_26196_5018# 0.0733f
C8974 CLK CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.00302f
C8975 a_37328_6265# dec3x8_ibr_mag_0.and_3_ibr_5.nand3_mag_ibr_0.OUT 0.0779f
C8976 RST a_30341_5062# 9.66e-19
C8977 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.122f
C8978 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 a_52003_n2199# 0.0157f
C8979 RST a_54947_n5721# 3.75e-19
C8980 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_30244_398# 0.012f
C8981 VDD110 a_54033_n15587# 3.14e-19
C8982 a_49640_2768# Vdiv110 6.45e-19
C8983 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN 0.0275f
C8984 CLK CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 7.07e-21
C8985 a_51193_n19793# CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.069f
C8986 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.343f
C8987 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 a_31506_5018# 1.86e-20
C8988 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C8989 VDD108 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1f
C8990 VDD110 a_48623_n13424# 5.08e-19
C8991 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_54004_5143# 2.88e-20
C8992 a_47264_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 1.17e-20
C8993 RST a_44517_n10160# 0.00212f
C8994 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.109f
C8995 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_48380_6284# 2.96e-19
C8996 RST CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 0.169f
C8997 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 4.95e-20
C8998 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_53304_n18696# 0.0101f
C8999 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_25800_n18723# 1.86e-20
C9000 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 7.24e-19
C9001 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 1.93e-20
C9002 CLK CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.00673f
C9003 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 2.51e-19
C9004 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.487f
C9005 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_45927_6284# 0.00118f
C9006 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 0.0529f
C9007 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_23249_11196# 2.88e-20
C9008 CLK_div_96_mag_0.JK_FF_mag_2.QB a_26778_n1855# 2.96e-19
C9009 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 a_43826_n7684# 0.0134f
C9010 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 3.25e-20
C9011 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 1.08f
C9012 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 7.11e-19
C9013 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_35614_n16636# 0.00696f
C9014 VDD105 VDD96 0.059f
C9015 VDD110 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 2.3e-20
C9016 CLK_div_96_mag_0.JK_FF_mag_3.Q a_25375_354# 0.0101f
C9017 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_33334_n18723# 0.00372f
C9018 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 0.392f
C9019 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB a_45075_n9063# 1.41e-20
C9020 RST CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 9.24e-20
C9021 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 4.52e-20
C9022 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.0635f
C9023 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_47704_n1102# 3.25e-19
C9024 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.642f
C9025 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_47492_n5176# 8.64e-19
C9026 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 a_50880_10154# 0.0101f
C9027 CLK CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 1.31f
C9028 VDD99 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 1.08e-20
C9029 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 a_28268_n6266# 0.0108f
C9030 a_33245_7558# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 9.21e-20
C9031 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0343f
C9032 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT 0.573f
C9033 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB 0.92f
C9034 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0334f
C9035 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.321f
C9036 Vdiv108 a_44841_n2243# 6.67e-19
C9037 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_45251_n1102# 0.011f
C9038 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 a_26932_n2952# 0.069f
C9039 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 0.00393f
C9040 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 8.87e-19
C9041 a_21896_n9884# m3_20882_n11188# 6.94e-19
C9042 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 a_28490_11196# 0.0157f
C9043 a_29208_10099# CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 4.9e-20
C9044 a_48587_10154# a_48747_10154# 0.0504f
C9045 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 a_37999_880# 2.44e-19
C9046 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_53850_6284# 0.00378f
C9047 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_50875_n2243# 2.88e-20
C9048 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 1.5e-20
C9049 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 1.12e-19
C9050 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0215f
C9051 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_28392_354# 0.0203f
C9052 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 4.08f
C9053 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 6.69e-19
C9054 a_28463_n15537# a_28623_n15537# 0.0504f
C9055 a_50903_n5# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 2.36e-22
C9056 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 a_30050_n13332# 3.35e-20
C9057 VDD105 a_48587_10154# 0.00891f
C9058 a_51803_n5724# CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 4.52e-20
C9059 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN a_53129_n19793# 5.1e-20
C9060 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 5.18e-20
C9061 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_28657_n18723# 8.77e-21
C9062 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_29905_n16590# 0.00964f
C9063 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT a_51481_n9064# 0.0732f
C9064 a_24784_n8778# a_24944_n8778# 0.0504f
C9065 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_40818_n8887# 0.00118f
C9066 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.IN1 0.728f
C9067 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 6.62e-20
C9068 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 2.11e-19
C9069 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_25619_n7107# 1.43e-19
C9070 CLK a_23179_5018# 5.65e-19
C9071 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_53286_6240# 0.00486f
C9072 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_53174_n1146# 0.0732f
C9073 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 1.99e-19
C9074 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_29270_n743# 0.0733f
C9075 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_54004_5143# 0.00696f
C9076 VDD110 a_47270_n18696# 3.78e-19
C9077 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 2.37f
C9078 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.JK_FF_mag_0.Q 2.64e-20
C9079 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 9.75e-19
C9080 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.768f
C9081 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN a_43826_n7684# 0.132f
C9082 a_29834_n699# CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 4.58e-20
C9083 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT 0.163f
C9084 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.16f
C9085 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_48056_n5176# 0.00378f
C9086 a_47332_n5176# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.00695f
C9087 RST a_29144_n8735# 6.56e-19
C9088 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 9.73e-19
C9089 CLK_div_96_mag_0.JK_FF_mag_3.Q a_30025_n2952# 0.00859f
C9090 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 2.84e-20
C9091 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 8.76e-20
C9092 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 2.08e-20
C9093 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 0.904f
C9094 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.00183f
C9095 VDD93 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 4.37e-19
C9096 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.00356f
C9097 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 3.55e-20
C9098 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 a_27850_n9876# 0.00335f
C9099 VDD96 a_24968_3016# 3.14e-19
C9100 RST a_47299_10154# 9.41e-19
C9101 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 a_25420_n13385# 0.00589f
C9102 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 dec3x8_ibr_mag_0.and_3_ibr_5.nand3_mag_ibr_0.OUT 0.00136f
C9103 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_45753_n15583# 0.0114f
C9104 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT a_22559_n7106# 0.00378f
C9105 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00158f
C9106 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 8.64e-20
C9107 RST CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 0.169f
C9108 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 2.81e-20
C9109 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.122f
C9110 CLK_div_96_mag_0.JK_FF_mag_0.Q a_25650_n1899# 0.00939f
C9111 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 CLK_div_108_new_mag_0.JK_FF_mag_1.QB 2.61e-19
C9112 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_53014_n1146# 0.00111f
C9113 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_32225_10099# 0.011f
C9114 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN 8.99e-19
C9115 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN 0.00102f
C9116 RST CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 0.337f
C9117 VDD Vdiv108 0.508f
C9118 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.0432f
C9119 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0622f
C9120 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_44793_5143# 0.0203f
C9121 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_37801_n8887# 0.00118f
C9122 VDD96 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_4.IN2 0.391f
C9123 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN a_33652_n13270# 3.59e-19
C9124 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 7.16e-20
C9125 RST a_45695_n17599# 0.0015f
C9126 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_22988_n1789# 0.0697f
C9127 RST a_22559_n7106# 6.28e-19
C9128 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT 0.649f
C9129 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 0.124f
C9130 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.233f
C9131 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_27334_n16588# 0.0811f
C9132 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.0877f
C9133 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 a_21431_n7106# 4.52e-20
C9134 a_40375_n7552# CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.00168f
C9135 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 0.235f
C9136 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_22264_n1833# 0.0203f
C9137 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 a_46755_574# 0.0084f
C9138 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 6.02e-20
C9139 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 0.329f
C9140 RST CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.196f
C9141 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_28489_5018# 1.5e-20
C9142 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C9143 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.768f
C9144 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.IN1 m3_20882_n11188# 0.00979f
C9145 a_27180_n15491# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 4.52e-20
C9146 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_28817_n18723# 0.0203f
C9147 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN a_22544_n13819# 0.069f
C9148 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0611f
C9149 RST CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.0148f
C9150 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0592f
C9151 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 0.276f
C9152 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 a_50103_5143# 0.00119f
C9153 a_39420_6821# F0 5.62e-19
C9154 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 1.03f
C9155 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN 9.25e-19
C9156 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB 9.89e-20
C9157 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.122f
C9158 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_54022_n17599# 3.6e-22
C9159 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 6.28e-19
C9160 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.338f
C9161 VDD105 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 0.0665f
C9162 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 m3_20882_n11188# 1.73e-20
C9163 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.00975f
C9164 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 3.38e-20
C9165 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.0894f
C9166 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_30317_n18723# 4.52e-20
C9167 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.742f
C9168 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT a_47994_n18696# 0.00378f
C9169 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_50833_6284# 3.25e-19
C9170 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K a_53309_n15631# 0.00472f
C9171 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_52115_5187# 0.0811f
C9172 VDD108 a_48252_n9063# 5.99e-19
C9173 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 a_49906_9057# 9.26e-19
C9174 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 0.0105f
C9175 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0635f
C9176 Vdiv100 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 0.0189f
C9177 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.0445f
C9178 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT 0.122f
C9179 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_24270_n2886# 0.00372f
C9180 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.739f
C9181 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 2.98e-19
C9182 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_25702_11196# 0.00964f
C9183 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 0.0622f
C9184 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.206f
C9185 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.398f
C9186 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 0.0016f
C9187 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.0763f
C9188 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 0.0501f
C9189 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.198f
C9190 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 0.159f
C9191 F0 a_35747_280# 6.89e-19
C9192 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_25535_354# 0.0732f
C9193 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 1.39e-19
C9194 F1 a_39420_6265# 0.00741f
C9195 CLK a_53469_n15631# 0.00939f
C9196 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_50287_n18696# 0.0101f
C9197 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 a_26811_n17626# 2.34e-20
C9198 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 6.91e-20
C9199 RST a_47528_n9019# 2.23e-19
C9200 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 0.0529f
C9201 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN 2.86e-19
C9202 VDD90 a_22275_10099# 3.56e-19
C9203 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C9204 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C9205 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_50157_n1146# 0.00392f
C9206 a_29213_n7028# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 3.66e-20
C9207 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 5.69e-19
C9208 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 2.03e-20
C9209 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00254f
C9210 CLK_div_96_mag_0.JK_FF_mag_5.Q a_22258_n2930# 0.00117f
C9211 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN a_43901_n15627# 1.29e-20
C9212 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_28663_n17626# 0.0731f
C9213 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 8.93e-19
C9214 a_23249_11196# a_23409_11196# 0.0504f
C9215 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_50874_n15583# 0.0195f
C9216 RST a_50721_n1102# 1.23e-20
C9217 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.00102f
C9218 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_25076_n18723# 1.75e-19
C9219 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_51592_n16680# 0.00378f
C9220 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 7.14e-19
C9221 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 2.76e-19
C9222 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_54615_9057# 0.00119f
C9223 RST a_44253_n18696# 9.37e-19
C9224 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT a_50316_10154# 0.00378f
C9225 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_29087_8532# 1.4e-19
C9226 VDD93 a_25619_n7107# 3.14e-19
C9227 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 a_47341_1671# 6.06e-21
C9228 CLK_div_105_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 0.00442f
C9229 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 0.00238f
C9230 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 0.647f
C9231 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.0343f
C9232 a_22982_n2930# a_23142_n2930# 0.0504f
C9233 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.652f
C9234 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN 1.03e-19
C9235 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN 0.108f
C9236 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 a_24922_n17626# 0.0101f
C9237 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.359f
C9238 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1.01f
C9239 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 a_44235_6240# 2.79e-20
C9240 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN m3_20882_n11188# 1.63e-21
C9241 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 6.62e-20
C9242 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_31512_6115# 1.41e-20
C9243 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 a_47086_5143# 0.001f
C9244 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT a_53934_n9020# 0.00378f
C9245 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_54022_n17599# 9.1e-19
C9246 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_53487_9057# 0.069f
C9247 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_49945_n6865# 1.17e-20
C9248 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 a_33429_n15491# 0.069f
C9249 VDD100 a_51285_n1102# 3.14e-19
C9250 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.0134f
C9251 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.426f
C9252 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C9253 CLK_div_108_new_mag_0.JK_FF_mag_1.QB CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.25f
C9254 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 0.0127f
C9255 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 0.00115f
C9256 VDD108 a_45081_n10160# 0.00305f
C9257 Vdiv110 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 0.075f
C9258 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 1.83e-20
C9259 a_37168_6265# dec3x8_ibr_mag_0.and_3_ibr_5.nand3_mag_ibr_0.OUT 0.0249f
C9260 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_26036_5018# 0.0203f
C9261 a_53014_n1146# a_53174_n1146# 0.0504f
C9262 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 4.36e-20
C9263 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 8.27e-19
C9264 RST a_29777_5062# 9.41e-19
C9265 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 0.026f
C9266 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.122f
C9267 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 a_51439_n2199# 0.00859f
C9268 RST a_54383_n5721# 3.75e-19
C9269 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 1.17e-19
C9270 VDD93 a_21736_n9884# 0.00108f
C9271 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_29680_398# 2.96e-19
C9272 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.198f
C9273 CLK_div_108_new_mag_0.JK_FF_mag_0.QB CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.198f
C9274 VDD110 a_54027_n16728# 2.21e-19
C9275 a_23948_n13382# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 0.132f
C9276 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 a_31346_5018# 2.55e-20
C9277 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT 0.306f
C9278 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.199f
C9279 VDD110 a_41117_n13911# 3.14e-19
C9280 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 8.58e-20
C9281 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_53844_5143# 9.1e-19
C9282 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 0.00393f
C9283 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00397f
C9284 RST a_44357_n10160# 0.00204f
C9285 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00545f
C9286 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 3.53e-19
C9287 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_47816_6284# 3.25e-19
C9288 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_25640_n18723# 1.41e-20
C9289 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 1.33e-20
C9290 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_52139_n18696# 9.45e-19
C9291 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 4.08f
C9292 a_38294_6821# a_38454_6821# 0.0504f
C9293 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_45363_6284# 0.011f
C9294 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.25f
C9295 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 9.98e-19
C9296 CLK_div_96_mag_0.JK_FF_mag_2.QB a_26214_n1855# 3.33e-19
C9297 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT 0.647f
C9298 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB a_35454_n16636# 0.00695f
C9299 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K 0.00102f
C9300 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 8.94e-19
C9301 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 6.22e-20
C9302 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0622f
C9303 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 9.85e-20
C9304 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_47140_n1146# 0.00392f
C9305 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.178f
C9306 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 2.18e-21
C9307 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 a_37328_6821# 0.00194f
C9308 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 a_50316_10154# 0.00859f
C9309 RST CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.21f
C9310 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C9311 RST CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 0.11f
C9312 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 a_39402_n7788# 0.01f
C9313 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 5.18e-20
C9314 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.64f
C9315 CLK CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 0.00391f
C9316 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 5.05f
C9317 VDD Vdiv93 0.237f
C9318 CLK_div_96_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 6.02e-20
C9319 Vdiv108 a_44681_n2243# 6.67e-19
C9320 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_44687_n1102# 1.43e-19
C9321 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 2.04e-19
C9322 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.306f
C9323 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 6.24e-20
C9324 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 a_30164_n7017# 9.22e-21
C9325 CLK_div_108_new_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 0.00559f
C9326 a_21736_n9884# m3_20882_n11188# 6.94e-19
C9327 CLK CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.00481f
C9328 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_0.OUT a_29307_n1855# 0.00378f
C9329 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.00356f
C9330 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 1.54e-21
C9331 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 a_37436_880# 1.04e-19
C9332 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_53286_6240# 0.0732f
C9333 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_50715_n2243# 9.1e-19
C9334 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 3.21e-20
C9335 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_25806_n17626# 1.17e-20
C9336 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00183f
C9337 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_0.OUT CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 5.51e-20
C9338 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 a_36873_n1822# 0.00372f
C9339 VDD100 a_47723_574# 6e-19
C9340 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 CLK_div_90_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00311f
C9341 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 0.622f
C9342 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 7.14e-19
C9343 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 1.98e-19
C9344 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 a_22544_n13819# 0.00544f
C9345 VDD105 a_48023_10154# 0.00123f
C9346 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 2.19f
C9347 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_29341_n16634# 0.00696f
C9348 CLK_div_96_mag_0.JK_FF_mag_2.QB CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.28f
C9349 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT a_50917_n9020# 0.00378f
C9350 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 a_28580_n8735# 6.43e-21
C9351 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_40254_n8887# 0.011f
C9352 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 2.34f
C9353 RST CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.0222f
C9354 VDD mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 0.46f
C9355 CLK a_23019_5018# 5.65e-19
C9356 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_25055_n7107# 0.011f
C9357 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0129f
C9358 RST CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0353f
C9359 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 0.235f
C9360 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00776f
C9361 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_53126_6240# 0.00111f
C9362 RST CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0134f
C9363 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_53014_n1146# 0.0203f
C9364 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 9.8e-19
C9365 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_29110_n743# 0.0203f
C9366 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_53844_5143# 0.00695f
C9367 VDD110 a_46105_n18696# 3.56e-19
C9368 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT 0.0693f
C9369 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0622f
C9370 RST a_28580_n8735# 5.43e-19
C9371 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0854f
C9372 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_26965_n18723# 4.52e-20
C9373 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0951f
C9374 CLK_div_96_mag_0.JK_FF_mag_3.Q a_29461_n2996# 0.0101f
C9375 VDD96 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 0.0687f
C9376 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.739f
C9377 VDD90 VDD93 0.399f
C9378 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 3.85e-20
C9379 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 0.66f
C9380 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_32230_5018# 2.88e-20
C9381 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB 0.103f
C9382 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN 0.107f
C9383 RST CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0202f
C9384 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00262f
C9385 a_33204_6159# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 4.52e-20
C9386 RST a_46735_10154# 9.66e-19
C9387 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_45189_n15583# 2.96e-19
C9388 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT a_29187_n15493# 0.00378f
C9389 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 a_37328_6265# 3.18e-19
C9390 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 a_28268_n6266# 0.00389f
C9391 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_50441_n17599# 3.66e-20
C9392 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C9393 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT 0.0622f
C9394 CLK CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.242f
C9395 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 1.32f
C9396 CLK_div_96_mag_0.JK_FF_mag_0.Q a_25490_n1899# 0.0101f
C9397 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 4.16f
C9398 VDD90 F0 0.168f
C9399 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.103f
C9400 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0779f
C9401 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_51849_n1102# 7.4e-19
C9402 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 2.62e-20
C9403 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT a_26206_n16632# 2.88e-20
C9404 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_31661_10099# 0.00118f
C9405 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 0.36f
C9406 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_43993_n13477# 8.64e-19
C9407 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.274f
C9408 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_37237_n8887# 0.011f
C9409 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_44229_5143# 1.5e-20
C9410 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C9411 CLK_div_100_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 0.00442f
C9412 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 0.0379f
C9413 CLK_div_93_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 2.34e-19
C9414 RST a_21995_n7106# 6.04e-19
C9415 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 3.81e-19
C9416 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT 0.00669f
C9417 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.122f
C9418 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 0.048f
C9419 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_26770_n16588# 0.00964f
C9420 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 2.06e-19
C9421 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 0.139f
C9422 CLK CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 1.29e-19
C9423 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 3.46e-19
C9424 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_28329_5018# 1.17e-20
C9425 Vdiv108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K 0.0613f
C9426 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 6.04e-21
C9427 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_28657_n18723# 0.0732f
C9428 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 0.25f
C9429 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 a_51598_9057# 0.00119f
C9430 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.36f
C9431 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 a_47252_6240# 2.79e-20
C9432 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.CLK 0.0036f
C9433 RST a_32750_n7675# 0.00703f
C9434 Vdiv110 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.00782f
C9435 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 a_49098_5187# 0.0157f
C9436 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 2.63f
C9437 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.VOUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00384f
C9438 RST CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 0.277f
C9439 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 8.94e-19
C9440 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_33204_6159# 0.0114f
C9441 CLK CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.235f
C9442 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_53458_n17599# 1.86e-20
C9443 RST CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN 0.0417f
C9444 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 2.07e-20
C9445 CLK_div_96_mag_0.JK_FF_mag_0.Q CLK_div_96_mag_0.JK_FF_mag_2.Q 0.155f
C9446 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_50269_6240# 0.00392f
C9447 RST a_43831_7266# 0.00198f
C9448 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.359f
C9449 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_51551_5187# 0.00964f
C9450 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C9451 VDD108 a_48092_n9063# 2.65e-19
C9452 Vdiv100 a_37999_280# 4.15e-20
C9453 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 5.95e-20
C9454 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K a_53303_n16728# 8.64e-19
C9455 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_23706_n2886# 0.069f
C9456 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_25138_11196# 0.0811f
C9457 CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 a_31733_n19822# 7.48e-20
C9458 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.359f
C9459 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.69f
C9460 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00118f
C9461 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0622f
C9462 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 1.54e-19
C9463 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.0161f
C9464 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_25375_354# 0.0203f
C9465 CLK a_53309_n15631# 0.0101f
C9466 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_49122_n18696# 0.069f
C9467 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.235f
C9468 CLK a_53463_n16728# 0.00164f
C9469 CLK_div_100_mag_0.CLK_div_10_mag_1.CLK CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 6.64e-19
C9470 RST a_46964_n9019# 0.00121f
C9471 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN a_46755_574# 0.069f
C9472 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_26778_n1855# 4.52e-20
C9473 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 8.16e-20
C9474 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 1.58e-20
C9475 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.105f
C9476 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 9e-20
C9477 RST a_25625_n6010# 8.64e-19
C9478 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00183f
C9479 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_28099_n17626# 9.1e-19
C9480 VDD90 a_22685_11196# 3.14e-19
C9481 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 0.593f
C9482 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I1 Vdiv108 0.00305f
C9483 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_24512_n18723# 2.96e-19
C9484 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0871f
C9485 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_51028_n16724# 0.0733f
C9486 VDD110 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 0.00159f
C9487 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.00166f
C9488 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_54051_9057# 1.43e-19
C9489 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.0591f
C9490 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT a_26052_n15491# 0.00378f
C9491 VDD93 a_25055_n7107# 3.14e-19
C9492 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 6.7e-19
C9493 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 a_46777_1671# 9.45e-19
C9494 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.748f
C9495 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K m3_20882_n11188# 0.00526f
C9496 CLK_div_105_mag_0.CLK_div_10_mag_1.CLK CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 1.48e-20
C9497 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.00183f
C9498 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 7.75e-19
C9499 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.00384f
C9500 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_0.OUT 0.122f
C9501 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN 0.00141f
C9502 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_29213_5018# 8.64e-19
C9503 dec3x8_ibr_mag_0.and_3_ibr_5.IN3 dec3x8_ibr_mag_0.and_3_ibr_1.nand3_mag_ibr_0.OUT 0.119f
C9504 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 a_24358_n17626# 0.00859f
C9505 VDD108 a_54947_n5721# 3.56e-19
C9506 a_39580_6265# dec3x8_ibr_mag_0.and_3_ibr_7.nand3_mag_ibr_0.OUT 0.0779f
C9507 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_0.OUT 7.24e-19
C9508 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 dec3x8_ibr_mag_0.and_3_ibr_0.nand3_mag_ibr_0.OUT 0.263f
C9509 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 9.5e-19
C9510 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0345f
C9511 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT a_45815_n1102# 2.05e-19
C9512 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_31352_6115# 1.86e-20
C9513 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.121f
C9514 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 a_46081_5187# 0.0157f
C9515 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0345f
C9516 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_53458_n17599# 0.0731f
C9517 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.122f
C9518 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 8.51e-22
C9519 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 a_26636_n8734# 4.6e-19
C9520 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.00109f
C9521 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.0175f
C9522 VDD96 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.653f
C9523 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_52923_9057# 0.00372f
C9524 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0569f
C9525 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 0.00121f
C9526 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.103f
C9527 VDD100 a_50721_n1102# 3.14e-19
C9528 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 Vdiv 0.0632f
C9529 VDD93 a_40375_n7552# 0.172f
C9530 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_24358_n17626# 0.0036f
C9531 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 0.103f
C9532 VDD a_39124_880# 0.00444f
C9533 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN 0.0758f
C9534 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 m3_20882_n11188# 0.00101f
C9535 CLK CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.268f
C9536 VDD108 a_44517_n10160# 2.21e-19
C9537 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0705f
C9538 a_37168_6265# a_37328_6265# 0.0504f
C9539 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_25472_5018# 1.5e-20
C9540 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB 0.28f
C9541 CLK_div_90_mag_0.CLK_div_10_mag_0.CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.267f
C9542 CLK_div_90_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.00117f
C9543 RST a_29213_5018# 0.00186f
C9544 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 5.11e-19
C9545 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 a_50875_n2243# 0.0101f
C9546 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C9547 RST a_53819_n5721# 4.3e-19
C9548 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_2.OUT a_26980_3016# 0.0202f
C9549 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.289f
C9550 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 0.00238f
C9551 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_29116_398# 1.75e-19
C9552 VDD110 a_53309_n15631# 2.21e-19
C9553 Vdiv96 Vdiv100 0.0715f
C9554 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 2.39f
C9555 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB 0.912f
C9556 Vdiv99 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 0.117f
C9557 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 0.00761f
C9558 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 a_30341_5062# 0.0157f
C9559 Vdiv108 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.108f
C9560 F0 dec3x8_ibr_mag_0.and_3_ibr_7.nand3_mag_ibr_0.OUT 0.354f
C9561 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 a_22711_n14504# 8.95e-19
C9562 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.JK_FF_mag_2.QB 1.61e-19
C9563 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 a_33583_n16588# 0.00372f
C9564 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_53280_5143# 0.0731f
C9565 RST CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN 0.0227f
C9566 RST a_43793_n10116# 0.00122f
C9567 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_47252_6240# 0.00392f
C9568 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_4.IN2 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT 0.122f
C9569 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_49098_5187# 0.0811f
C9570 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_51575_n18696# 6.06e-21
C9571 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.00127f
C9572 RST CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 1.03f
C9573 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.251f
C9574 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 0.0496f
C9575 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_44799_6284# 1.43e-19
C9576 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 0.386f
C9577 CLK_div_96_mag_0.JK_FF_mag_2.QB a_25650_n1899# 0.00392f
C9578 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK 0.25f
C9579 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT 0.257f
C9580 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.0592f
C9581 Vdiv100 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 0.0115f
C9582 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.064f
C9583 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB a_51040_10154# 0.00695f
C9584 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0306f
C9585 dec3x8_ibr_mag_0.and_3_ibr_0.nand3_mag_ibr_0.OUT a_36202_6821# 0.0779f
C9586 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 a_37168_6821# 0.00182f
C9587 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 a_49752_10154# 0.0157f
C9588 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT Vdiv110 0.00521f
C9589 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.113f
C9590 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN a_30165_n6282# 1.05e-20
C9591 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0274f
C9592 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.125f
C9593 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.343f
C9594 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_29871_n1855# 0.0059f
C9595 Vdiv108 a_44117_n2243# 0.00158f
C9596 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_44123_n1146# 0.00119f
C9597 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 1.4e-20
C9598 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 9.98e-19
C9599 CLK_div_100_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 a_54866_n1102# 2.1e-20
C9600 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 a_31731_n16632# 4.66e-19
C9601 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 8.16e-20
C9602 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 4.92e-21
C9603 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00118f
C9604 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 7.08e-20
C9605 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0156f
C9606 CLK CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.00302f
C9607 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_0.OUT a_28743_n1899# 0.0732f
C9608 a_47050_n7372# CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 3.16e-19
C9609 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 a_36873_880# 2.44e-19
C9610 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 0.128f
C9611 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN 0.11f
C9612 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_53126_6240# 0.0203f
C9613 RST a_23691_9000# 5e-19
C9614 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_50151_n2243# 0.0731f
C9615 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT 0.343f
C9616 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.0881f
C9617 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 0.0222f
C9618 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 1.2e-19
C9619 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB m3_20882_n11188# 0.00404f
C9620 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 0.69f
C9621 CLK_div_108_new_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 6.11e-19
C9622 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_25646_n17626# 1.5e-20
C9623 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 2.64e-19
C9624 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 2e-19
C9625 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 6.82e-19
C9626 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 a_36310_n1822# 0.069f
C9627 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN 0.00907f
C9628 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 1f
C9629 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.122f
C9630 VDD105 a_47863_10154# 0.00101f
C9631 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.198f
C9632 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB a_29181_n16634# 0.00695f
C9633 CLK_div_96_mag_0.JK_FF_mag_3.QB a_30589_n2952# 0.0811f
C9634 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.131f
C9635 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 a_28016_n8779# 0.00939f
C9636 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_39690_n8887# 1.43e-19
C9637 RST a_28823_n17626# 0.00466f
C9638 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 a_48581_9057# 0.00119f
C9639 CLK a_22455_5018# 0.00134f
C9640 a_45899_7960# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 8.17e-21
C9641 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_24491_n7107# 0.00118f
C9642 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00617f
C9643 a_47424_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 1.46e-19
C9644 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.0496f
C9645 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 0.0635f
C9646 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_51961_6284# 7.4e-19
C9647 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0697f
C9648 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_28546_n743# 1.5e-20
C9649 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.121f
C9650 VDD110 a_45541_n18696# 3.14e-19
C9651 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 0.781f
C9652 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 0.00212f
C9653 RST a_28016_n8779# 0.00154f
C9654 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 1f
C9655 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 0.342f
C9656 CLK_div_96_mag_0.JK_FF_mag_3.Q a_29301_n2996# 0.0102f
C9657 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.36f
C9658 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_32070_5018# 9.1e-19
C9659 CLK CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 0.149f
C9660 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 a_23956_n14213# 0.00379f
C9661 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.269f
C9662 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 a_37168_6265# 5.51e-19
C9663 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT a_28623_n15537# 0.0732f
C9664 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_44625_n15583# 3.33e-19
C9665 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_23967_10099# 0.00119f
C9666 a_53120_5143# a_53280_5143# 0.0504f
C9667 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.392f
C9668 CLK_div_96_mag_0.JK_FF_mag_0.Q a_24116_n1789# 0.069f
C9669 VDD dec3x8_ibr_mag_0.and_3_ibr_6.nand3_mag_ibr_0.OUT 0.693f
C9670 VDD90 a_30187_6159# 3.56e-19
C9671 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.103f
C9672 VDD96 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT 0.999f
C9673 CLK CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 3.23e-19
C9674 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_51285_n1102# 7.4e-19
C9675 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT a_26046_n16632# 9.1e-19
C9676 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_36673_n8887# 1.43e-19
C9677 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_44069_5143# 1.17e-20
C9678 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C9679 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0622f
C9680 CLK_div_96_mag_0.JK_FF_mag_4.QB CLK_div_96_mag_0.JK_FF_mag_3.Q 3.23e-19
C9681 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 7.08e-20
C9682 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 1.64e-20
C9683 RST a_21431_n7106# 6.04e-19
C9684 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.457f
C9685 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT 0.00543f
C9686 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 7.63e-19
C9687 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 1.2f
C9688 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_45815_n1102# 0.00372f
C9689 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT 6.99e-20
C9690 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_26206_n16632# 0.00696f
C9691 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN a_31128_n7028# 8.67e-20
C9692 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0129f
C9693 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.JK_FF_mag_1.Q 0.0179f
C9694 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 4.67e-22
C9695 CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 0.0445f
C9696 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.0979f
C9697 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 0.321f
C9698 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 1.54e-19
C9699 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.00481f
C9700 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 a_51034_9057# 1.43e-19
C9701 Vdiv90 Vdiv99 1.63e-19
C9702 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_28093_n18723# 0.00378f
C9703 Vdiv105 CLK_div_105_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00258f
C9704 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 a_48534_5187# 0.00859f
C9705 RST CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.0581f
C9706 VDD93 a_23594_n8743# 3.56e-19
C9707 a_38294_6821# F0 5.62e-19
C9708 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 0.242f
C9709 a_30317_n18723# CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 4.94e-20
C9710 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 0.0582f
C9711 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_32640_6159# 2.96e-19
C9712 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 a_36742_n16592# 0.00372f
C9713 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_53298_n17599# 2.55e-20
C9714 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 7.24e-19
C9715 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0384f
C9716 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB 2.15e-19
C9717 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.122f
C9718 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 0.623f
C9719 RST a_43671_7266# 0.00189f
C9720 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_4.QB 0.28f
C9721 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I1 0.109f
C9722 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB 3.48e-19
C9723 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.103f
C9724 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_50987_5143# 0.00696f
C9725 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.122f
C9726 VDD108 a_47528_n9019# 3.14e-19
C9727 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 a_35747_880# 0.00372f
C9728 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K a_52156_n16680# 2.75e-21
C9729 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 2.01e-19
C9730 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00137f
C9731 a_28457_n16634# a_28617_n16634# 0.0504f
C9732 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.122f
C9733 a_40818_n8887# CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 4.52e-20
C9734 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK a_44407_n17599# 0.00164f
C9735 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_51652_2768# 2.81e-19
C9736 CLK a_52002_n15583# 9.36e-19
C9737 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_48558_n18696# 6.06e-21
C9738 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.177f
C9739 CLK a_53303_n16728# 0.00117f
C9740 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.313f
C9741 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 0.107f
C9742 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 0.00602f
C9743 VDD99 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 0.00152f
C9744 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT 0.00982f
C9745 RST a_46400_n9019# 0.00154f
C9746 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN 0.0549f
C9747 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_26214_n1855# 0.0202f
C9748 RST a_25465_n6010# 0.00173f
C9749 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 0.321f
C9750 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN 0.00102f
C9751 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_53973_n6862# 8.64e-19
C9752 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 1.19f
C9753 CLK_div_105_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 7.14e-19
C9754 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_33583_n16588# 0.0811f
C9755 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_27939_n17626# 2.88e-20
C9756 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 0.266f
C9757 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_32789_10099# 0.0202f
C9758 VDD90 a_22121_11196# 3.14e-19
C9759 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 1.82e-19
C9760 a_43872_9057# CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 1.54e-19
C9761 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 2.01e-19
C9762 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_44953_5143# 8.64e-19
C9763 VDD100 a_43831_7266# 0.00249f
C9764 RST CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.302f
C9765 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_23948_n18723# 0.012f
C9766 Vdiv105 F1 0.166f
C9767 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 a_39402_n7788# 7.48e-20
C9768 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.VOUT CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN 1.56e-19
C9769 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_50868_n16724# 0.0203f
C9770 CLK CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT 1.29e-19
C9771 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB 0.103f
C9772 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_53487_9057# 0.011f
C9773 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.99e-19
C9774 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT a_33812_n13270# 8.64e-19
C9775 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.237f
C9776 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_26072_n8734# 4.52e-20
C9777 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_33513_10099# 8.64e-19
C9778 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.768f
C9779 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT a_25488_n15535# 0.0732f
C9780 VDD93 a_24491_n7107# 3.56e-19
C9781 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 2.75e-19
C9782 VDD96 CLK_div_90_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 4.43e-19
C9783 CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.209f
C9784 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 0.0591f
C9785 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0854f
C9786 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 a_23794_n17626# 0.0157f
C9787 RST CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.322f
C9788 F0 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT 0.00165f
C9789 VDD108 a_54383_n5721# 3.14e-19
C9790 a_39420_6265# dec3x8_ibr_mag_0.and_3_ibr_7.nand3_mag_ibr_0.OUT 0.0249f
C9791 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 1.87e-19
C9792 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 a_45517_5187# 0.00859f
C9793 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 a_54182_n17599# 0.0101f
C9794 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_53298_n17599# 0.0202f
C9795 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_33744_n17626# 0.069f
C9796 dec3x8_ibr_mag_0.and_3_ibr_2.nand3_mag_ibr_0.OUT a_39580_6821# 3.58e-20
C9797 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.00143f
C9798 RST CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00797f
C9799 VDD100 a_50157_n1146# 2.66e-19
C9800 VDD a_38561_880# 3.14e-19
C9801 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 Vdiv110 0.00376f
C9802 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.11f
C9803 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT a_45787_574# 0.00138f
C9804 VDD99 a_35186_n18723# 5.99e-19
C9805 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.16f
C9806 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.468f
C9807 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.343f
C9808 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_25312_5018# 1.17e-20
C9809 RST a_29053_5018# 0.00169f
C9810 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_53304_n18696# 6.36e-19
C9811 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 0.128f
C9812 a_51983_7381# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 1.45e-20
C9813 RST a_53255_n5765# 0.00122f
C9814 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_2.OUT a_26820_3016# 0.0731f
C9815 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 a_50715_n2243# 0.0102f
C9816 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB 0.198f
C9817 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_28552_354# 0.00392f
C9818 VDD110 a_52002_n15583# 3.56e-19
C9819 a_50144_n16724# a_50304_n16724# 0.0504f
C9820 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 0.416f
C9821 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.289f
C9822 VDD110 a_53303_n16728# 2.21e-19
C9823 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K 0.487f
C9824 F0 a_39580_6265# 0.00168f
C9825 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 a_29777_5062# 0.00859f
C9826 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.CLK 0.00887f
C9827 Vdiv90 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.IN2 0.0686f
C9828 Vdiv100 Vdiv108 1.37f
C9829 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 a_33019_n16588# 0.069f
C9830 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.415f
C9831 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 0.149f
C9832 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_53120_5143# 0.0202f
C9833 a_47264_n17599# a_47424_n17599# 0.0504f
C9834 RST a_43229_n10116# 0.00114f
C9835 RST a_27227_398# 0.00155f
C9836 RST CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 0.0465f
C9837 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_48534_5187# 0.00964f
C9838 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.352f
C9839 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 a_27170_6159# 9.26e-19
C9840 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 3.68e-19
C9841 VDD93 F0 0.228f
C9842 a_54182_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.00696f
C9843 CLK a_28267_n7033# 2.26e-19
C9844 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_43826_n7684# 2.51e-19
C9845 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 0.642f
C9846 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_44235_6240# 0.00119f
C9847 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.00157f
C9848 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.28f
C9849 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 a_51438_n15583# 0.0059f
C9850 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.352f
C9851 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C9852 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_33513_10099# 0.0203f
C9853 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 5.08e-20
C9854 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C9855 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.106f
C9856 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 3.49e-19
C9857 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB a_51646_1671# 1.86e-20
C9858 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 a_30165_n6282# 0.00347f
C9859 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.105f
C9860 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 0.492f
C9861 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.374f
C9862 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB 3.28e-19
C9863 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00183f
C9864 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 5.79e-20
C9865 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB a_50880_10154# 0.00696f
C9866 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0346f
C9867 dec3x8_ibr_mag_0.and_3_ibr_0.nand3_mag_ibr_0.OUT a_36042_6821# 0.0249f
C9868 F1 dec3x8_ibr_mag_0.and_3_ibr_2.nand3_mag_ibr_0.OUT 8.63e-19
C9869 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.0659f
C9870 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0948f
C9871 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 3.87e-19
C9872 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 1.96f
C9873 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 4.27e-20
C9874 RST CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.00239f
C9875 a_34730_n16636# a_34890_n16636# 0.0504f
C9876 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.175f
C9877 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 0.399f
C9878 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN a_29214_n6271# 0.069f
C9879 RST CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.082f
C9880 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 0.121f
C9881 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_50447_n18696# 0.00392f
C9882 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.065f
C9883 Vdiv108 a_43957_n2243# 0.00158f
C9884 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_29307_n1855# 0.0697f
C9885 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 1.93f
C9886 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 a_31571_n16632# 6.02e-19
C9887 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 1.87e-19
C9888 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0151f
C9889 a_43826_n7684# CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 0.00168f
C9890 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 4.78e-20
C9891 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 1.17e-19
C9892 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_0.OUT a_28583_n1899# 0.0203f
C9893 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 a_36310_880# 0.00211f
C9894 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 m3_20882_n11188# 8.75e-19
C9895 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_49991_n2243# 0.0202f
C9896 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 0.983f
C9897 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0622f
C9898 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_25082_n17626# 0.0203f
C9899 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 1.59e-20
C9900 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.267f
C9901 a_28267_n7033# CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 1.91e-21
C9902 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_29213_n7028# 3.85e-20
C9903 VDD108 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.31f
C9904 VDD93 m3_20882_n11188# 0.0993f
C9905 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.IN2 1.19e-20
C9906 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_26196_5018# 8.64e-19
C9907 CLK CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 2.31f
C9908 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 8.02e-19
C9909 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0899f
C9910 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 a_29708_n8735# 0.0695f
C9911 CLK_div_96_mag_0.JK_FF_mag_2.QB CLK_div_96_mag_0.JK_FF_mag_2.Q 1.96f
C9912 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.121f
C9913 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 0.00164f
C9914 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB 6.93e-19
C9915 VDD105 a_47299_10154# 0.00152f
C9916 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.647f
C9917 CLK_div_96_mag_0.JK_FF_mag_3.QB a_30025_n2952# 0.00964f
C9918 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.121f
C9919 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.103f
C9920 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.00434f
C9921 RST CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00365f
C9922 CLK CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 3.43e-19
C9923 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 a_27856_n8779# 0.0101f
C9924 a_31346_5018# a_31506_5018# 0.0504f
C9925 RST CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 0.277f
C9926 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_39126_n8931# 0.00119f
C9927 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 5.05f
C9928 RST CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.258f
C9929 RST a_28663_n17626# 0.00464f
C9930 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 a_48017_9057# 1.43e-19
C9931 CLK a_22295_5018# 0.00134f
C9932 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT 0.0121f
C9933 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT 0.00154f
C9934 CLK_div_96_mag_0.JK_FF_mag_5.Q CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 1.48e-20
C9935 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 6.01e-19
C9936 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.359f
C9937 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_51397_6284# 7.4e-19
C9938 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C9939 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN 6.88e-21
C9940 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_28386_n743# 1.17e-20
C9941 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.415f
C9942 VDD110 a_44977_n18696# 3.14e-19
C9943 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT a_48741_9057# 0.0203f
C9944 RST CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 0.015f
C9945 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.0286f
C9946 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0715f
C9947 RST a_27856_n8779# 0.00185f
C9948 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 CLK_div_96_mag_0.JK_FF_mag_3.Q 2.25e-19
C9949 CLK_div_96_mag_0.JK_FF_mag_3.Q a_28737_n2996# 0.00789f
C9950 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_45927_6284# 0.00372f
C9951 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_31506_5018# 0.0731f
C9952 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT a_28463_n15537# 0.0203f
C9953 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_44061_n15627# 0.00392f
C9954 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 6.51e-19
C9955 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_23403_10099# 1.43e-19
C9956 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_45907_n16680# 0.0811f
C9957 VDD90 a_29623_6159# 3.14e-19
C9958 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 1.82e-19
C9959 VDD99 a_28823_n17626# 0.0132f
C9960 RST CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 0.0465f
C9961 CLK_div_96_mag_0.JK_FF_mag_0.Q a_23552_n1789# 1.63e-20
C9962 a_45081_n10160# a_45241_n10160# 0.0504f
C9963 CLK a_55132_5187# 5.03e-19
C9964 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 a_22551_n16006# 0.00347f
C9965 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT a_25482_n16632# 0.0731f
C9966 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_50721_n1102# 3.12e-19
C9967 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_23973_11196# 1.46e-19
C9968 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.VOUT 5.82e-21
C9969 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_36109_n8931# 0.00119f
C9970 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 7.24e-19
C9971 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 8.58e-20
C9972 CLK a_30060_9000# 0.0103f
C9973 CLK CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.00481f
C9974 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00335f
C9975 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.0285f
C9976 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 CLK_div_100_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00311f
C9977 VDD105 a_46867_7960# 3.14e-19
C9978 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0432f
C9979 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.122f
C9980 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_45251_n1102# 0.069f
C9981 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_26046_n16632# 0.00695f
C9982 CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 2.37f
C9983 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 0.338f
C9984 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 0.36f
C9985 F1 mux_8x1_ibr_0.mux_2x1_ibr_0.I1 0.011f
C9986 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K 0.0484f
C9987 CLK_div_108_new_mag_0.JK_FF_mag_1.Q CLK_div_108_new_mag_0.CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 0.00528f
C9988 CLK CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 6.19e-21
C9989 a_45787_574# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 8.17e-21
C9990 RST CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.146f
C9991 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.765f
C9992 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 a_50470_9057# 0.011f
C9993 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.065f
C9994 RST CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.0198f
C9995 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 a_47970_5143# 0.0101f
C9996 VDD93 a_23030_n8743# 3.14e-19
C9997 RST a_32175_n17626# 0.00498f
C9998 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 a_48832_n1102# 9.26e-19
C9999 RST CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.163f
C10000 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_42521_n13474# 0.00718f
C10001 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 a_36178_n16592# 0.069f
C10002 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_32076_6159# 3.25e-19
C10003 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 1.41e-20
C10004 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C10005 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_40818_n8887# 0.00372f
C10006 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN 0.0169f
C10007 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_25619_n7107# 0.0202f
C10008 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_50827_5143# 0.00695f
C10009 VDD108 a_46964_n9019# 3.14e-19
C10010 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_108_new_mag_0.JK_FF_mag_1.CLK 0.00199f
C10011 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 a_35184_880# 0.069f
C10012 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K a_51592_n16680# 5.58e-22
C10013 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_0.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.00392f
C10014 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 4.44e-20
C10015 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT 1.11e-20
C10016 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_29270_n743# 8.64e-19
C10017 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT 0.103f
C10018 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C10019 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0622f
C10020 CLK_div_108_new_mag_0.JK_FF_mag_1.Q CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.338f
C10021 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 8.16e-20
C10022 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.16f
C10023 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 2.59e-19
C10024 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.768f
C10025 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.0894f
C10026 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_48056_n5176# 0.0036f
C10027 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN 2.86e-19
C10028 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 2.97e-20
C10029 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK a_44247_n17599# 0.00117f
C10030 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_0.OUT 0.267f
C10031 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C10032 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.395f
C10033 CLK a_51438_n15583# 9.24e-19
C10034 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.338f
C10035 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 7.08e-20
C10036 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 a_41124_n16098# 4.44e-20
C10037 RST a_45235_n9063# 0.00211f
C10038 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 a_48092_n9063# 3.49e-20
C10039 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT 0.305f
C10040 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.321f
C10041 CLK_div_105_mag_0.CLK_div_10_mag_1.CLK CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.42f
C10042 VDD a_37999_n1822# 0.00444f
C10043 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 0.0529f
C10044 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.IN2 0.00216f
C10045 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00118f
C10046 RST a_24901_n6010# 8.06e-19
C10047 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_33019_n16588# 0.00964f
C10048 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.0758f
C10049 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 8.02e-20
C10050 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_32225_10099# 4.52e-20
C10051 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB 7.08e-20
C10052 RST CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT 0.0042f
C10053 CLK CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.315f
C10054 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 0.0609f
C10055 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.122f
C10056 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 9.52e-19
C10057 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C10058 VDD100 a_43671_7266# 0.00556f
C10059 RST a_48620_n5176# 5.85e-19
C10060 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_37801_n8887# 0.00372f
C10061 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.02f
C10062 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.0881f
C10063 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_50304_n16724# 1.5e-20
C10064 RST CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_2.OUT 0.0876f
C10065 a_29801_1733# CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.4e-19
C10066 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT a_33652_n13270# 0.0105f
C10067 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_52923_9057# 0.00118f
C10068 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_25508_n8734# 0.0202f
C10069 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_45131_n17599# 8.64e-19
C10070 CLK CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 1.05e-20
C10071 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT a_25328_n15535# 0.0203f
C10072 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.0622f
C10073 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00183f
C10074 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.175f
C10075 CLK_div_96_mag_0.JK_FF_mag_5.Q CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_0.OUT 8.73e-19
C10076 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 1.36e-19
C10077 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 5.36e-20
C10078 RST CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.136f
C10079 CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 a_40375_n7552# 0.0134f
C10080 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.0521f
C10081 a_43826_n7684# CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 1.4e-19
C10082 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB a_48629_1671# 1.86e-20
C10083 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 0.00392f
C10084 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.322f
C10085 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 Vdiv100 0.00396f
C10086 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 5.36e-20
C10087 RST a_44475_n5176# 0.00189f
C10088 a_39420_6265# a_39580_6265# 0.0504f
C10089 VDD108 a_53819_n5721# 3.14e-19
C10090 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.263f
C10091 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 a_44953_5143# 0.0101f
C10092 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_45241_n10160# 0.0202f
C10093 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_33180_n17626# 0.00372f
C10094 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 a_54022_n17599# 0.0102f
C10095 dec3x8_ibr_mag_0.and_3_ibr_2.nand3_mag_ibr_0.OUT a_39420_6821# 6.08e-20
C10096 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 5.36e-20
C10097 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 a_25508_n8734# 6.43e-21
C10098 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 1f
C10099 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 0.0599f
C10100 VDD90 a_33513_10099# 5.99e-19
C10101 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 a_31737_n15535# 2.79e-20
C10102 VDD100 a_49997_n1146# 0.00746f
C10103 RST CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_2.OUT 0.0544f
C10104 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 0.321f
C10105 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00122f
C10106 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 2.85e-20
C10107 VDD a_37999_880# 0.00444f
C10108 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.0622f
C10109 CLK_div_105_mag_0.CLK_div_10_mag_1.CLK CLK_div_105_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 2.16e-19
C10110 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT 3.2e-19
C10111 VDD99 a_35026_n18723# 2.65e-19
C10112 VDD108 a_43793_n10116# 3.14e-19
C10113 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_47430_n18696# 0.00392f
C10114 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 0.412f
C10115 RST a_28489_5018# 0.00186f
C10116 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_52139_n18696# 0.069f
C10117 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 a_50151_n2243# 0.00789f
C10118 RST a_53095_n5765# 0.00147f
C10119 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_2.OUT a_26256_3016# 9.1e-19
C10120 VDD110 a_51438_n15583# 3.14e-19
C10121 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 0.122f
C10122 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 5.7e-19
C10123 VDD110 a_52156_n16680# 3.14e-19
C10124 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT 0.343f
C10125 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.129f
C10126 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 0.00525f
C10127 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 a_29213_5018# 0.0101f
C10128 F0 a_39420_6265# 0.00181f
C10129 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT 0.0334f
C10130 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.266f
C10131 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.198f
C10132 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT 0.0854f
C10133 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 0.765f
C10134 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_5.QB 0.28f
C10135 RST a_40972_n9984# 1.17e-19
C10136 RST a_26663_398# 7.14e-19
C10137 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 3.27e-20
C10138 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_25619_n7107# 0.0697f
C10139 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_47970_5143# 0.00696f
C10140 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.391f
C10141 a_54022_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.00695f
C10142 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_54746_n17599# 0.00378f
C10143 CLK a_26343_n7107# 0.0118f
C10144 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.0063f
C10145 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0106f
C10146 RST CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 0.00589f
C10147 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00213f
C10148 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 a_50874_n15583# 0.0697f
C10149 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_33353_10099# 0.0732f
C10150 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 a_50358_1671# 0.069f
C10151 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB a_51486_1671# 1.41e-20
C10152 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 a_47905_1671# 0.0697f
C10153 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB a_50316_10154# 0.00964f
C10154 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN a_31177_7256# 5.1e-20
C10155 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_46259_n17599# 0.0157f
C10156 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 8.2e-19
C10157 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.346f
C10158 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB 1.96f
C10159 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 0.0172f
C10160 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_29777_5062# 0.0036f
C10161 CLK_div_108_new_mag_0.JK_FF_mag_1.QB CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 2.72e-19
C10162 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.765f
C10163 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 0.19f
C10164 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.23f
C10165 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.14f
C10166 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 1.31f
C10167 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.66f
C10168 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 8.16e-20
C10169 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 a_30469_n16590# 0.0157f
C10170 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.768f
C10171 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK 0.00254f
C10172 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 0.00846f
C10173 a_47863_10154# a_48023_10154# 0.0504f
C10174 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 a_35747_880# 0.069f
C10175 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C10176 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_24922_n17626# 0.0733f
C10177 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 8.98e-19
C10178 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB a_54498_n9064# 0.00392f
C10179 a_22559_n7106# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 5e-20
C10180 VDD105 a_46735_10154# 0.00152f
C10181 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 a_31128_n7028# 4.35e-19
C10182 a_26093_n743# a_26253_n743# 0.0504f
C10183 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 0.0108f
C10184 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 7.07e-20
C10185 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_51165_n17599# 2.88e-20
C10186 CLK_div_96_mag_0.JK_FF_mag_3.QB a_29461_n2996# 0.00696f
C10187 F0 m1_42708_4265# 4.37e-19
C10188 RST a_28099_n17626# 0.00311f
C10189 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 a_47453_9057# 0.011f
C10190 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 0.177f
C10191 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K a_34730_n16636# 8.64e-19
C10192 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_41284_n14596# 6.63e-20
C10193 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 7.14e-19
C10194 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 0.338f
C10195 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 9.62e-20
C10196 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0281f
C10197 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0209f
C10198 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0187f
C10199 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 5.53e-19
C10200 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_50833_6284# 3.12e-19
C10201 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 2.81e-20
C10202 RST a_31128_n7028# 9.29e-19
C10203 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT a_48581_9057# 0.0732f
C10204 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 0.0568f
C10205 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT 4.42e-19
C10206 a_46259_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.0811f
C10207 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.298f
C10208 a_23123_n7106# a_23283_n7106# 0.0504f
C10209 CLK_div_96_mag_0.JK_FF_mag_3.Q a_28577_n2996# 0.00335f
C10210 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.0378f
C10211 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_45363_6284# 0.069f
C10212 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_31346_5018# 0.0202f
C10213 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 0.108f
C10214 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00764f
C10215 Vdiv93 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.VOUT 0.0808f
C10216 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.346f
C10217 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT a_52839_n5# 0.00138f
C10218 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 0.415f
C10219 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_22839_10099# 0.011f
C10220 CLK CLK_div_96_mag_0.JK_FF_mag_4.Q 0.169f
C10221 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_45343_n16680# 0.00964f
C10222 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_52811_1671# 4.52e-20
C10223 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.0894f
C10224 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C10225 VDD a_38294_6265# 2.21e-19
C10226 VDD90 a_29059_6159# 3.14e-19
C10227 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.416f
C10228 VDD99 a_28663_n17626# 0.00888f
C10229 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.122f
C10230 CLK a_54568_5187# 4.86e-19
C10231 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.399f
C10232 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 1.77e-19
C10233 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_50157_n1146# 9.32e-19
C10234 RST CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 0.0455f
C10235 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT a_25322_n16632# 0.0202f
C10236 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.08f
C10237 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT 0.0238f
C10238 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 0.118f
C10239 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.0495f
C10240 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 4.66e-21
C10241 RST CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.156f
C10242 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_44413_n18696# 2.79e-20
C10243 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_54509_2768# 1.46e-19
C10244 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C10245 RST CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.179f
C10246 CLK_div_96_mag_0.JK_FF_mag_4.QB a_26814_1919# 0.00392f
C10247 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_32076_6159# 0.00378f
C10248 CLK_div_96_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 3.67e-20
C10249 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.00116f
C10250 VDD105 a_43831_7266# 0.234f
C10251 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 0.0635f
C10252 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 0.0598f
C10253 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN 8.03e-20
C10254 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN 0.11f
C10255 CLK CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 0.362f
C10256 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.338f
C10257 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.00243f
C10258 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 4.08e-20
C10259 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.0914f
C10260 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 a_33812_n13270# 0.0504f
C10261 CLK_div_93_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 3.34e-19
C10262 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00169f
C10263 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0175f
C10264 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_44475_n5176# 8.64e-19
C10265 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 a_49906_9057# 0.00118f
C10266 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 0.399f
C10267 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_55101_n6818# 0.00372f
C10268 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 a_47810_5143# 0.0102f
C10269 RST a_27150_11196# 0.00446f
C10270 RST a_32015_n17626# 0.00495f
C10271 VDD93 a_22466_n8743# 3.14e-19
C10272 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 7.24e-19
C10273 VDD100 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 0.0305f
C10274 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 7.24e-19
C10275 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_31512_6115# 0.00486f
C10276 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.362f
C10277 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN 0.00253f
C10278 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_40254_n8887# 0.069f
C10279 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 3.04f
C10280 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 3.25e-20
C10281 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.0683f
C10282 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_25055_n7107# 4.52e-20
C10283 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.0151f
C10284 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 1.83e-19
C10285 VDD108 a_46400_n9019# 3.56e-19
C10286 a_43383_n9019# CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 4.52e-20
C10287 a_48620_n5176# CLK_div_108_new_mag_0.JK_FF_mag_1.CLK 4.77e-20
C10288 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 4.25e-20
C10289 CLK_div_96_mag_0.JK_FF_mag_2.Q a_28737_n2996# 0.00212f
C10290 CLK CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.00673f
C10291 VDD Vdiv110 0.649f
C10292 a_55179_7683# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 3.02e-19
C10293 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 3.32e-20
C10294 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT 0.75f
C10295 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.00586f
C10296 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.122f
C10297 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.00518f
C10298 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 6.22e-20
C10299 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.647f
C10300 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0622f
C10301 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN a_45899_7960# 0.069f
C10302 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 3.81e-19
C10303 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_26253_n743# 2.88e-20
C10304 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 7.55e-19
C10305 Vdiv100 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT 6.29e-20
C10306 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 2.66f
C10307 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_0.Q 0.0171f
C10308 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_44413_n18696# 0.00392f
C10309 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 1.28e-20
C10310 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 1.16f
C10311 CLK a_50874_n15583# 3.8e-19
C10312 VDD99 a_32175_n17626# 0.00743f
C10313 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.268f
C10314 VDD a_39124_280# 0.00444f
C10315 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_41284_n14596# 0.0177f
C10316 RST a_45075_n9063# 0.00152f
C10317 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 Vdiv108 0.00531f
C10318 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 0.00212f
C10319 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 0.177f
C10320 VDD a_37436_n1822# 3.14e-19
C10321 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00183f
C10322 RST a_24337_n6010# 8.24e-19
C10323 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.00118f
C10324 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C10325 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.768f
C10326 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_32455_n16632# 0.00696f
C10327 VDD99 a_37328_6821# 0.00116f
C10328 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.00182f
C10329 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00126f
C10330 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 CLK_div_100_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 0.00442f
C10331 RST a_48056_n5176# 5.66e-19
C10332 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_37237_n8887# 0.069f
C10333 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1f
C10334 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0334f
C10335 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_50144_n16724# 1.17e-20
C10336 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.289f
C10337 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 4.11e-19
C10338 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT a_30915_n13291# 6.43e-19
C10339 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.175f
C10340 RST a_33898_n18723# 3.62e-19
C10341 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.399f
C10342 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_51193_n19793# 2.36e-22
C10343 CLK CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 3.76e-19
C10344 RST CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.0573f
C10345 a_48092_n9063# a_48252_n9063# 0.0504f
C10346 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.132f
C10347 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 4.66e-21
C10348 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_47140_n1146# 1.41e-20
C10349 a_22258_n2930# a_22418_n2930# 0.0504f
C10350 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 4.66e-21
C10351 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_51193_n19793# 0.00929f
C10352 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB a_48469_1671# 1.41e-20
C10353 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT 1.61e-19
C10354 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 7.47e-19
C10355 VDD dec3x8_ibr_mag_0.and_3_ibr_1.nand3_mag_ibr_0.OUT 0.72f
C10356 RST a_44315_n5176# 0.0014f
C10357 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB 2.59e-21
C10358 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 a_27375_n17626# 2.34e-20
C10359 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT 0.00123f
C10360 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 a_44793_5143# 0.0102f
C10361 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 a_53458_n17599# 0.00789f
C10362 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_45081_n10160# 0.0731f
C10363 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 a_24944_n8778# 0.00939f
C10364 dec3x8_ibr_mag_0.and_3_ibr_2.nand3_mag_ibr_0.OUT a_38454_6821# 0.0779f
C10365 VDD90 a_33353_10099# 2.65e-19
C10366 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 6.18e-19
C10367 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.913f
C10368 CLK_div_96_mag_0.JK_FF_mag_2.QB CLK_div_96_mag_0.JK_FF_mag_3.QB 2.36e-21
C10369 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 4.44e-20
C10370 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_2.Q 0.0343f
C10371 VDD99 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_2.OUT 0.0115f
C10372 VDD100 a_48832_n1102# 3.56e-19
C10373 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT m3_20882_n11188# 0.00257f
C10374 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 1.29f
C10375 VDD a_37436_880# 3.14e-19
C10376 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_51575_n18696# 0.0059f
C10377 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 7.03e-21
C10378 Vdiv96 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.OUT 0.00113f
C10379 VDD99 a_34462_n18723# 3.14e-19
C10380 VDD108 a_43229_n10116# 3.14e-19
C10381 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_30025_n2952# 0.00378f
C10382 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 8.16e-20
C10383 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 0.321f
C10384 VDD108 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 0.00127f
C10385 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 2.96e-19
C10386 RST a_28329_5018# 0.00186f
C10387 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 3.17e-19
C10388 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 a_49991_n2243# 0.00335f
C10389 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.00166f
C10390 RST a_51803_n5724# 9.71e-19
C10391 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_2.OUT a_26096_3016# 2.88e-20
C10392 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 0.065f
C10393 VDD110 a_50874_n15583# 3.14e-19
C10394 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.053f
C10395 VDD96 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.765f
C10396 VDD110 a_51592_n16680# 3.14e-19
C10397 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 a_29053_5018# 0.0102f
C10398 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 0.647f
C10399 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C10400 a_50715_n2243# a_50875_n2243# 0.0504f
C10401 CLK F1 0.31f
C10402 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.198f
C10403 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0352f
C10404 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.122f
C10405 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 1f
C10406 CLK_div_105_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00182f
C10407 Vdiv90 a_35184_880# 2.63e-21
C10408 a_44413_n18696# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0732f
C10409 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.00137f
C10410 CLK_div_96_mag_0.JK_FF_mag_5.QB CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_1.IN2 0.0592f
C10411 CLK_div_96_mag_0.JK_FF_mag_3.QB CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.198f
C10412 CLK_div_100_mag_0.CLK_div_10_mag_1.CLK CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB 0.307f
C10413 VDD110 a_39580_6821# 0.00156f
C10414 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 8.26e-20
C10415 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_25055_n7107# 0.0059f
C10416 Vdiv Vdiv108 0.00685f
C10417 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00183f
C10418 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_47810_5143# 0.00695f
C10419 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 a_26042_6159# 6.43e-21
C10420 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 5.49e-19
C10421 CLK a_26183_n7107# 0.0106f
C10422 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 3.09e-19
C10423 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_35186_n18723# 0.0203f
C10424 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.0654f
C10425 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.OUT 0.25f
C10426 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB a_33353_10099# 0.00392f
C10427 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K a_31571_n16632# 8.64e-19
C10428 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_45517_5187# 0.0036f
C10429 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_32789_10099# 0.00378f
C10430 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 a_49794_1671# 0.00372f
C10431 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 a_51028_n16724# 8.64e-19
C10432 VDD108 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.748f
C10433 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_49488_n13383# 0.015f
C10434 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_54051_9057# 0.0202f
C10435 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 a_47341_1671# 0.0059f
C10436 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.121f
C10437 VDD99 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.79e-19
C10438 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB a_49752_10154# 0.0811f
C10439 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 3.43e-19
C10440 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.104f
C10441 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C10442 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_43597_n6273# 8.64e-19
C10443 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 a_45695_n17599# 0.00859f
C10444 VDD96 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.397f
C10445 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.305f
C10446 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 1.31e-20
C10447 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.321f
C10448 RST a_45618_2768# 0.00186f
C10449 CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 m3_20882_n11188# 0.0251f
C10450 CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN a_49789_n9020# 4.94e-20
C10451 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 4.3e-20
C10452 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0345f
C10453 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT 0.0854f
C10454 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 1.17e-19
C10455 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 a_49794_1671# 4.52e-20
C10456 CLK_div_93_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.00384f
C10457 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 a_29905_n16590# 0.00859f
C10458 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00381f
C10459 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 3.6e-21
C10460 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00183f
C10461 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00157f
C10462 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0263f
C10463 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 8.16e-20
C10464 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB 0.198f
C10465 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 2.35e-20
C10466 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.0343f
C10467 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 a_47751_2768# 8.64e-19
C10468 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 a_51598_9057# 2.79e-20
C10469 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.109f
C10470 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 6.02e-20
C10471 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0343f
C10472 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 a_53464_n18696# 2.79e-20
C10473 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 2.48f
C10474 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_24358_n17626# 0.00378f
C10475 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT m3_20882_n11188# 0.00166f
C10476 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB a_53934_n9020# 3.33e-19
C10477 VDD mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT 0.648f
C10478 RST CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN 0.0388f
C10479 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 1.38e-19
C10480 RST CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00437f
C10481 VDD110 F1 0.111f
C10482 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB 0.25f
C10483 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C10484 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C10485 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.529f
C10486 VDD mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT 0.663f
C10487 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.2f
C10488 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.13f
C10489 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 1.54e-19
C10490 CLK_div_96_mag_0.JK_FF_mag_3.QB a_29301_n2996# 0.00695f
C10491 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_51005_n17599# 9.1e-19
C10492 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.CLK 1.71e-21
C10493 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 2.61f
C10494 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 0.395f
C10495 Vdiv90 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 0.00483f
C10496 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.16f
C10497 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 6.36e-19
C10498 RST a_27939_n17626# 0.00359f
C10499 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 a_46889_9057# 0.00118f
C10500 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_41124_n14596# 4.15e-19
C10501 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_44734_2768# 8.64e-19
C10502 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0622f
C10503 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_50269_6240# 9.32e-19
C10504 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT a_48017_9057# 0.00378f
C10505 VDD108 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 2.07e-19
C10506 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 1.51e-19
C10507 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.283f
C10508 a_45695_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.00964f
C10509 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT a_28580_n8735# 0.00378f
C10510 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 0.427f
C10511 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_52002_n15583# 0.00118f
C10512 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 a_48629_1671# 0.0101f
C10513 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_53464_n18696# 0.00486f
C10514 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.23f
C10515 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.765f
C10516 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 a_31129_n6271# 4.35e-19
C10517 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT 4.42e-19
C10518 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT a_55067_297# 0.00894f
C10519 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_22275_10099# 0.00118f
C10520 VDD99 a_25364_n19822# 5.92e-19
C10521 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_44779_n16724# 0.00696f
C10522 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_36024_n15495# 4.52e-20
C10523 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 1.49e-21
C10524 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.209f
C10525 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 6.23e-19
C10526 VDD99 a_28099_n17626# 0.0012f
C10527 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0622f
C10528 CLK_div_96_mag_0.JK_FF_mag_0.Q a_22424_n1833# 2.79e-20
C10529 VDD90 a_28495_6115# 2.66e-19
C10530 VDD100 a_51646_1671# 3.78e-19
C10531 CLK a_54004_5143# 4.68e-19
C10532 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_49997_n1146# 0.00111f
C10533 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0881f
C10534 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 8.36e-19
C10535 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 a_32750_n7675# 8.64e-19
C10536 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 0.652f
C10537 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.654f
C10538 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.338f
C10539 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT a_29298_n9832# 0.00378f
C10540 CLK_div_96_mag_0.JK_FF_mag_4.QB a_26250_1919# 3.08e-19
C10541 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_54051_9057# 0.0697f
C10542 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C10543 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_29307_n1855# 1.76e-20
C10544 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_31512_6115# 0.0732f
C10545 VDD99 dec3x8_ibr_mag_0.and_3_ibr_0.nand3_mag_ibr_0.OUT 8.06e-20
C10546 VDD105 a_43671_7266# 0.0407f
C10547 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN 0.00138f
C10548 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_0.OUT 0.0622f
C10549 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 a_48635_2768# 0.00119f
C10550 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 9.55e-20
C10551 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN a_29708_n8735# 6.6e-20
C10552 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.00739f
C10553 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 0.0134f
C10554 CLK CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 2.28f
C10555 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT a_48635_2768# 0.0202f
C10556 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 0.0314f
C10557 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 a_33652_n13270# 0.0186f
C10558 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.305f
C10559 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.00101f
C10560 CLK_div_93_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_40375_n7552# 3.25e-19
C10561 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.103f
C10562 CLK_div_108_new_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 2.34e-19
C10563 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.338f
C10564 a_33583_n16588# CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 2.58e-20
C10565 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.00165f
C10566 CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0345f
C10567 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_26760_5062# 0.0036f
C10568 RST a_26990_11196# 0.00446f
C10569 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 a_47246_5143# 0.00789f
C10570 VDD105 a_54775_9057# 0.00752f
C10571 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_54537_n6818# 0.069f
C10572 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.653f
C10573 RST a_31451_n17626# 0.00343f
C10574 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.107f
C10575 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.00183f
C10576 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 4.27e-20
C10577 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 a_47704_n1102# 6.43e-21
C10578 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K a_43901_n15627# 0.00472f
C10579 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 0.0765f
C10580 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_31352_6115# 0.00111f
C10581 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.0635f
C10582 RST a_55310_n17599# 2.58e-19
C10583 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.0107f
C10584 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.0859f
C10585 a_48056_n5176# CLK_div_108_new_mag_0.JK_FF_mag_1.CLK 1.73e-20
C10586 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_45618_2768# 0.0202f
C10587 VDD108 a_45235_n9063# 2.21e-19
C10588 CLK_div_96_mag_0.JK_FF_mag_2.Q a_28577_n2996# 0.00179f
C10589 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.122f
C10590 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 1.36e-19
C10591 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00157f
C10592 RST CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN 0.0185f
C10593 a_55019_7683# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 9.21e-20
C10594 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_26932_n2952# 0.0036f
C10595 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 0.00488f
C10596 CLK_div_100_mag_0.CLK_div_10_mag_1.CLK CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 0.256f
C10597 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.00447f
C10598 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 1.5e-20
C10599 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT 0.653f
C10600 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_26093_n743# 9.1e-19
C10601 VDD108 a_48620_n5176# 3.14e-19
C10602 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 8.16e-20
C10603 CLK a_50310_n15627# 0.0105f
C10604 VDD99 a_32015_n17626# 0.00305f
C10605 RST a_51165_n17599# 0.00211f
C10606 RST a_53487_9057# 6.14e-19
C10607 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 a_28268_n6266# 0.00353f
C10608 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.233f
C10609 CLK_div_108_new_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN a_43826_n7684# 3.25e-19
C10610 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_41124_n14596# 0.00765f
C10611 RST a_44511_n9019# 5.58e-19
C10612 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1f
C10613 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.468f
C10614 VDD a_36873_n1822# 0.00444f
C10615 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 3.98e-19
C10616 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_47252_6240# 1.41e-20
C10617 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 a_29059_6159# 1.25e-20
C10618 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00118f
C10619 Vdiv110 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K 0.0131f
C10620 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.00441f
C10621 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.046f
C10622 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_32295_n16632# 0.00695f
C10623 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_1.IN2 0.053f
C10624 VDD99 a_37168_6821# 0.00118f
C10625 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 a_33812_n13270# 2.84e-20
C10626 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K a_53126_6240# 8.64e-19
C10627 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_24133_11196# 1.17e-20
C10628 CLK_div_105_mag_0.CLK_div_10_mag_1.CLK CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 0.256f
C10629 Vdiv90 a_35747_n1222# 0.00298f
C10630 RST a_47704_n1102# 1.23e-20
C10631 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.103f
C10632 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT 0.298f
C10633 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0894f
C10634 VDD108 a_44475_n5176# 9.82e-19
C10635 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.0126f
C10636 CLK CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.298f
C10637 CLK_div_108_new_mag_0.JK_FF_mag_1.QB a_53255_n5765# 1.08e-20
C10638 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.998f
C10639 RST a_33334_n18723# 7.24e-19
C10640 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 0.657f
C10641 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0345f
C10642 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 2.63e-19
C10643 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 0.622f
C10644 Vdiv105 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT 3e-19
C10645 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.359f
C10646 RST a_30502_11196# 0.0049f
C10647 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 8.16e-20
C10648 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_46980_n1146# 1.86e-20
C10649 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 2.57f
C10650 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 0.797f
C10651 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 5.73e-19
C10652 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.013f
C10653 RST a_43751_n5176# 0.00127f
C10654 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT a_51034_9057# 0.0202f
C10655 VDD108 a_53095_n5765# 0.00514f
C10656 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 1.3f
C10657 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 a_44229_5143# 0.00789f
C10658 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 a_53298_n17599# 0.00335f
C10659 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_44517_n10160# 9.1e-19
C10660 dec3x8_ibr_mag_0.and_3_ibr_2.nand3_mag_ibr_0.OUT a_38294_6821# 0.0249f
C10661 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 a_24784_n8778# 0.0101f
C10662 VDD90 a_32789_10099# 3.14e-19
C10663 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN 0.00832f
C10664 VDD110 a_52293_n17599# 0.00152f
C10665 VDD100 a_48268_n1102# 3.14e-19
C10666 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.28f
C10667 VDD a_36873_880# 0.00444f
C10668 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_51011_n18696# 0.0697f
C10669 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 9.9e-19
C10670 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.103f
C10671 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_29461_n2996# 0.0733f
C10672 VDD99 a_33898_n18723# 3.14e-19
C10673 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 0.197f
C10674 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB a_26183_n7107# 0.00392f
C10675 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.321f
C10676 RST a_27324_5062# 9.66e-19
C10677 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 a_46777_1671# 4.52e-20
C10678 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 6.88e-21
C10679 a_54978_6284# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 4.52e-20
C10680 RST a_51239_n5724# 9.71e-19
C10681 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 5.08e-20
C10682 Vdiv110 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I1 0.0131f
C10683 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_29834_n699# 0.0036f
C10684 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN 0.112f
C10685 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1f
C10686 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0894f
C10687 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 a_28489_5018# 0.00789f
C10688 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_48620_n5176# 0.00372f
C10689 CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 Vdiv108 0.0668f
C10690 VDD110 a_48148_n17599# 0.00101f
C10691 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 a_23967_10099# 2.79e-20
C10692 VDD93 Vdiv105 0.632f
C10693 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0568f
C10694 a_44253_n18696# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0203f
C10695 RST a_39844_n10028# 0.00103f
C10696 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_10_mag_0.CLK 4.46e-19
C10697 VDD110 a_39420_6821# 0.00153f
C10698 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.122f
C10699 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 1.96f
C10700 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 a_24133_11196# 0.00335f
C10701 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_51439_n2199# 0.00378f
C10702 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 a_25478_6115# 0.00939f
C10703 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 8.16e-20
C10704 CLK a_25619_n7107# 3.01e-19
C10705 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 a_47187_2768# 0.069f
C10706 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.0794f
C10707 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 dec3x8_ibr_mag_0.and_3_ibr_6.nand3_mag_ibr_0.OUT 0.11f
C10708 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT 3.91e-20
C10709 RST CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT 0.0843f
C10710 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB 0.179f
C10711 Vdiv105 F0 2.84f
C10712 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 1.29e-19
C10713 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_35026_n18723# 0.0732f
C10714 CLK CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 2.61e-19
C10715 Vdiv99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 1.71e-21
C10716 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 0.122f
C10717 F2 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 0.136f
C10718 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB a_32789_10099# 3.33e-19
C10719 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.101f
C10720 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_48783_n13424# 5.19e-20
C10721 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 0.0693f
C10722 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.235f
C10723 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_53487_9057# 4.52e-20
C10724 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 1.53e-19
C10725 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_26072_n8734# 0.0059f
C10726 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 6.91e-20
C10727 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.28f
C10728 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.233f
C10729 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 0.424f
C10730 CLK_div_100_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 4.85e-20
C10731 CLK_div_108_new_mag_0.JK_FF_mag_1.Q CLK_div_108_new_mag_0.JK_FF_mag_0.QB 0.307f
C10732 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 0.0163f
C10733 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 a_47050_n7372# 0.01f
C10734 RST a_45458_2768# 0.00186f
C10735 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 0.321f
C10736 RST CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.142f
C10737 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00219f
C10738 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.338f
C10739 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C10740 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 a_29341_n16634# 0.0101f
C10741 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 a_39124_880# 0.00372f
C10742 CLK CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.0323f
C10743 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_29680_398# 4.52e-20
C10744 a_25420_n13385# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.132f
C10745 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.655f
C10746 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.343f
C10747 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C10748 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 6.22e-20
C10749 RST CLK_div_100_mag_0.CLK_div_10_mag_1.CLK 0.00173f
C10750 CLK CLK_div_100_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 3.06e-20
C10751 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT Vdiv110 0.0073f
C10752 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I1 a_37436_880# 0.00372f
C10753 F2 dec3x8_ibr_mag_0.and_3_ibr_0.nand3_mag_ibr_0.OUT 0.0275f
C10754 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00118f
C10755 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.231f
C10756 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 0.0264f
C10757 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 8.75e-19
C10758 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 4.49e-20
C10759 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 a_24116_n1789# 2.73e-19
C10760 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 a_28016_n8779# 2.79e-20
C10761 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_48558_n18696# 4.52e-20
C10762 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 a_50721_n1102# 1.25e-20
C10763 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 1.84e-19
C10764 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 9.87e-20
C10765 RST a_30589_n2952# 2.09e-19
C10766 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_50441_n17599# 0.0731f
C10767 RST a_50922_1671# 1.23e-20
C10768 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN a_52385_n13362# 2.31e-19
C10769 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT 0.00118f
C10770 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 2.77e-19
C10771 VDD100 a_45618_2768# 0.00727f
C10772 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 1.23f
C10773 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 2.48e-19
C10774 RST a_27375_n17626# 0.00439f
C10775 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_50109_6240# 0.00111f
C10776 RST CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.00223f
C10777 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 9.61e-21
C10778 CLK_div_96_mag_0.JK_FF_mag_0.QB CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 5.83e-19
C10779 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 0.0305f
C10780 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 5.87e-19
C10781 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT a_28016_n8779# 0.0732f
C10782 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.647f
C10783 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 0.111f
C10784 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 7.55e-19
C10785 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_51438_n15583# 0.011f
C10786 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 0.0592f
C10787 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 a_48469_1671# 0.00939f
C10788 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K 0.487f
C10789 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 8.16e-20
C10790 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_53304_n18696# 0.00111f
C10791 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 0.124f
C10792 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 a_30165_n6282# 0.0193f
C10793 dec3x8_ibr_mag_0.and_3_ibr_2.nand3_mag_ibr_0.OUT F0 0.0013f
C10794 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT a_54907_297# 0.0294f
C10795 VDD110 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.00721f
C10796 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.257f
C10797 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.0156f
C10798 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 a_44619_n16724# 0.00695f
C10799 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT a_35460_n15495# 0.0195f
C10800 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.VOUT CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN 0.00174f
C10801 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.0635f
C10802 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 0.00442f
C10803 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.00403f
C10804 VDD99 a_27939_n17626# 9.82e-19
C10805 VDD90 a_28335_6115# 0.00746f
C10806 VDD100 a_51486_1671# 2.66e-19
C10807 CLK a_53844_5143# 4.68e-19
C10808 CLK_div_108_new_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 1.35e-20
C10809 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_48832_n1102# 7.4e-19
C10810 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_22685_11196# 0.0036f
C10811 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_23123_n7106# 0.00119f
C10812 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.343f
C10813 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN 4.36e-20
C10814 VDD Vdiv99 0.387f
C10815 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.105f
C10816 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT a_28734_n9876# 0.0733f
C10817 CLK_div_96_mag_0.JK_FF_mag_4.QB a_25686_1919# 2.96e-19
C10818 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_53487_9057# 0.0059f
C10819 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT 8.94e-19
C10820 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_31352_6115# 0.0203f
C10821 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00178f
C10822 a_27170_6159# CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 4.52e-20
C10823 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 a_48475_2768# 0.00166f
C10824 Vdiv a_39124_880# 0.069f
C10825 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN a_29144_n8735# 2.72e-20
C10826 a_28657_n18723# a_28817_n18723# 0.0504f
C10827 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 1.96f
C10828 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT a_48475_2768# 0.0731f
C10829 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 m3_20882_n11188# 0.00101f
C10830 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 1.54e-21
C10831 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0854f
C10832 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 5.51e-20
C10833 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_25082_n17626# 0.00695f
C10834 RST Vdiv108 2.25f
C10835 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 0.198f
C10836 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT 0.259f
C10837 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_32009_n18723# 0.00119f
C10838 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 0.0432f
C10839 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT a_54978_6284# 1.54e-19
C10840 VDD105 a_54615_9057# 2.66e-19
C10841 RST a_26426_11196# 0.00311f
C10842 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 a_47086_5143# 0.00335f
C10843 RST a_31291_n17626# 0.00327f
C10844 VDD93 a_21742_n8787# 0.00533f
C10845 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00157f
C10846 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 5.07e-21
C10847 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 a_28817_n18723# 3.69e-19
C10848 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 a_47140_n1146# 0.00939f
C10849 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.CLK 9.71e-20
C10850 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 3.22e-20
C10851 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00118f
C10852 RST a_54746_n17599# 2.47e-19
C10853 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.471f
C10854 VDD90 CLK 3.08f
C10855 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0983f
C10856 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.768f
C10857 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT a_48017_9057# 0.0202f
C10858 RST CLK_div_105_mag_0.CLK_div_10_mag_1.CLK 0.00314f
C10859 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_45458_2768# 0.0731f
C10860 CLK_div_96_mag_0.JK_FF_mag_2.Q a_27496_n2952# 0.0157f
C10861 VDD99 Vdiv96 0.00674f
C10862 a_46867_7960# CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN 5.1e-20
C10863 VDD96 a_27227_398# 3.56e-19
C10864 CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 0.149f
C10865 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.122f
C10866 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_48741_9057# 0.00111f
C10867 CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 0.0445f
C10868 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_25529_n743# 0.0731f
C10869 VDD108 a_48056_n5176# 3.14e-19
C10870 VDD99 a_31451_n17626# 2.21e-19
C10871 CLK a_50150_n15627# 0.0114f
C10872 RST a_51005_n17599# 0.00198f
C10873 RST a_52923_9057# 6.14e-19
C10874 RST a_43947_n9019# 5.01e-19
C10875 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 1.14f
C10876 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0231f
C10877 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 1.08e-20
C10878 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_23403_10099# 0.0202f
C10879 VDD99 a_24391_n20290# 0.165f
C10880 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0948f
C10881 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 a_28495_6115# 0.00939f
C10882 VDD a_36310_n1822# 3.14e-19
C10883 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT a_53850_6284# 5.94e-20
C10884 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_47092_6240# 1.86e-20
C10885 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN a_45363_6284# 8.17e-21
C10886 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 a_30164_n7017# 7.37e-19
C10887 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 5.32e-19
C10888 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 a_33652_n13270# 9.09e-19
C10889 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_23973_11196# 1.5e-20
C10890 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN 0.00525f
C10891 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_55067_297# 0.00261f
C10892 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_46774_n6273# 0.00119f
C10893 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 2.37f
C10894 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_54669_2768# 1.17e-20
C10895 CLK CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 0.362f
C10896 VDD108 a_44315_n5176# 0.0012f
C10897 RST CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT 0.0284f
C10898 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.394f
C10899 Vdiv108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 1.26e-19
C10900 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 0.00236f
C10901 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN 4.17e-19
C10902 CLK_div_108_new_mag_0.JK_FF_mag_1.QB a_53095_n5765# 1.38e-20
C10903 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0175f
C10904 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0905f
C10905 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.198f
C10906 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 8.16e-20
C10907 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.995f
C10908 F0 mux_8x1_ibr_0.mux_2x1_ibr_0.I1 2.08e-19
C10909 RST a_30342_11196# 0.00487f
C10910 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 0.00274f
C10911 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_45815_n1102# 0.0114f
C10912 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_54775_9057# 0.0203f
C10913 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.999f
C10914 RST CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00498f
C10915 RST a_43591_n5176# 0.00127f
C10916 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.739f
C10917 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT a_50470_9057# 4.52e-20
C10918 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.231f
C10919 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT a_55357_n20487# 0.00894f
C10920 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 0.0116f
C10921 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00178f
C10922 VDD108 a_51803_n5724# 3.56e-19
C10923 a_26189_n6010# a_26349_n6010# 0.0504f
C10924 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.296f
C10925 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 a_44069_5143# 0.00335f
C10926 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_44357_n10160# 2.88e-20
C10927 a_45815_n1102# CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 4.52e-20
C10928 VDD mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.IN2 0.404f
C10929 VDD90 a_32225_10099# 3.14e-19
C10930 VDD110 a_51729_n17599# 0.00152f
C10931 VDD100 a_47704_n1102# 3.14e-19
C10932 VDD a_36310_880# 3.14e-19
C10933 VDD99 a_33334_n18723# 3.56e-19
C10934 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_29301_n2996# 0.0203f
C10935 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 0.98f
C10936 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB a_25619_n7107# 3.29e-19
C10937 RST a_26760_5062# 9.41e-19
C10938 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 0.299f
C10939 VDD96 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.662f
C10940 RST a_50675_n5724# 1.71e-19
C10941 VDD110 a_50150_n15627# 2.21e-19
C10942 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 2.59e-19
C10943 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_55132_5187# 0.00372f
C10944 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.122f
C10945 VDD110 a_50868_n16724# 2.21e-19
C10946 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C10947 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 0.233f
C10948 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 5.25e-20
C10949 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 a_28329_5018# 0.00335f
C10950 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.122f
C10951 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 5.08e-20
C10952 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_48056_n5176# 0.069f
C10953 VDD110 a_47988_n17599# 0.00123f
C10954 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.741f
C10955 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 8.71e-20
C10956 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 8.75e-20
C10957 CLK CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 7.92e-20
C10958 RST a_39684_n10028# 0.00119f
C10959 a_44253_n18696# a_44413_n18696# 0.0504f
C10960 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.00183f
C10961 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 5.98e-20
C10962 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_49276_n17599# 0.0157f
C10963 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_45541_n18696# 4.52e-20
C10964 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 8.16e-20
C10965 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 a_23973_11196# 0.00789f
C10966 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I1 0.328f
C10967 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 8.58e-20
C10968 CLK_div_105_mag_0.CLK_div_10_mag_1.CLK CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 6.64e-19
C10969 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_50875_n2243# 0.0733f
C10970 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 a_25318_6115# 0.0101f
C10971 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 a_46623_2768# 0.00372f
C10972 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 a_38454_6265# 0.00297f
C10973 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.321f
C10974 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_34462_n18723# 0.00378f
C10975 a_55019_7683# a_55179_7683# 0.186f
C10976 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT m3_20882_n11188# 0.00523f
C10977 VDD110 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.00665f
C10978 F2 a_37999_280# 2.16e-19
C10979 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0894f
C10980 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.121f
C10981 VDD99 a_33812_n13270# 0.0418f
C10982 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 0.265f
C10983 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_48623_n13424# 3.35e-20
C10984 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT m3_20882_n11188# 0.0024f
C10985 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_25508_n8734# 0.0697f
C10986 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 0.205f
C10987 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.343f
C10988 CLK_div_96_mag_0.JK_FF_mag_0.QB a_25650_n1899# 1.09e-20
C10989 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.0635f
C10990 RST a_44894_2768# 0.00169f
C10991 RST CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00543f
C10992 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.361f
C10993 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_28489_5018# 1.46e-19
C10994 CLK dec3x8_ibr_mag_0.and_3_ibr_7.nand3_mag_ibr_0.OUT 0.0017f
C10995 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 a_52003_n2199# 0.00372f
C10996 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.866f
C10997 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB 0.117f
C10998 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 a_38561_880# 0.069f
C10999 Vdiv110 Vdiv100 0.00673f
C11000 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 0.197f
C11001 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 0.0782f
C11002 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 a_29181_n16634# 0.0102f
C11003 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 0.00335f
C11004 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 8.39e-21
C11005 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.338f
C11006 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_29116_398# 0.0202f
C11007 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 0.0635f
C11008 VDD93 a_23289_n6009# 0.00108f
C11009 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 a_50470_9057# 6.06e-21
C11010 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB 0.913f
C11011 RST CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 9.76e-19
C11012 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.321f
C11013 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 1.03f
C11014 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 8.16e-20
C11015 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 7.16e-20
C11016 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.352f
C11017 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 0.00579f
C11018 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 3.39e-20
C11019 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I1 a_36873_880# 0.069f
C11020 F1 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 0.00219f
C11021 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB a_52806_n9020# 0.0112f
C11022 Vdiv105 m1_42708_4265# 0.00338f
C11023 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.994f
C11024 Vdiv100 a_39124_280# 4.15e-20
C11025 RST CLK_div_96_mag_0.JK_FF_mag_0.Q 0.152f
C11026 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_47994_n18696# 0.0202f
C11027 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN 0.00126f
C11028 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00163f
C11029 a_42529_n14305# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 3.01e-20
C11030 RST Vdiv93 0.264f
C11031 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 a_50157_n1146# 0.00939f
C11032 RST a_30025_n2952# 2e-19
C11033 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_54302_n1102# 4.52e-20
C11034 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_50281_n17599# 0.0202f
C11035 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.0188f
C11036 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.0631f
C11037 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN a_52225_n13362# 3.59e-19
C11038 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.399f
C11039 VDD100 a_45458_2768# 0.00299f
C11040 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 0.101f
C11041 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.177f
C11042 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB 0.0835f
C11043 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT 2.86e-19
C11044 RST a_26811_n17626# 0.00379f
C11045 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT 0.122f
C11046 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_28657_n18723# 0.00119f
C11047 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_48944_6284# 7.4e-19
C11048 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 3.54e-20
C11049 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 0.0646f
C11050 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 0.242f
C11051 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 0.338f
C11052 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 0.0766f
C11053 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_54746_n17599# 0.0036f
C11054 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0052f
C11055 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.CLK 1.47f
C11056 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 a_25686_1919# 0.069f
C11057 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT a_27856_n8779# 0.0203f
C11058 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN a_41117_n13911# 0.069f
C11059 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN a_23510_n15620# 1.14e-19
C11060 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_50874_n15583# 1.43e-19
C11061 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 6.11e-20
C11062 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 5.7e-20
C11063 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_52139_n18696# 7.4e-19
C11064 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 a_47905_1671# 1.25e-20
C11065 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 1.18f
C11066 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 5.98e-20
C11067 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_51592_n16680# 0.0036f
C11068 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.CLK 9.71e-20
C11069 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 a_29214_n6271# 0.0114f
C11070 VDD110 a_40375_n7552# 0.00131f
C11071 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_32071_11196# 0.069f
C11072 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB a_54615_9057# 0.00392f
C11073 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 0.0314f
C11074 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C11075 VDD96 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_2.OUT 0.752f
C11076 VDD110 dec3x8_ibr_mag_0.and_3_ibr_7.nand3_mag_ibr_0.OUT 0.182f
C11077 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.103f
C11078 VDD90 a_27170_6159# 3.56e-19
C11079 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_48422_n2199# 0.00378f
C11080 VDD99 a_27375_n17626# 0.00149f
C11081 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_29087_8532# 0.00168f
C11082 CLK a_53280_5143# 0.00111f
C11083 a_44357_n10160# a_44517_n10160# 0.0504f
C11084 VDD100 a_50922_1671# 3.14e-19
C11085 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_48268_n1102# 7.4e-19
C11086 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_22559_n7106# 1.43e-19
C11087 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 9.64e-19
C11088 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 4.27e-20
C11089 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 0.221f
C11090 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_53221_2768# 0.0036f
C11091 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 0.0016f
C11092 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT a_28574_n9876# 0.0203f
C11093 CLK_div_96_mag_0.JK_FF_mag_4.QB a_25122_1919# 0.0114f
C11094 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 3.23f
C11095 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.0435f
C11096 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.159f
C11097 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.398f
C11098 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.01f
C11099 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 a_47911_2768# 3.6e-22
C11100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.159f
C11101 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK 0.235f
C11102 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 6.3e-20
C11103 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 0.812f
C11104 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT a_47911_2768# 9.1e-19
C11105 a_28644_10099# CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 4.94e-20
C11106 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.00107f
C11107 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT m3_20882_n11188# 0.00189f
C11108 RST CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 0.158f
C11109 Vdiv110 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 2.4e-20
C11110 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_43757_n6273# 0.00119f
C11111 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K Vdiv105 4.19e-19
C11112 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_24922_n17626# 0.00696f
C11113 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.0725f
C11114 CLK CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.013f
C11115 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00335f
C11116 VDD96 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_2.OUT 0.751f
C11117 VDD100 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 1.05e-19
C11118 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 a_49122_n18696# 0.00372f
C11119 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_31445_n18723# 1.43e-19
C11120 VDD105 a_54051_9057# 3.14e-19
C11121 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 2.62e-20
C11122 RST a_26266_11196# 0.00359f
C11123 RST a_30727_n17626# 0.00382f
C11124 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 0.166f
C11125 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 a_46980_n1146# 0.0101f
C11126 RST CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 0.258f
C11127 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 0.652f
C11128 RST CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 0.133f
C11129 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.655f
C11130 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_26266_11196# 8.64e-19
C11131 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT a_47453_9057# 4.52e-20
C11132 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT 0.0758f
C11133 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.0948f
C11134 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_44894_2768# 9.1e-19
C11135 VDD108 a_44511_n9019# 3.14e-19
C11136 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 Vdiv110 0.00436f
C11137 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 6.35e-19
C11138 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.113f
C11139 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00103f
C11140 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 3.58e-19
C11141 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 0.11f
C11142 CLK_div_96_mag_0.JK_FF_mag_2.Q a_26932_n2952# 0.00859f
C11143 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 a_30915_n13291# 0.00476f
C11144 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_26663_398# 4.52e-20
C11145 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 5.37e-19
C11146 VDD96 a_26663_398# 3.14e-19
C11147 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 0.266f
C11148 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_48581_9057# 9.32e-19
C11149 VDD a_37999_n1222# 0.00444f
C11150 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_54947_n5721# 0.00118f
C11151 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_25369_n743# 0.0202f
C11152 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0156f
C11153 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.28f
C11154 VDD100 Vdiv108 0.529f
C11155 CLK a_48888_n15585# 9.33e-19
C11156 RST a_50441_n17599# 0.00247f
C11157 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00334f
C11158 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 m3_20882_n11188# 0.00142f
C11159 CLK a_50304_n16724# 0.00164f
C11160 CLK_div_96_mag_0.JK_FF_mag_2.Q CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.338f
C11161 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 8.16e-20
C11162 RST a_43383_n9019# 5.01e-19
C11163 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_22839_10099# 4.52e-20
C11164 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.417f
C11165 VDD a_35747_n1822# 0.00444f
C11166 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_54592_n18696# 4.52e-20
C11167 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_45927_6284# 0.0114f
C11168 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 a_28335_6115# 0.0101f
C11169 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.0622f
C11170 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 1.48e-20
C11171 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0854f
C11172 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C11173 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.00183f
C11174 CLK CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB 1.69e-20
C11175 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_23409_11196# 0.0203f
C11176 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00434f
C11177 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_54907_297# 0.00239f
C11178 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.995f
C11179 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 a_37328_6821# 0.00193f
C11180 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 a_48620_n5176# 0.0157f
C11181 RST CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00252f
C11182 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_54509_2768# 1.5e-20
C11183 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C11184 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C11185 VDD108 a_43751_n5176# 0.00888f
C11186 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.768f
C11187 CLK_div_108_new_mag_0.JK_FF_mag_1.Q CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 6.64e-19
C11188 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT Vdiv100 0.0153f
C11189 RST a_23510_n15620# 4.17e-19
C11190 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_29871_n1855# 1.63e-20
C11191 CLK_div_108_new_mag_0.JK_FF_mag_1.QB a_51803_n5724# 0.0114f
C11192 a_42521_n13474# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 0.132f
C11193 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT Vdiv100 0.0143f
C11194 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 9.55e-20
C11195 RST CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.0843f
C11196 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK a_50675_n5724# 6.43e-21
C11197 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 7.36e-21
C11198 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 7.89e-20
C11199 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_33019_n16588# 0.00378f
C11200 RST a_29778_11196# 0.00343f
C11201 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.768f
C11202 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.00481f
C11203 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_45251_n1102# 2.96e-19
C11204 Vdiv99 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 2.37e-20
C11205 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_54615_9057# 0.0732f
C11206 RST a_46774_n6273# 0.0012f
C11207 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0343f
C11208 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT a_55197_n20487# 0.0294f
C11209 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00183f
C11210 VDD108 a_51239_n5724# 3.14e-19
C11211 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.741f
C11212 VDD90 a_31661_10099# 3.56e-19
C11213 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 Vdiv110 0.00326f
C11214 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 0.0188f
C11215 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 0.411f
C11216 VDD100 a_47140_n1146# 2.66e-19
C11217 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_27150_11196# 0.0202f
C11218 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.16f
C11219 VDD a_35747_880# 0.00444f
C11220 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 0.00101f
C11221 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_28737_n2996# 1.5e-20
C11222 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB a_25055_n7107# 2.96e-19
C11223 RST a_26196_5018# 0.00186f
C11224 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00943f
C11225 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 0.0107f
C11226 RST a_50111_n5768# 4.58e-19
C11227 VDD110 a_48888_n15585# 3.56e-19
C11228 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_54568_5187# 0.069f
C11229 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 0.0294f
C11230 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 0.342f
C11231 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00115f
C11232 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT 0.802f
C11233 CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_99_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.124f
C11234 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 4.04e-19
C11235 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN 0.418f
C11236 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0886f
C11237 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C11238 RST CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 2.96e-19
C11239 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 a_23703_n287# 0.00119f
C11240 a_28392_354# a_28552_354# 0.0504f
C11241 VDD96 dec3x8_ibr_mag_0.and_3_ibr_0.nand3_mag_ibr_0.OUT 8.14e-19
C11242 VDD110 a_47424_n17599# 0.00863f
C11243 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 0.397f
C11244 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0555f
C11245 RST CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 0.133f
C11246 RST a_39120_n10028# 0.00218f
C11247 CLK CLK_div_108_new_mag_0.CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 0.0983f
C11248 CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K 0.00761f
C11249 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 a_48712_n17599# 0.00859f
C11250 CLK CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00433f
C11251 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.00452f
C11252 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_44977_n18696# 0.0202f
C11253 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_50715_n2243# 0.0203f
C11254 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 a_23409_11196# 0.0102f
C11255 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT 0.0758f
C11256 F1 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 4.51e-21
C11257 CLK CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT 9.25e-19
C11258 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 1.27f
C11259 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 2.13e-20
C11260 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 a_24153_6159# 0.069f
C11261 CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 7.06e-20
C11262 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.121f
C11263 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 a_38294_6265# 0.00699f
C11264 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K a_27334_n16588# 1.44e-21
C11265 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB a_31661_10099# 0.0112f
C11266 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB 7.08e-20
C11267 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_44229_5143# 1.46e-19
C11268 VDD99 a_33652_n13270# 0.235f
C11269 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 7.24e-19
C11270 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.0432f
C11271 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.01f
C11272 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K a_52951_7381# 0.0027f
C11273 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_41117_n13911# 0.00544f
C11274 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 0.0593f
C11275 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_51871_n5# 5.1e-20
C11276 RST CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB 0.696f
C11277 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN 1.15e-19
C11278 CLK_div_96_mag_0.JK_FF_mag_0.QB a_25490_n1899# 1.37e-20
C11279 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_37801_n8887# 0.0112f
C11280 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 0.0128f
C11281 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 mux_8x1_ibr_0.mux_2x1_ibr_0.I0 0.051f
C11282 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN 3.59e-20
C11283 CLK_div_96_mag_0.JK_FF_mag_2.Q CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.41f
C11284 RST a_44734_2768# 0.00128f
C11285 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 3.14e-20
C11286 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 9.8e-19
C11287 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 1.03e-19
C11288 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_54414_6284# 4.52e-20
C11289 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 a_51439_n2199# 0.069f
C11290 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB a_51598_9057# 0.00392f
C11291 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.103f
C11292 RST CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 3.05f
C11293 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 a_23283_n7106# 0.0101f
C11294 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 a_28617_n16634# 0.00789f
C11295 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 3.61e-21
C11296 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 a_49906_9057# 0.069f
C11297 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 0.994f
C11298 VDD93 CLK 3.63f
C11299 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 8.16e-20
C11300 RST CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT 0.0284f
C11301 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB a_51641_n9064# 1.86e-20
C11302 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 8.16e-20
C11303 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 0.00145f
C11304 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 3.38e-19
C11305 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 a_49997_n1146# 0.0101f
C11306 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.0576f
C11307 a_25369_n743# a_25529_n743# 0.0504f
C11308 RST CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.00355f
C11309 CLK F0 0.213f
C11310 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_53738_n1102# 0.0202f
C11311 RST a_29461_n2996# 0.00178f
C11312 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0576f
C11313 VDD100 a_44894_2768# 2.21e-19
C11314 a_48581_9057# a_48741_9057# 0.0504f
C11315 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00545f
C11316 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0894f
C11317 VDD99 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB 9.92e-19
C11318 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 1.03f
C11319 CLK_div_96_mag_0.JK_FF_mag_0.QB CLK_div_96_mag_0.JK_FF_mag_2.Q 7.83e-20
C11320 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_28093_n18723# 1.43e-19
C11321 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN 5.7e-20
C11322 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_48380_6284# 7.4e-19
C11323 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_53333_10154# 0.069f
C11324 VDD99 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 0.00264f
C11325 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 a_36873_280# 8.2e-19
C11326 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_33358_5062# 0.00372f
C11327 RST CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00936f
C11328 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 0.21f
C11329 CLK CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.00673f
C11330 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 a_23948_n13382# 0.00186f
C11331 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 a_25122_1919# 0.00372f
C11332 RST CLK_div_110_mag_0.CLK_div_10_mag_0.CLK 0.671f
C11333 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.398f
C11334 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 7.63e-19
C11335 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_50310_n15627# 0.00119f
C11336 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 0.385f
C11337 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_51575_n18696# 7.4e-19
C11338 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_51193_n19793# 3.38e-20
C11339 a_50109_6240# a_50269_6240# 0.0504f
C11340 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 a_27334_n16588# 0.00372f
C11341 Vdiv96 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT 8.22e-21
C11342 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 2.11e-19
C11343 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_31507_11196# 0.00372f
C11344 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.432f
C11345 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB a_54051_9057# 3.33e-19
C11346 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.00183f
C11347 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 1.49e-21
C11348 RST CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.0625f
C11349 F2 Vdiv108 0.0469f
C11350 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_26636_n8734# 0.00118f
C11351 VDD110 a_39580_6265# 0.00172f
C11352 VDD99 a_26811_n17626# 0.00149f
C11353 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 1.12e-19
C11354 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_47858_n2243# 0.0733f
C11355 VDD90 a_26606_6159# 3.14e-19
C11356 VDD100 a_50358_1671# 3.14e-19
C11357 CLK a_53120_5143# 0.00111f
C11358 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 3.66e-20
C11359 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 a_51647_n10161# 0.00335f
C11360 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_47704_n1102# 3.12e-19
C11361 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_21995_n7106# 0.011f
C11362 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 2.12e-19
C11363 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 a_42083_n15712# 0.0178f
C11364 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 1.9e-20
C11365 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.122f
C11366 VDD108 Vdiv108 1.63f
C11367 a_36873_880# Vdiv100 5.55e-19
C11368 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT a_28010_n9876# 1.5e-20
C11369 CLK m3_20882_n11188# 0.0033f
C11370 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.0152f
C11371 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 dec3x8_ibr_mag_0.and_3_ibr_1.nand3_mag_ibr_0.OUT 0.0808f
C11372 CLK CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 7.81e-19
C11373 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 0.129f
C11374 VDD93 VDD110 0.648f
C11375 a_55197_n20487# a_55357_n20487# 0.186f
C11376 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_51575_n18696# 4.52e-20
C11377 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00393f
C11378 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 2.81e-20
C11379 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 dec3x8_ibr_mag_0.and_3_ibr_0.nand3_mag_ibr_0.OUT 0.271f
C11380 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT 0.0622f
C11381 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0246f
C11382 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.768f
C11383 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00118f
C11384 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C11385 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 6.71e-19
C11386 CLK_div_96_mag_0.JK_FF_mag_5.QB CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 4.51e-20
C11387 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 2.62e-19
C11388 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0945f
C11389 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 2.37f
C11390 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT a_47751_2768# 2.88e-20
C11391 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.0161f
C11392 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 9.86e-19
C11393 a_54664_n10161# m3_20882_n11188# 0.00102f
C11394 RST CLK_div_90_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.00352f
C11395 CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 a_23691_9000# 7.48e-20
C11396 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00335f
C11397 VDD90 a_29087_8532# 0.165f
C11398 CLK_div_93_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 8.04e-19
C11399 a_32750_n7675# CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.132f
C11400 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_33358_5062# 0.0811f
C11401 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_27144_10099# 1.09e-20
C11402 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_24358_n17626# 0.00964f
C11403 VDD110 F0 1.12f
C11404 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 3.92e-19
C11405 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_25472_5018# 1.46e-19
C11406 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_30881_n18723# 0.011f
C11407 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 a_48558_n18696# 0.069f
C11408 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.106f
C11409 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C11410 RST a_25702_11196# 0.00439f
C11411 VDD105 a_53487_9057# 3.14e-19
C11412 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 5.08e-20
C11413 RST a_30163_n17626# 0.00373f
C11414 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.126f
C11415 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_49122_n18696# 0.00118f
C11416 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 a_45815_n1102# 0.069f
C11417 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 0.159f
C11418 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_25856_10099# 0.069f
C11419 a_25686_1919# CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 2.05e-20
C11420 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K 6.13e-20
C11421 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB 0.28f
C11422 Vdiv90 F1 0.00151f
C11423 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 0.00116f
C11424 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_44734_2768# 2.88e-20
C11425 VDD108 a_43947_n9019# 3.14e-19
C11426 a_48635_2768# Vdiv110 0.00138f
C11427 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.398f
C11428 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 0.122f
C11429 a_50232_n7685# CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K 0.00168f
C11430 CLK_div_96_mag_0.JK_FF_mag_2.Q a_26368_n2996# 0.0101f
C11431 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 5.05e-20
C11432 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 a_30210_n13332# 0.00107f
C11433 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_26099_398# 0.0202f
C11434 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C11435 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_23743_5062# 0.00378f
C11436 VDD96 a_26099_398# 3.14e-19
C11437 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 a_29214_n6271# 6.36e-20
C11438 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_25644_n2996# 1.46e-19
C11439 CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 5.32e-19
C11440 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.199f
C11441 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_48017_9057# 3.12e-19
C11442 VDD a_36873_n1222# 0.00444f
C11443 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.00157f
C11444 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_54383_n5721# 0.011f
C11445 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 0.0189f
C11446 CLK a_48324_n15585# 9.25e-19
C11447 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 a_52002_n15583# 0.00372f
C11448 VDD99 a_30727_n17626# 3.14e-19
C11449 RST a_50281_n17599# 0.00247f
C11450 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00545f
C11451 VDD99 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 0.0987f
C11452 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.0435f
C11453 CLK a_50144_n16724# 0.00117f
C11454 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.159f
C11455 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.378f
C11456 VDD a_35184_n1822# 3.14e-19
C11457 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_54028_n18696# 0.0202f
C11458 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 6.82e-19
C11459 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_45363_6284# 2.96e-19
C11460 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 a_27170_6159# 0.069f
C11461 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 a_36024_n15495# 0.00605f
C11462 VDD110 m3_20882_n11188# 0.732f
C11463 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.122f
C11464 CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0343f
C11465 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 a_26790_n9831# 0.0157f
C11466 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 4.08f
C11467 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_23249_11196# 0.0733f
C11468 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 a_37168_6821# 0.00175f
C11469 RST a_45815_n1102# 0.00104f
C11470 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT 0.768f
C11471 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 a_48056_n5176# 0.00859f
C11472 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_53945_2768# 0.0203f
C11473 VDD108 a_43591_n5176# 0.0132f
C11474 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.647f
C11475 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 1.04e-19
C11476 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 1.33e-20
C11477 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.251f
C11478 CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.338f
C11479 CLK_div_108_new_mag_0.JK_FF_mag_1.QB a_51239_n5724# 2.96e-19
C11480 RST CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN 9.43e-19
C11481 F1 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 0.0874f
C11482 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK a_53458_n17599# 0.0024f
C11483 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 8.16e-20
C11484 RST a_26790_n9831# 9.82e-19
C11485 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK a_50111_n5768# 0.00939f
C11486 RST CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0602f
C11487 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_32455_n16632# 0.0733f
C11488 RST a_29618_11196# 0.00327f
C11489 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 7.24e-19
C11490 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_35032_n17626# 1.46e-19
C11491 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_54182_n17599# 8.64e-19
C11492 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_44687_n1102# 3.33e-19
C11493 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_54051_9057# 0.00378f
C11494 RST a_46614_n6273# 0.00163f
C11495 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0432f
C11496 CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00393f
C11497 VDD108 a_50675_n5724# 3.14e-19
C11498 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 7.89e-19
C11499 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 1.03f
C11500 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00125f
C11501 RST CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN 0.0275f
C11502 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.349f
C11503 CLK_div_100_mag_0.CLK_div_10_mag_1.CLK CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 4.19e-19
C11504 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.768f
C11505 RST CLK_div_96_mag_0.JK_FF_mag_2.QB 0.257f
C11506 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.00163f
C11507 VDD100 a_46980_n1146# 3.78e-19
C11508 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 4.36e-20
C11509 VDD99 a_23510_n15620# 0.167f
C11510 Vdiv110 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 0.00873f
C11511 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 2.12e-19
C11512 CLK_div_96_mag_0.JK_FF_mag_3.Q a_30435_n1855# 0.0696f
C11513 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_26990_11196# 0.0731f
C11514 VDD a_35184_880# 3.14e-19
C11515 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 0.502f
C11516 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_28577_n2996# 1.17e-20
C11517 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB a_48581_9057# 0.00392f
C11518 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB a_24491_n7107# 0.0114f
C11519 a_47036_n15629# a_47196_n15629# 0.0504f
C11520 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.122f
C11521 RST a_26036_5018# 0.00169f
C11522 RST a_49951_n5768# 5.6e-19
C11523 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.11f
C11524 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.00183f
C11525 VDD110 a_48324_n15585# 3.14e-19
C11526 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_28546_n743# 1.46e-19
C11527 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00118f
C11528 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.0285f
C11529 VDD110 a_50144_n16724# 2.76e-19
C11530 CLK CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 0.00163f
C11531 CLK CLK_div_108_new_mag_0.JK_FF_mag_1.Q 0.014f
C11532 a_49991_n2243# a_50151_n2243# 0.0504f
C11533 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 a_23139_n287# 1.43e-19
C11534 VDD110 a_47264_n17599# 0.0123f
C11535 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 a_22275_10099# 0.069f
C11536 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT a_32175_n17626# 5.54e-20
C11537 VDD93 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 0.00125f
C11538 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 9.98e-19
C11539 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C11540 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 0.00127f
C11541 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00118f
C11542 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.768f
C11543 RST a_38960_n10028# 0.00218f
C11544 RST CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.00208f
C11545 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1f
C11546 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 a_23249_11196# 0.0101f
C11547 F1 dec3x8_ibr_mag_0.and_3_ibr_4.nand3_mag_ibr_0.OUT 0.0359f
C11548 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_50151_n2243# 1.5e-20
C11549 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_23967_10099# 0.00392f
C11550 a_33353_10099# a_33513_10099# 0.0504f
C11551 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 a_23589_6159# 6.06e-21
C11552 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 3.6e-19
C11553 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_34896_n15539# 1.19e-20
C11554 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C11555 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 1.2e-19
C11556 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT a_33812_n13270# 0.198f
C11557 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_53463_n16728# 4.28e-19
C11558 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K a_26770_n16588# 4.96e-22
C11559 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 0.0172f
C11560 RST CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00229f
C11561 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.235f
C11562 VDD99 a_30915_n13291# 3.14e-19
C11563 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 0.392f
C11564 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 0.149f
C11565 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 3.38e-19
C11566 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 1.99e-20
C11567 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB 0.915f
C11568 VDD99 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 7.57e-21
C11569 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_2.OUT CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT 0.121f
C11570 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_5.QB 0.0385f
C11571 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00392f
C11572 CLK_div_96_mag_0.JK_FF_mag_0.QB a_24116_n1789# 0.0114f
C11573 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 2.57e-19
C11574 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN 2.35e-19
C11575 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C11576 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K Vdiv90 2.52e-19
C11577 a_21742_n8787# a_21902_n8787# 0.0504f
C11578 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0934f
C11579 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK a_53464_n18696# 2.06e-19
C11580 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_3.Q 1.07e-19
C11581 VDD96 Vdiv96 0.503f
C11582 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.31f
C11583 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_53850_6284# 0.0202f
C11584 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB a_51034_9057# 3.25e-19
C11585 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 0.11f
C11586 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.273f
C11587 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_54568_5187# 0.00378f
C11588 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 0.00481f
C11589 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 a_28457_n16634# 0.00335f
C11590 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 a_23123_n7106# 0.00939f
C11591 VDD108 Vdiv93 0.0363f
C11592 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.272f
C11593 VDD93 a_22565_n6009# 2.21e-19
C11594 Vdiv96 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I1 0.00214f
C11595 RST CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00218f
C11596 VDD mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 0.405f
C11597 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 1.48e-20
C11598 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_31445_n18723# 0.0697f
C11599 Vdiv110 Vdiv 0.203f
C11600 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0135f
C11601 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0592f
C11602 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.OUT a_37999_n1822# 0.00949f
C11603 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 5.11e-19
C11604 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I1 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.11f
C11605 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB a_51481_n9064# 1.41e-20
C11606 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.133f
C11607 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT Vdiv90 0.12f
C11608 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.VOUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 1.53e-22
C11609 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K 0.00825f
C11610 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 a_22424_n1833# 3.23e-20
C11611 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.783f
C11612 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 a_48832_n1102# 0.069f
C11613 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00183f
C11614 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.654f
C11615 a_50232_n7685# CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 1.4e-19
C11616 RST a_29301_n2996# 0.00193f
C11617 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 5.05e-20
C11618 CLK_div_99_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN a_31733_n19822# 0.069f
C11619 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_24127_10099# 1.86e-20
C11620 RST CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN 0.0116f
C11621 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0345f
C11622 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 0.233f
C11623 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 0.00103f
C11624 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 9.24e-20
C11625 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_27529_n18723# 0.011f
C11626 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_47816_6284# 3.12e-19
C11627 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_51729_n17599# 5.02e-20
C11628 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.175f
C11629 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_52769_10154# 0.00372f
C11630 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_46105_n18696# 0.00118f
C11631 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I1 0.00146f
C11632 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_32794_5062# 0.069f
C11633 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.00395f
C11634 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_29751_n15493# 4.52e-20
C11635 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT 0.58f
C11636 RST CLK_div_96_mag_0.JK_FF_mag_4.QB 0.242f
C11637 CLK_div_90_mag_0.CLK_div_10_mag_0.CLK a_23025_6159# 6.43e-21
C11638 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 5.42e-20
C11639 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 5.2e-20
C11640 Vdiv108 CLK_div_108_new_mag_0.JK_FF_mag_1.QB 1.43e-19
C11641 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_51011_n18696# 3.12e-19
C11642 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 a_26770_n16588# 0.069f
C11643 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.414f
C11644 VDD93 a_29213_n7028# 3.14e-19
C11645 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB a_53487_9057# 2.96e-19
C11646 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 5.52e-20
C11647 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.192f
C11648 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_26072_n8734# 0.011f
C11649 CLK_div_108_new_mag_0.JK_FF_mag_0.QB CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.25f
C11650 VDD110 a_39420_6265# 0.00153f
C11651 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 0.00132f
C11652 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT Vdiv108 1.51e-19
C11653 VDD90 a_26042_6159# 3.14e-19
C11654 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_47698_n2243# 0.0203f
C11655 VDD100 a_49794_1671# 3.56e-19
C11656 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 a_26349_n6010# 0.0117f
C11657 CLK a_52115_5187# 5.03e-19
C11658 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 6.82e-19
C11659 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_47140_n1146# 9.32e-19
C11660 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 a_51487_n10161# 0.00789f
C11661 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_29461_n2996# 2.88e-20
C11662 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_21431_n7106# 0.00118f
C11663 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 0.149f
C11664 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.122f
C11665 a_36310_880# Vdiv100 4.07e-19
C11666 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.0789f
C11667 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT a_27850_n9876# 1.17e-20
C11668 VDD93 a_39402_n7788# 5.95e-19
C11669 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 0.122f
C11670 CLK m1_42708_4265# 0.206f
C11671 Vdiv96 mux_8x1_ibr_0.mux_2x1_ibr_0.I0 4.93e-19
C11672 RST CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0614f
C11673 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_51011_n18696# 0.0202f
C11674 Vdiv90 a_35747_280# 3.43e-19
C11675 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 9.14e-19
C11676 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 2.59e-21
C11677 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.CLK 1.47f
C11678 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT 0.053f
C11679 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_29680_398# 0.0059f
C11680 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.756f
C11681 mux_8x1_ibr_0.mux_2x1_ibr_0.I0 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.11f
C11682 dec3x8_ibr_mag_0.and_3_ibr_5.IN3 F1 0.384f
C11683 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 2.46e-20
C11684 a_50447_n18696# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.0732f
C11685 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0833f
C11686 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_1.IN2 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00352f
C11687 a_54504_n10161# m3_20882_n11188# 0.00102f
C11688 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 0.0106f
C11689 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 a_22544_n13819# 0.00572f
C11690 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 a_37801_n8887# 0.069f
C11691 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_32794_5062# 0.00964f
C11692 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_23794_n17626# 0.0811f
C11693 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_26984_10099# 8.77e-21
C11694 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB Vdiv110 0.0113f
C11695 a_43760_1671# CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 1.54e-19
C11696 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00213f
C11697 CLK_div_96_mag_0.JK_FF_mag_4.QB a_26256_3016# 0.00695f
C11698 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0635f
C11699 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.159f
C11700 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_30317_n18723# 0.00118f
C11701 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 1.19f
C11702 VDD105 a_52923_9057# 3.56e-19
C11703 RST a_25138_11196# 0.00379f
C11704 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_48558_n18696# 0.011f
C11705 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 4.69e-20
C11706 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 a_45251_n1102# 6.06e-21
C11707 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.25f
C11708 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 4.01e-20
C11709 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_25292_10099# 0.00372f
C11710 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 0.295f
C11711 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K a_43895_n16724# 8.64e-19
C11712 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT 0.00166f
C11713 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 3.81e-19
C11714 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 1.29f
C11715 mux_8x1_ibr_0.mux_2x1_ibr_0.I0 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 0.0449f
C11716 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.648f
C11717 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT a_52385_n13362# 8.64e-19
C11718 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.0172f
C11719 VDD108 a_43383_n9019# 3.56e-19
C11720 a_48475_2768# Vdiv110 0.00138f
C11721 Vdiv93 a_43597_n6273# 4.38e-19
C11722 VDD90 a_27144_10099# 5.99e-19
C11723 CLK_div_96_mag_0.JK_FF_mag_2.Q a_26208_n2996# 0.0102f
C11724 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 5.55e-21
C11725 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 a_30050_n13332# 0.00271f
C11726 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 2.6e-20
C11727 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_23179_5018# 0.0733f
C11728 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT 0.58f
C11729 VDD99 dec3x8_ibr_mag_0.and_3_ibr_6.nand3_mag_ibr_0.OUT 0.0321f
C11730 VDD96 a_25535_354# 2.65e-19
C11731 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_47453_9057# 7.4e-19
C11732 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_55310_n17599# 0.00372f
C11733 VDD a_35747_n1222# 0.00444f
C11734 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0622f
C11735 Vdiv99 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.VOUT 1.19f
C11736 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_53819_n5721# 1.43e-19
C11737 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN a_31129_n6271# 8.67e-20
C11738 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 a_35747_280# 1.5e-19
C11739 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 a_51438_n15583# 0.069f
C11740 CLK a_47760_n15585# 3.81e-19
C11741 VDD99 a_30163_n17626# 3.14e-19
C11742 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 9.69e-19
C11743 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 1.05e-19
C11744 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.118f
C11745 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.108f
C11746 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 a_26606_6159# 6.06e-21
C11747 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 a_35460_n15495# 0.0697f
C11748 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_44799_6284# 3.33e-19
C11749 VDD110 m1_42708_4265# 3.2e-19
C11750 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0309f
C11751 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 a_26226_n9831# 0.00859f
C11752 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_22685_11196# 0.00378f
C11753 CLK_div_108_new_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 7.3e-19
C11754 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_26616_n15491# 4.52e-20
C11755 RST a_45251_n1102# 0.00167f
C11756 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_53785_2768# 0.0733f
C11757 Vdiv105 mux_8x1_ibr_0.mux_2x1_ibr_0.I1 1.08e-19
C11758 CLK CLK_div_90_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.0983f
C11759 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 a_28734_n9876# 8.64e-19
C11760 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 0.995f
C11761 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 3.38e-19
C11762 CLK_div_96_mag_0.JK_FF_mag_3.QB CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.28f
C11763 CLK_div_108_new_mag_0.JK_FF_mag_1.QB a_50675_n5724# 3.33e-19
C11764 RST a_45787_574# 4.48e-19
C11765 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK a_53298_n17599# 0.0024f
C11766 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 0.0635f
C11767 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK a_49951_n5768# 0.0101f
C11768 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT Vdiv 0.346f
C11769 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 1.41e-20
C11770 RST a_26226_n9831# 9.62e-19
C11771 a_29087_8532# CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 5.89e-19
C11772 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 1.97f
C11773 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT m3_20882_n11188# 0.00166f
C11774 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_32295_n16632# 0.0203f
C11775 RST a_29054_11196# 0.00382f
C11776 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 9.72f
C11777 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_44123_n1146# 0.00392f
C11778 CLK CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 0.0256f
C11779 RST a_45449_n6273# 0.00208f
C11780 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.487f
C11781 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 0.162f
C11782 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 2.59e-21
C11783 a_23123_n7106# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 3.87e-20
C11784 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.0894f
C11785 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_28644_10099# 4.52e-20
C11786 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 0.0286f
C11787 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00118f
C11788 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_30915_n13291# 3.04e-20
C11789 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.CLK 0.235f
C11790 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 2.11e-19
C11791 VDD100 a_45815_n1102# 3.56e-19
C11792 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_26426_11196# 9.1e-19
C11793 VDD96 a_30589_n2952# 3.14e-19
C11794 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 2.81e-20
C11795 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB a_48017_9057# 3.25e-19
C11796 RST a_25472_5018# 0.00186f
C11797 CLK_div_96_mag_0.JK_FF_mag_0.Q CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.267f
C11798 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 2.92f
C11799 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN 0.431f
C11800 VDD110 a_47760_n15585# 3.14e-19
C11801 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 0.888f
C11802 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 0.0496f
C11803 VDD110 a_49042_n16682# 3.14e-19
C11804 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 8.36e-19
C11805 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_28268_n6266# 0.069f
C11806 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 a_22575_n287# 0.011f
C11807 RST a_37955_n9984# 0.00114f
C11808 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN 0.00517f
C11809 F1 a_36202_6265# 3.58e-20
C11810 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.994f
C11811 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 6.18e-19
C11812 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 a_22685_11196# 0.00859f
C11813 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB 0.876f
C11814 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_23403_10099# 1.75e-19
C11815 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_49991_n2243# 1.17e-20
C11816 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 0.00656f
C11817 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT a_51646_1671# 0.0203f
C11818 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_55156_n18696# 0.00118f
C11819 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 a_34736_n15539# 1.52e-20
C11820 a_48023_n7840# CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 2.51e-19
C11821 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 Vdiv108 0.00531f
C11822 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_52002_n15583# 0.069f
C11823 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 3.81e-19
C11824 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT a_33652_n13270# 0.0135f
C11825 F2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 7.34e-20
C11826 a_41284_n14596# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT 0.0732f
C11827 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 7.24e-19
C11828 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.VOUT CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN 0.106f
C11829 RST a_45730_10154# 0.00186f
C11830 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_53303_n16728# 5.5e-19
C11831 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 5.63e-21
C11832 Vdiv108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 4.81e-22
C11833 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 1.88e-19
C11834 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.338f
C11835 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.107f
C11836 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 5.55e-21
C11837 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.00488f
C11838 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 1.03f
C11839 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_36673_n8887# 3.33e-19
C11840 CLK_div_96_mag_0.JK_FF_mag_0.QB a_23552_n1789# 2.96e-19
C11841 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.652f
C11842 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 1.89e-21
C11843 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_51983_7381# 5.1e-20
C11844 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_33405_7558# 3.16e-19
C11845 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT 3.39e-20
C11846 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK a_53304_n18696# 2.94e-19
C11847 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.652f
C11848 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB a_50470_9057# 2.96e-19
C11849 a_51492_2768# a_51652_2768# 0.0504f
C11850 a_23956_n14213# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN 0.069f
C11851 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_54004_5143# 0.0733f
C11852 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 6.37e-19
C11853 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.122f
C11854 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 a_22559_n7106# 6.43e-21
C11855 Vdiv110 CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 0.0959f
C11856 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 CLK_div_96_mag_0.JK_FF_mag_2.Q 0.00113f
C11857 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.398f
C11858 RST a_25800_n18723# 7.78e-19
C11859 Vdiv100 a_37999_n1222# 3.41e-19
C11860 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_30881_n18723# 0.0059f
C11861 Vdiv96 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_1.IN2 0.0056f
C11862 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0626f
C11863 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 5.09e-24
C11864 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 a_35747_280# 0.00372f
C11865 VDD90 Vdiv90 0.117f
C11866 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT a_33405_7558# 0.00894f
C11867 a_25328_n15535# a_25488_n15535# 0.0504f
C11868 VDD108 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.399f
C11869 RST CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.0238f
C11870 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.41f
C11871 CLK_div_100_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 5.13e-19
C11872 a_30210_n13332# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 4.33e-21
C11873 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 a_48268_n1102# 6.06e-21
C11874 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 0.149f
C11875 RST CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 0.00425f
C11876 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0894f
C11877 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C11878 RST a_28737_n2996# 0.00243f
C11879 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 0.0101f
C11880 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.0622f
C11881 VDD100 a_44170_2768# 3.14e-19
C11882 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_23967_10099# 1.41e-20
C11883 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 2.25e-19
C11884 CLK CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 1.29e-19
C11885 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_26965_n18723# 0.00118f
C11886 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 2.51e-19
C11887 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.397f
C11888 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_47252_6240# 9.32e-19
C11889 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0634f
C11890 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.394f
C11891 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_45541_n18696# 0.011f
C11892 RST CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.147f
C11893 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_50875_n2243# 8.64e-19
C11894 CLK_div_105_mag_0.CLK_div_10_mag_1.CLK CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB 0.307f
C11895 RST CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.0783f
C11896 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 6.03e-20
C11897 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK 0.341f
C11898 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT a_29187_n15493# 0.0195f
C11899 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_1.IN2 0.109f
C11900 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 8.16e-20
C11901 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K 0.487f
C11902 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 m3_20882_n11188# 0.00197f
C11903 CLK CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.00364f
C11904 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_54503_1671# 0.00119f
C11905 CLK_div_90_mag_0.CLK_div_10_mag_0.CLK a_22461_6115# 0.00939f
C11906 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C11907 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.0881f
C11908 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 5.05f
C11909 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_50304_n16724# 1.46e-19
C11910 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 0.198f
C11911 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.153f
C11912 F2 dec3x8_ibr_mag_0.and_3_ibr_6.nand3_mag_ibr_0.OUT 0.299f
C11913 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.00182f
C11914 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 0.16f
C11915 VDD110 CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 0.329f
C11916 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB a_52923_9057# 0.0114f
C11917 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00105f
C11918 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_25508_n8734# 1.43e-19
C11919 a_50827_5143# a_50987_5143# 0.0504f
C11920 VDD90 a_25478_6115# 2.66e-19
C11921 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN 1.56e-21
C11922 CLK_div_93_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 6.11e-19
C11923 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_47134_n2243# 1.5e-20
C11924 CLK a_51551_5187# 4.86e-19
C11925 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 a_26189_n6010# 0.016f
C11926 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_51239_n5724# 4.52e-20
C11927 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT 0.0357f
C11928 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_46980_n1146# 0.00876f
C11929 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.159f
C11930 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_29301_n2996# 9.1e-19
C11931 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 a_50923_n10161# 0.0102f
C11932 RST CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 6.71e-19
C11933 RST CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 8.93e-19
C11934 CLK a_55357_n20487# 0.00233f
C11935 VDD93 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 5.5e-19
C11936 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 1.19e-19
C11937 Vdiv108 mux_8x1_ibr_0.mux_2x1_ibr_0.I0 0.0259f
C11938 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 0.338f
C11939 VDD99 CLK_div_96_mag_0.JK_FF_mag_4.QB 0.0523f
C11940 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_29116_398# 0.0697f
C11941 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 1.41e-20
C11942 a_50287_n18696# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.0203f
C11943 CLK_div_96_mag_0.JK_FF_mag_3.Q a_28828_1497# 0.0103f
C11944 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.343f
C11945 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 8.16e-20
C11946 a_53940_n10161# m3_20882_n11188# 4.3e-19
C11947 F0 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 0.395f
C11948 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 a_47863_10154# 8.64e-19
C11949 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 1f
C11950 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_32230_5018# 0.00696f
C11951 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 a_54615_9057# 2.79e-20
C11952 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 2.17e-19
C11953 RST CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.288f
C11954 CLK CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 0.151f
C11955 CLK_div_96_mag_0.JK_FF_mag_4.QB a_26096_3016# 0.00696f
C11956 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K 0.0685f
C11957 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT 0.0622f
C11958 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.652f
C11959 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_47994_n18696# 1.43e-19
C11960 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 5.98e-20
C11961 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT 0.338f
C11962 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 6.82e-19
C11963 a_48148_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.00696f
C11964 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_54302_n1102# 0.0059f
C11965 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.00205f
C11966 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 0.3f
C11967 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.055f
C11968 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT 0.0622f
C11969 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT a_52225_n13362# 0.0105f
C11970 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0854f
C11971 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_25292_10099# 4.52e-20
C11972 VDD90 a_26984_10099# 2.65e-19
C11973 a_47911_2768# Vdiv110 5.84e-19
C11974 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 1.48e-19
C11975 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_44846_10154# 8.64e-19
C11976 CLK_div_96_mag_0.JK_FF_mag_2.Q a_25644_n2996# 0.00789f
C11977 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 1.74e-19
C11978 a_43671_7266# a_43831_7266# 0.186f
C11979 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_23019_5018# 0.0203f
C11980 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 4.44e-20
C11981 VDD99 a_38454_6265# 0.00137f
C11982 VDD96 a_25375_354# 5.99e-19
C11983 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00183f
C11984 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_46889_9057# 7.4e-19
C11985 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN 1.61e-19
C11986 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_54746_n17599# 0.069f
C11987 CLK_div_105_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN 4.85e-20
C11988 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_53255_n5765# 0.00119f
C11989 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.121f
C11990 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.529f
C11991 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN a_30165_n6282# 0.069f
C11992 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.125f
C11993 CLK a_47196_n15629# 0.0105f
C11994 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.00137f
C11995 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_105_mag_0.CLK_div_10_mag_1.CLK 0.235f
C11996 RST a_39690_n8887# 1.9e-19
C11997 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 3.8e-20
C11998 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 a_51646_1671# 0.0101f
C11999 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_2.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 1.14e-20
C12000 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 0.00574f
C12001 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_44235_6240# 0.00392f
C12002 VDD110 a_55357_n20487# 0.0407f
C12003 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 1.93e-19
C12004 RST Vdiv110 4.79f
C12005 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 a_25662_n9875# 0.0101f
C12006 CLK a_33513_10099# 0.0101f
C12007 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 0.0126f
C12008 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.00132f
C12009 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN 1.36e-19
C12010 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 2.59e-21
C12011 a_47050_n7372# CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 4.98e-20
C12012 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 0.0018f
C12013 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_22559_n7106# 0.0202f
C12014 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK 0.937f
C12015 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT a_26052_n15491# 0.0195f
C12016 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN a_43719_n120# 2.85e-20
C12017 RST a_44687_n1102# 0.0012f
C12018 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_53221_2768# 0.00378f
C12019 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.395f
C12020 VDD108 a_46614_n6273# 2.21e-19
C12021 CLK_div_105_mag_0.CLK_div_10_mag_1.CLK CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.267f
C12022 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.231f
C12023 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C12024 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.69f
C12025 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.404f
C12026 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_52139_n18696# 0.00118f
C12027 CLK_div_108_new_mag_0.JK_FF_mag_1.QB a_50111_n5768# 0.00392f
C12028 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.00975f
C12029 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 2.81e-20
C12030 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.231f
C12031 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 a_48747_10154# 0.00119f
C12032 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 a_47723_574# 2.36e-22
C12033 RST a_25662_n9875# 0.00187f
C12034 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_30341_5062# 0.0811f
C12035 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 7.35e-19
C12036 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_31731_n16632# 1.5e-20
C12037 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 a_29144_n8735# 3.59e-20
C12038 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.122f
C12039 RST a_28490_11196# 0.00371f
C12040 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT a_48747_10154# 0.0202f
C12041 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_46810_n10116# 0.069f
C12042 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.16f
C12043 VDD96 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 0.49f
C12044 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0893f
C12045 CLK CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.235f
C12046 RST a_44885_n6273# 8.99e-19
C12047 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 7.24e-19
C12048 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 0.198f
C12049 VDD100 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0077f
C12050 VDD108 a_49951_n5768# 0.00484f
C12051 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_31445_n18723# 0.0202f
C12052 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 4.08f
C12053 a_25465_n6010# a_25625_n6010# 0.0504f
C12054 CLK CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 6.64e-19
C12055 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_30210_n13332# 8.5e-20
C12056 F2 a_38561_880# 0.0144f
C12057 VDD96 CLK_div_96_mag_0.JK_FF_mag_0.Q 2.07f
C12058 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT 0.768f
C12059 CLK_div_90_mag_0.CLK_div_10_mag_0.CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 6.64e-19
C12060 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00118f
C12061 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 1.5e-20
C12062 VDD100 a_45251_n1102# 3.14e-19
C12063 CLK CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_0.OUT 0.267f
C12064 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_26266_11196# 2.88e-20
C12065 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.75f
C12066 VDD96 a_30025_n2952# 3.14e-19
C12067 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB a_47453_9057# 2.96e-19
C12068 CLK_div_96_mag_0.JK_FF_mag_5.QB a_23145_810# 0.00695f
C12069 a_49997_n1146# a_50157_n1146# 0.0504f
C12070 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_22620_n9884# 2.88e-20
C12071 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 a_31129_n6271# 2.43e-19
C12072 RST a_25312_5018# 0.00186f
C12073 a_47050_n7372# CLK_div_108_new_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.069f
C12074 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 3.48e-19
C12075 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0822f
C12076 CLK_div_100_mag_0.CLK_div_10_mag_1.CLK CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 3.1e-22
C12077 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_45730_10154# 0.0202f
C12078 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_26663_398# 0.0059f
C12079 VDD100 a_45787_574# 3.14e-19
C12080 a_47754_n16726# a_47914_n16726# 0.0504f
C12081 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.JK_FF_mag_5.QB 0.307f
C12082 VDD110 a_48478_n16682# 3.14e-19
C12083 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB 0.179f
C12084 Vdiv110 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 3.13e-20
C12085 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 a_27342_n1855# 0.00372f
C12086 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 1.53e-19
C12087 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.0591f
C12088 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 a_22011_n287# 0.00118f
C12089 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 4.44e-20
C12090 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_1.IN2 a_22575_n287# 0.069f
C12091 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 a_27227_398# 0.069f
C12092 a_35026_n18723# a_35186_n18723# 0.0504f
C12093 RST a_37391_n9984# 0.00164f
C12094 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0038f
C12095 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K 2.37f
C12096 F1 a_36042_6265# 0.00132f
C12097 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB 6.93e-19
C12098 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 a_22121_11196# 0.0157f
C12099 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_22839_10099# 2.96e-19
C12100 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0219f
C12101 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_54592_n18696# 0.011f
C12102 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT a_51486_1671# 0.0732f
C12103 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_36588_n15495# 0.00118f
C12104 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 a_22461_6115# 2.79e-20
C12105 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.122f
C12106 VDD mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 0.405f
C12107 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C12108 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C12109 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C12110 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.00105f
C12111 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 3.01e-20
C12112 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT a_52951_7381# 3.92e-20
C12113 a_41124_n14596# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT 0.0202f
C12114 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_52156_n16680# 0.0157f
C12115 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_23409_11196# 0.00695f
C12116 RST a_45570_10154# 0.00186f
C12117 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_54028_n18696# 0.00378f
C12118 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 2.36f
C12119 VDD99 a_30050_n13332# 5.08e-19
C12120 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C12121 CLK_div_96_mag_0.JK_FF_mag_3.Q a_28546_n743# 0.0108f
C12122 RST CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 0.0546f
C12123 CLK_div_96_mag_0.JK_FF_mag_5.Q CLK_div_96_mag_0.JK_FF_mag_5.QB 1.97f
C12124 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 9.24e-20
C12125 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 Vdiv110 0.00131f
C12126 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 8.27e-19
C12127 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 4.68e-20
C12128 CLK_div_96_mag_0.JK_FF_mag_0.QB a_22988_n1789# 3.33e-19
C12129 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_36109_n8931# 0.00392f
C12130 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.0591f
C12131 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_51015_7381# 0.069f
C12132 Vdiv99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 0.0303f
C12133 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.JK_FF_mag_3.Q 0.0449f
C12134 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_33245_7558# 3.16e-19
C12135 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 a_51486_1671# 0.00119f
C12136 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 0.179f
C12137 VDD90 dec3x8_ibr_mag_0.and_3_ibr_5.IN3 0.118f
C12138 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_35192_n17626# 1.17e-20
C12139 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C12140 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 4.36e-20
C12141 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0129f
C12142 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 2.86e-19
C12143 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB a_49906_9057# 0.0114f
C12144 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 2.37f
C12145 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_53844_5143# 0.0203f
C12146 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 8.58e-20
C12147 CLK_div_108_new_mag_0.JK_FF_mag_1.QB CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0592f
C12148 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT 2.57e-20
C12149 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 3.72e-19
C12150 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 1.3f
C12151 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 4.44e-20
C12152 dec3x8_ibr_mag_0.and_3_ibr_5.nand3_mag_ibr_0.OUT dec3x8_ibr_mag_0.and_3_ibr_6.nand3_mag_ibr_0.OUT 6.7e-19
C12153 VDD93 a_21841_n6009# 3.14e-19
C12154 RST a_25640_n18723# 6.43e-19
C12155 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 0.0579f
C12156 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT Vdiv110 0.00521f
C12157 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.69f
C12158 VDD90 a_33405_7558# 0.0407f
C12159 CLK Vdiv105 0.298f
C12160 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT a_33245_7558# 0.0294f
C12161 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 0.00158f
C12162 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.741f
C12163 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 5.7e-19
C12164 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 a_32076_6159# 6.43e-21
C12165 a_55156_n18696# CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 2.1e-20
C12166 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.00518f
C12167 RST a_28577_n2996# 0.00243f
C12168 RST a_54028_n18696# 2.78e-19
C12169 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 0.0231f
C12170 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.122f
C12171 a_29053_5018# a_29213_5018# 0.0504f
C12172 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 1.33e-20
C12173 VDD100 a_43606_2768# 3.14e-19
C12174 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.0189f
C12175 F0 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 0.378f
C12176 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 0.25f
C12177 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_47092_6240# 0.00876f
C12178 RST a_55161_n15587# 6.17e-19
C12179 VDD99 a_25800_n18723# 2.21e-19
C12180 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_44977_n18696# 1.43e-19
C12181 RST a_55315_n16684# 0.00106f
C12182 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 9.4e-19
C12183 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_52385_n13362# 0.0504f
C12184 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.99e-19
C12185 CLK_div_96_mag_0.JK_FF_mag_0.QB CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.28f
C12186 CLK_div_90_mag_0.CLK_div_10_mag_0.CLK a_22301_6115# 0.0101f
C12187 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_53939_1671# 1.43e-19
C12188 a_43872_9057# CLK_div_105_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 2.1e-20
C12189 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.303f
C12190 CLK_div_108_new_mag_0.JK_FF_mag_0.QB a_55101_n6818# 0.0811f
C12191 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 1.08f
C12192 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.198f
C12193 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.395f
C12194 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0501f
C12195 VDD105 dec3x8_ibr_mag_0.and_3_ibr_6.nand3_mag_ibr_0.OUT 0.15f
C12196 VDD99 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 3.45e-20
C12197 F2 a_38454_6265# 0.00981f
C12198 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_44953_5143# 2.88e-20
C12199 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C12200 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_24944_n8778# 0.00119f
C12201 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 9.24e-20
C12202 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.106f
C12203 VDD90 a_25318_6115# 3.78e-19
C12204 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.16f
C12205 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_46974_n2243# 1.17e-20
C12206 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.00418f
C12207 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_50675_n5724# 0.0202f
C12208 CLK a_50987_5143# 4.68e-19
C12209 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 a_25625_n6010# 0.0102f
C12210 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 0.296f
C12211 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 4.67e-22
C12212 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 a_50763_n10161# 0.0101f
C12213 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_28737_n2996# 0.0731f
C12214 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 0.0683f
C12215 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.643f
C12216 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.653f
C12217 CLK a_55197_n20487# 0.00204f
C12218 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 0.79f
C12219 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.119f
C12220 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.105f
C12221 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_54414_6284# 0.0059f
C12222 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.192f
C12223 VDD110 Vdiv105 0.123f
C12224 RST CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.602f
C12225 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 0.109f
C12226 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 1.54e-19
C12227 VDD mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 0.405f
C12228 a_50287_n18696# a_50447_n18696# 0.0504f
C12229 a_53780_n10161# m3_20882_n11188# 4.3e-19
C12230 RST CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.132f
C12231 Vdiv105 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 0.131f
C12232 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 0.66f
C12233 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K a_32070_5018# 0.00695f
C12234 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 1.29e-19
C12235 CLK_div_96_mag_0.JK_FF_mag_4.QB a_25532_3016# 0.00964f
C12236 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_44885_n6273# 0.0059f
C12237 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0343f
C12238 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 0.0126f
C12239 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB 2.1e-19
C12240 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 0.00656f
C12241 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 2.86e-19
C12242 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 0.198f
C12243 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 a_44123_n1146# 2.79e-20
C12244 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K 8.05e-19
C12245 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_48712_n17599# 0.00378f
C12246 a_47988_n17599# CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.00695f
C12247 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 a_45618_2768# 0.00117f
C12248 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT 8.48e-20
C12249 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 2.33e-19
C12250 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 9.05e-22
C12251 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_53738_n1102# 0.0697f
C12252 CLK_div_96_mag_0.JK_FF_mag_2.QB CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.343f
C12253 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_44888_1671# 0.0697f
C12254 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0209f
C12255 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.768f
C12256 VDD110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.395f
C12257 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT a_49488_n13383# 6.43e-19
C12258 RST CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0119f
C12259 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 0.175f
C12260 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_28093_n18723# 0.0202f
C12261 a_47751_2768# Vdiv110 5.84e-19
C12262 VDD90 a_26420_10099# 3.14e-19
C12263 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_27381_n699# 0.00372f
C12264 CLK_div_96_mag_0.JK_FF_mag_2.Q a_25484_n2996# 0.00335f
C12265 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB 0.169f
C12266 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_22455_5018# 1.5e-20
C12267 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0622f
C12268 VDD99 a_38294_6265# 0.00174f
C12269 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.298f
C12270 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 0.0175f
C12271 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 0.0147f
C12272 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.132f
C12273 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_45000_9057# 0.0697f
C12274 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_28817_n18723# 8.64e-19
C12275 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN a_29214_n6271# 4.56e-21
C12276 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB 1.76e-21
C12277 CLK a_47036_n15629# 0.0114f
C12278 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 7.08e-20
C12279 CLK_div_90_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN a_29087_8532# 3.25e-19
C12280 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 a_22551_n16006# 0.0111f
C12281 RST CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 3.84e-20
C12282 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 0.00916f
C12283 RST a_39126_n8931# 6.43e-19
C12284 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.468f
C12285 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 a_51486_1671# 0.00939f
C12286 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 a_25478_6115# 2.79e-20
C12287 VDD99 a_33429_n15491# 3.56e-19
C12288 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 0.00121f
C12289 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_26636_n8734# 0.00372f
C12290 VDD110 a_55197_n20487# 0.234f
C12291 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 a_25502_n9875# 0.0102f
C12292 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 a_34890_n16636# 4.28e-19
C12293 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_46081_5187# 0.0811f
C12294 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_47858_n2243# 8.64e-19
C12295 CLK a_33353_10099# 0.00939f
C12296 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 0.671f
C12297 Vdiv100 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 0.00288f
C12298 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT a_21995_n7106# 4.52e-20
C12299 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN 0.125f
C12300 RST a_44123_n1146# 9.5e-19
C12301 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 1.83e-19
C12302 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_23552_n1789# 4.52e-20
C12303 VDD108 a_45449_n6273# 3.56e-19
C12304 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0263f
C12305 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_51575_n18696# 0.011f
C12306 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 1.88e-19
C12307 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 0.0725f
C12308 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT 0.343f
C12309 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.159f
C12310 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C12311 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 a_48587_10154# 0.00166f
C12312 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_30244_398# 0.00118f
C12313 RST a_25502_n9875# 0.00171f
C12314 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT 1.2e-19
C12315 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_29777_5062# 0.00964f
C12316 CLK_div_96_mag_0.JK_FF_mag_3.QB a_30435_n1855# 0.0114f
C12317 VDD96 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.00586f
C12318 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 CLK_div_96_mag_0.JK_FF_mag_3.QB 0.0015f
C12319 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 7.94e-20
C12320 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT a_31571_n16632# 1.17e-20
C12321 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_33744_n17626# 0.0036f
C12322 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT a_48587_10154# 0.0731f
C12323 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_46246_n10116# 0.00372f
C12324 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0169f
C12325 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.0521f
C12326 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 3.84e-20
C12327 VDD110 dec3x8_ibr_mag_0.and_3_ibr_2.nand3_mag_ibr_0.OUT 1.51e-19
C12328 VDD93 Vdiv90 1.55f
C12329 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 1.76f
C12330 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 3.53e-19
C12331 RST a_44321_n6273# 1.21e-19
C12332 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 a_46774_n6273# 2.79e-20
C12333 VDD99 Vdiv110 0.00752f
C12334 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 0.0241f
C12335 RST CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.00217f
C12336 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_30881_n18723# 4.52e-20
C12337 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C12338 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 1.83e-19
C12339 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.199f
C12340 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K 0.0432f
C12341 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 a_49122_n18696# 4.52e-20
C12342 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.0591f
C12343 VDD100 Vdiv110 0.546f
C12344 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0132f
C12345 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_30050_n13332# 1.32e-19
C12346 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 a_48469_1671# 0.00119f
C12347 Vdiv90 F0 0.0667f
C12348 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB 0.28f
C12349 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 9.22e-20
C12350 VDD100 a_44687_n1102# 3.14e-19
C12351 RST CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.155f
C12352 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 0.209f
C12353 CLK_div_96_mag_0.JK_FF_mag_3.Q a_28743_n1899# 2.79e-20
C12354 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB 0.25f
C12355 CLK_div_96_mag_0.JK_FF_mag_0.Q CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 9.71e-20
C12356 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB a_46889_9057# 0.0114f
C12357 CLK_div_96_mag_0.JK_FF_mag_5.QB a_22985_810# 0.00696f
C12358 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 0.395f
C12359 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_22460_n9884# 9.1e-19
C12360 RST a_24307_5062# 9.66e-19
C12361 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0894f
C12362 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_45570_10154# 0.0731f
C12363 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 a_50111_n5768# 1.07e-20
C12364 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_26099_398# 0.0697f
C12365 VDD110 a_47036_n15629# 2.21e-19
C12366 CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 1.82e-19
C12367 Vdiv93 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_1.IN2 0.109f
C12368 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.231f
C12369 Vdiv93 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK 3.81e-20
C12370 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 3.28e-19
C12371 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 a_26778_n1855# 0.069f
C12372 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00183f
C12373 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 1.96f
C12374 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 0.00121f
C12375 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 2.31e-19
C12376 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 a_48475_2768# 1.46e-19
C12377 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_1.IN2 a_22011_n287# 0.00372f
C12378 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 9.83e-19
C12379 VDD99 a_30760_n20290# 0.165f
C12380 RST a_36827_n10028# 0.00228f
C12381 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 0.391f
C12382 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.69f
C12383 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C12384 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.231f
C12385 a_28663_n17626# a_28823_n17626# 0.0504f
C12386 a_52811_1671# CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 2.05e-19
C12387 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_22275_10099# 0.012f
C12388 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.122f
C12389 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 9.62e-20
C12390 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 2.48e-20
C12391 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT a_50922_1671# 0.00378f
C12392 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_54028_n18696# 1.43e-19
C12393 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00174f
C12394 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_36024_n15495# 0.011f
C12395 VDD a_36873_280# 0.00444f
C12396 CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00335f
C12397 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0854f
C12398 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 0.0267f
C12399 a_41124_n14596# a_41284_n14596# 0.0504f
C12400 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_51592_n16680# 0.00859f
C12401 RST a_45006_10154# 0.00169f
C12402 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.121f
C12403 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_23249_11196# 0.00696f
C12404 VDD99 dec3x8_ibr_mag_0.and_3_ibr_1.nand3_mag_ibr_0.OUT 0.0247f
C12405 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB a_53945_2768# 0.00695f
C12406 VDD99 a_22544_n13819# 3.14e-19
C12407 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 8.58e-20
C12408 CLK_div_96_mag_0.JK_FF_mag_3.Q a_28386_n743# 0.00749f
C12409 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 4.88e-19
C12410 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 a_29298_n9832# 0.0036f
C12411 RST CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_1.IN2 0.00682f
C12412 a_28335_6115# a_28495_6115# 0.0504f
C12413 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB 0.307f
C12414 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.038f
C12415 VDD110 CLK_div_93_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 7.6e-19
C12416 F0 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 0.198f
C12417 RST a_45724_9057# 8.64e-19
C12418 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.487f
C12419 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_53892_n2243# 2.88e-20
C12420 CLK_div_96_mag_0.JK_FF_mag_0.QB a_22424_n1833# 0.00392f
C12421 RST CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.684f
C12422 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN a_33245_7558# 2.85e-20
C12423 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB 1e-19
C12424 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.378f
C12425 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 a_50922_1671# 1.43e-19
C12426 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 a_32455_n16632# 8.64e-19
C12427 a_27856_n8779# a_28016_n8779# 0.0504f
C12428 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0432f
C12429 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_35032_n17626# 1.5e-20
C12430 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 a_26250_1919# 0.0697f
C12431 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.0626f
C12432 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C12433 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.11f
C12434 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_53280_5143# 1.5e-20
C12435 CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0263f
C12436 CLK_div_96_mag_0.JK_FF_mag_2.Q a_29307_n1855# 6.43e-21
C12437 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.397f
C12438 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.43e-20
C12439 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 3.57e-20
C12440 VDD93 a_21277_n6009# 3.14e-19
C12441 dec3x8_ibr_mag_0.and_3_ibr_5.nand3_mag_ibr_0.OUT a_38454_6265# 3.58e-20
C12442 RST a_25076_n18723# 2.97e-19
C12443 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.00264f
C12444 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 0.16f
C12445 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN 2.44e-21
C12446 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.122f
C12447 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 a_47341_1671# 0.069f
C12448 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_44321_n6273# 0.00378f
C12449 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.00733f
C12450 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_27324_5062# 0.0811f
C12451 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 8.83e-19
C12452 VDD90 a_33245_7558# 0.234f
C12453 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 2.6e-19
C12454 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.999f
C12455 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.768f
C12456 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT a_30209_7256# 0.00138f
C12457 RST CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00722f
C12458 VDD110 a_50447_n18696# 2.66e-19
C12459 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 a_31512_6115# 0.00939f
C12460 VDD93 dec3x8_ibr_mag_0.and_3_ibr_4.nand3_mag_ibr_0.OUT 0.149f
C12461 CLK CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 3.92e-21
C12462 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0352f
C12463 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 1.54e-21
C12464 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.338f
C12465 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 a_47140_n1146# 2.79e-20
C12466 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 9.48e-20
C12467 RST a_27496_n2952# 0.00122f
C12468 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.122f
C12469 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 1.55e-19
C12470 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.338f
C12471 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 3.41e-19
C12472 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.00586f
C12473 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.125f
C12474 VDD110 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 7.81e-22
C12475 F0 dec3x8_ibr_mag_0.and_3_ibr_4.nand3_mag_ibr_0.OUT 0.285f
C12476 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.00118f
C12477 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C12478 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.768f
C12479 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.121f
C12480 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB 0.0386f
C12481 RST a_54597_n15587# 6.17e-19
C12482 VDD90 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.878f
C12483 RST a_54751_n16684# 0.00106f
C12484 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 6.82e-19
C12485 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 5.08e-20
C12486 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0135f
C12487 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 a_52225_n13362# 0.0186f
C12488 a_40375_n7552# CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.4e-19
C12489 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB 0.904f
C12490 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN 6.2e-19
C12491 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_43719_n120# 9.21e-20
C12492 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_53375_1671# 0.011f
C12493 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.00165f
C12494 CLK_div_108_new_mag_0.JK_FF_mag_0.QB a_54537_n6818# 0.00964f
C12495 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.579f
C12496 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 0.493f
C12497 VDD105 a_38454_6265# 0.00174f
C12498 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.0213f
C12499 VDD mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 0.405f
C12500 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB a_33245_7558# 5.07e-21
C12501 F2 a_38294_6265# 0.00237f
C12502 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 m3_20882_n11188# 1.48e-19
C12503 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_44793_5143# 9.1e-19
C12504 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.108f
C12505 a_23129_n6009# a_23289_n6009# 0.0504f
C12506 VDD100 a_54669_2768# 0.0132f
C12507 RST a_45612_1671# 8.64e-19
C12508 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0262f
C12509 VDD90 a_24153_6159# 3.56e-19
C12510 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_32640_6159# 4.52e-20
C12511 CLK a_23289_n6009# 0.00165f
C12512 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 2.48e-19
C12513 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 a_25465_n6010# 0.0101f
C12514 CLK a_50827_5143# 4.68e-19
C12515 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 0.00395f
C12516 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.16f
C12517 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 a_50199_n10117# 0.00859f
C12518 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_2.OUT a_28577_n2996# 0.0202f
C12519 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.0576f
C12520 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.00109f
C12521 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 a_43671_7266# 0.019f
C12522 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.11f
C12523 VDD96 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.754f
C12524 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 a_23283_n7106# 4.47e-19
C12525 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_53850_6284# 0.0697f
C12526 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0215f
C12527 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.457f
C12528 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 7.08e-20
C12529 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0718f
C12530 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB 0.348f
C12531 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 0.00656f
C12532 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 1.32f
C12533 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 0.102f
C12534 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_51764_10154# 2.81e-19
C12535 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN 0.0609f
C12536 VDD F1 5.05f
C12537 RST CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.023f
C12538 a_53216_n10117# m3_20882_n11188# 4.41e-19
C12539 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.235f
C12540 RST CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN 0.0239f
C12541 CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 0.0445f
C12542 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 a_36109_n8931# 2.79e-20
C12543 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 a_53487_9057# 6.06e-21
C12544 VDD96 CLK_div_96_mag_0.JK_FF_mag_2.QB 0.92f
C12545 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.529f
C12546 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT a_29059_6159# 0.00378f
C12547 CLK_div_96_mag_0.JK_FF_mag_4.QB a_24968_3016# 0.0811f
C12548 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_44321_n6273# 0.0697f
C12549 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.303f
C12550 Vdiv99 a_35949_n8931# 8.56e-19
C12551 RST Vdiv99 0.437f
C12552 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 0.397f
C12553 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_52161_n19793# 5.1e-20
C12554 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 a_52385_n13362# 2.84e-20
C12555 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 a_45458_2768# 0.00164f
C12556 VDD93 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 2.57e-19
C12557 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.22f
C12558 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_44324_1671# 0.0059f
C12559 RST a_32301_n15491# 3.68e-20
C12560 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 0.199f
C12561 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.122f
C12562 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00391f
C12563 F2 Vdiv110 0.0601f
C12564 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 3.21e-20
C12565 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN 8.18e-19
C12566 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB 7.08e-20
C12567 a_47187_2768# Vdiv110 6.25e-19
C12568 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_27529_n18723# 4.52e-20
C12569 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB a_46755_574# 1.45e-20
C12570 VDD90 a_25856_10099# 3.14e-19
C12571 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_26817_n699# 0.069f
C12572 F0 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 0.162f
C12573 RST a_51205_n7921# 7.58e-19
C12574 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0592f
C12575 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_46105_n18696# 4.52e-20
C12576 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 0.829f
C12577 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 1f
C12578 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_22295_5018# 1.17e-20
C12579 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.CLK 0.149f
C12580 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_51439_n2199# 0.0036f
C12581 VDD108 Vdiv110 0.212f
C12582 VDD96 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.391f
C12583 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT a_33204_6159# 1.54e-19
C12584 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.857f
C12585 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 a_29751_n15493# 0.0059f
C12586 CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 a_25364_n19822# 7.48e-20
C12587 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 dec3x8_ibr_mag_0.and_3_ibr_6.nand3_mag_ibr_0.OUT 3.53e-19
C12588 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_44436_9057# 0.0059f
C12589 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 0.321f
C12590 F2 a_39124_280# 2.62e-19
C12591 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 8.28e-20
C12592 CLK a_45753_n15583# 9.34e-19
C12593 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 0.0172f
C12594 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 1.49e-21
C12595 RST a_38966_n8931# 7.78e-19
C12596 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C12597 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0175f
C12598 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK a_39120_n10028# 0.00164f
C12599 Vdiv110 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 0.0263f
C12600 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.012f
C12601 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.0435f
C12602 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00166f
C12603 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 1.01e-20
C12604 CLK_div_96_mag_0.JK_FF_mag_4.Q CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 1.48e-20
C12605 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 a_50922_1671# 6.43e-21
C12606 VDD99 a_32865_n15491# 3.14e-19
C12607 RST CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0683f
C12608 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_26072_n8734# 0.069f
C12609 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN a_22551_n16006# 0.069f
C12610 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 2.25e-19
C12611 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 a_34730_n16636# 5.5e-19
C12612 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 5.45e-20
C12613 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 a_24938_n9875# 0.00789f
C12614 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_45517_5187# 0.00964f
C12615 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.0463f
C12616 CLK a_32789_10099# 6.43e-21
C12617 VDD93 dec3x8_ibr_mag_0.and_3_ibr_5.IN3 0.292f
C12618 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K a_45787_574# 0.0027f
C12619 RST a_43963_n1146# 8.88e-19
C12620 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.121f
C12621 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.103f
C12622 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_22988_n1789# 0.0202f
C12623 a_37801_n8887# CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 4.52e-20
C12624 VDD108 a_44885_n6273# 3.14e-19
C12625 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 CLK_div_96_mag_0.JK_FF_mag_3.Q 1.86e-21
C12626 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 CLK_div_90_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 8.04e-19
C12627 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB 0.198f
C12628 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 2.15e-20
C12629 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_23179_5018# 2.88e-20
C12630 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 a_51011_n18696# 1.43e-19
C12631 a_54615_9057# a_54775_9057# 0.0504f
C12632 dec3x8_ibr_mag_0.and_3_ibr_5.IN3 F0 0.293f
C12633 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 0.285f
C12634 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 a_48023_10154# 3.6e-22
C12635 CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 a_22718_8532# 8.64e-19
C12636 RST a_24938_n9875# 0.00189f
C12637 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_29680_398# 0.011f
C12638 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_29213_5018# 0.00696f
C12639 CLK_div_96_mag_0.JK_FF_mag_3.QB a_29871_n1855# 2.96e-19
C12640 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.233f
C12641 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_108_new_mag_0.JK_FF_mag_1.Q 7.24e-19
C12642 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C12643 F2 dec3x8_ibr_mag_0.and_3_ibr_1.nand3_mag_ibr_0.OUT 0.0191f
C12644 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0846f
C12645 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.401f
C12646 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.00955f
C12647 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT a_48023_10154# 9.1e-19
C12648 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 2.11e-20
C12649 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 1.33e-20
C12650 VDD93 a_33405_7558# 7.01e-19
C12651 a_22575_n287# CLK_div_96_mag_0.JK_FF_mag_0.QB 2.12e-20
C12652 a_21431_n7106# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 2.21e-19
C12653 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.765f
C12654 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.0854f
C12655 RST CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.00721f
C12656 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 8.16e-20
C12657 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 a_47905_1671# 1.43e-19
C12658 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.28f
C12659 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT a_52951_7381# 0.00138f
C12660 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_54866_n1102# 0.00118f
C12661 Vdiv108 a_54947_n5721# 0.069f
C12662 CLK_div_96_mag_0.JK_FF_mag_3.Q CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 2.09f
C12663 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.129f
C12664 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K 3.7f
C12665 VDD100 a_44123_n1146# 2.66e-19
C12666 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT 0.121f
C12667 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN 1e-19
C12668 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.101f
C12669 VDD96 a_29301_n2996# 2.21e-19
C12670 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 0.321f
C12671 CLK_div_96_mag_0.JK_FF_mag_5.QB a_22421_810# 0.00964f
C12672 VDD105 a_45730_10154# 0.00727f
C12673 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_21896_n9884# 0.0731f
C12674 RST a_23743_5062# 9.41e-19
C12675 RST CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN 0.00749f
C12676 a_48620_n5176# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.0811f
C12677 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 0.106f
C12678 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 a_29214_n6271# 3.11e-21
C12679 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT a_26042_6159# 0.00378f
C12680 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_45006_10154# 9.1e-19
C12681 VDD99 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.00219f
C12682 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 a_49951_n5768# 1.37e-20
C12683 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 2.22e-20
C12684 VDD110 a_45753_n15583# 3.56e-19
C12685 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_23179_5018# 8.64e-19
C12686 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.0654f
C12687 Vdiv96 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT 0.0434f
C12688 VDD110 a_47754_n16726# 2.21e-19
C12689 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.122f
C12690 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 1.14f
C12691 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.649f
C12692 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_52293_n17599# 5.02e-20
C12693 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.41f
C12694 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 8.16e-20
C12695 RST a_36667_n10028# 0.00187f
C12696 CLK_div_96_mag_0.JK_FF_mag_4.QB CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 4.46e-20
C12697 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 1.12e-19
C12698 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C12699 RST CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.IN2 9.19e-19
C12700 VDD96 CLK_div_96_mag_0.JK_FF_mag_4.QB 0.917f
C12701 a_43993_n13477# CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.132f
C12702 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 0.158f
C12703 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.0115f
C12704 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.653f
C12705 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_35460_n15495# 1.43e-19
C12706 a_27334_n16588# CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 2.34e-20
C12707 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C12708 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 0.11f
C12709 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_50310_n15627# 2.79e-20
C12710 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.194f
C12711 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_51028_n16724# 0.0101f
C12712 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_22685_11196# 0.00964f
C12713 CLK_div_108_new_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 3.76e-19
C12714 RST a_44846_10154# 0.00128f
C12715 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB a_23123_n7106# 0.00392f
C12716 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 a_26616_n15491# 0.0059f
C12717 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB a_53785_2768# 0.00696f
C12718 CLK_div_93_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_39402_n7788# 0.069f
C12719 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 0.438f
C12720 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.251f
C12721 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K 2.21e-19
C12722 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 0.651f
C12723 RST a_45564_9057# 9.22e-19
C12724 RST CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 0.055f
C12725 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 0.629f
C12726 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 1.51e-19
C12727 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_53732_n2243# 9.1e-19
C12728 a_44475_n5176# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0733f
C12729 Vdiv110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 0.00117f
C12730 RST a_22551_n16006# 3.77e-19
C12731 CLK_div_96_mag_0.JK_FF_mag_4.Q a_26814_1919# 2.79e-20
C12732 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 a_50358_1671# 0.011f
C12733 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_34468_n17626# 0.0203f
C12734 a_50105_n6865# CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 4.06e-19
C12735 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 a_25686_1919# 0.0059f
C12736 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.OUT a_37999_n1222# 0.0964f
C12737 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 0.0432f
C12738 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_53120_5143# 1.17e-20
C12739 CLK_div_96_mag_0.JK_FF_mag_2.Q a_28743_n1899# 0.00939f
C12740 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.0622f
C12741 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.11f
C12742 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_32009_n18723# 0.00392f
C12743 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.36f
C12744 dec3x8_ibr_mag_0.and_3_ibr_5.nand3_mag_ibr_0.OUT a_38294_6265# 6.08e-20
C12745 RST a_24512_n18723# 2.24e-19
C12746 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN 0.111f
C12747 F2 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT 0.00122f
C12748 RST CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 0.133f
C12749 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 a_46777_1671# 0.00372f
C12750 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_26760_5062# 0.00964f
C12751 VDD90 a_30209_7256# 3.14e-19
C12752 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_0.OUT CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0622f
C12753 F2 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT 0.11f
C12754 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 a_51165_n17599# 8.64e-19
C12755 VDD110 a_50287_n18696# 0.00746f
C12756 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN 0.112f
C12757 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 a_31352_6115# 0.0101f
C12758 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB 0.307f
C12759 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_51165_n17599# 0.0101f
C12760 VDD93 a_36202_6265# 0.00167f
C12761 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.0659f
C12762 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN 0.0248f
C12763 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_27227_398# 0.00118f
C12764 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT 2.67e-20
C12765 RST a_53945_2768# 8.64e-19
C12766 RST a_26932_n2952# 0.0012f
C12767 VDD a_39420_6821# 2.21e-19
C12768 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.VOUT CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN 0.00527f
C12769 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.458f
C12770 a_53095_n5765# a_53255_n5765# 0.0504f
C12771 F0 a_36202_6265# 8.64e-19
C12772 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.00481f
C12773 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT a_29144_n8735# 4.52e-20
C12774 VDD99 a_25076_n18723# 3.14e-19
C12775 RST a_54033_n15587# 2.67e-19
C12776 RST a_54187_n16728# 0.002f
C12777 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.0592f
C12778 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_55156_n18696# 4.52e-20
C12779 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT 7.24e-19
C12780 RST CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.0873f
C12781 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K 5.25e-20
C12782 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_33359_11196# 1.46e-19
C12783 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K a_43559_n120# 3.02e-19
C12784 a_26817_n699# CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 5.3e-20
C12785 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_52811_1671# 0.00118f
C12786 CLK_div_108_new_mag_0.JK_FF_mag_0.QB a_53973_n6862# 0.00696f
C12787 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 8.94e-19
C12788 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 0.768f
C12789 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.235f
C12790 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.742f
C12791 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 a_52839_n5# 0.01f
C12792 VDD105 a_38294_6265# 0.00139f
C12793 VDD a_35747_280# 0.00444f
C12794 Vdiv108 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 7.02e-21
C12795 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 5.62e-19
C12796 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_44229_5143# 0.0731f
C12797 VDD100 a_50903_n5# 6e-19
C12798 Vdiv110 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K 8.29e-19
C12799 VDD100 a_54509_2768# 0.00892f
C12800 RST a_45452_1671# 9.22e-19
C12801 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_32076_6159# 0.0202f
C12802 VDD90 a_23589_6159# 3.14e-19
C12803 CLK a_23129_n6009# 0.00165f
C12804 VDD93 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.08f
C12805 CLK a_50263_5143# 0.00111f
C12806 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 a_24901_n6010# 0.00859f
C12807 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.496f
C12808 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 0.018f
C12809 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 a_49635_n10117# 0.0157f
C12810 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB a_32169_n18723# 1.86e-20
C12811 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT 1.17e-19
C12812 a_30315_n15493# CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 4.52e-20
C12813 RST CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 0.139f
C12814 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.CLK 0.149f
C12815 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.107f
C12816 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 a_23123_n7106# 3.43e-19
C12817 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.OUT 4.55e-20
C12818 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 2.61e-20
C12819 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 0.0298f
C12820 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 1.07f
C12821 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_54004_5143# 8.64e-19
C12822 Vdiv105 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 0.1f
C12823 a_23139_n287# CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 3.64e-20
C12824 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.198f
C12825 CLK a_54664_n10161# 0.00117f
C12826 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 Vdiv96 2.53e-19
C12827 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 a_37999_880# 0.00372f
C12828 RST CLK_div_96_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.00347f
C12829 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 0.00127f
C12830 a_52652_n10117# m3_20882_n11188# 4.57e-19
C12831 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.0343f
C12832 RST CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 0.135f
C12833 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 a_52923_9057# 0.069f
C12834 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.0116f
C12835 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 9.8e-20
C12836 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT a_28495_6115# 0.0732f
C12837 VDD108 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.742f
C12838 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 0.0042f
C12839 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_48023_n7840# 1.4e-19
C12840 CLK_div_96_mag_0.JK_FF_mag_2.QB CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 0.0382f
C12841 RST CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.306f
C12842 VDD100 a_45612_1671# 2.21e-19
C12843 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 6.64e-19
C12844 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 4.39e-19
C12845 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 a_52225_n13362# 9.09e-19
C12846 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.267f
C12847 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 0.36f
C12848 Vdiv100 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 0.018f
C12849 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN 1.34e-20
C12850 RST CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.162f
C12851 VDD105 Vdiv110 0.00455f
C12852 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00109f
C12853 VDD93 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 0.391f
C12854 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT 2.11e-20
C12855 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 0.0014f
C12856 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT Vdiv110 0.0268f
C12857 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0014f
C12858 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_2.OUT CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 1.53e-20
C12859 dec3x8_ibr_mag_0.and_3_ibr_1.nand3_mag_ibr_0.OUT dec3x8_ibr_mag_0.and_3_ibr_5.nand3_mag_ibr_0.OUT 0.00141f
C12860 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.11f
C12861 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.768f
C12862 Vdiv108 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.00617f
C12863 VDD90 a_25292_10099# 3.56e-19
C12864 a_46623_2768# Vdiv110 6.45e-19
C12865 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 1.65e-21
C12866 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 2.56e-19
C12867 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C12868 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 5.32e-19
C12869 RST CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.103f
C12870 VDD90 a_33204_6159# 3.56e-19
C12871 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.121f
C12872 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN 7.44e-19
C12873 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 a_29187_n15493# 0.0697f
C12874 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.179f
C12875 CLK_div_105_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 CLK_div_105_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.11f
C12876 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00133f
C12877 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 m3_20882_n11188# 0.00225f
C12878 VDD99 Vdiv99 0.706f
C12879 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.121f
C12880 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB 2.81e-20
C12881 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.0263f
C12882 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K Vdiv110 4e-21
C12883 CLK a_45189_n15583# 9.23e-19
C12884 CLK a_47190_n16726# 0.00164f
C12885 RST CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.00825f
C12886 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00281f
C12887 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_55161_n15587# 0.069f
C12888 RST CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 0.00535f
C12889 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN 2.02e-19
C12890 VDD110 CLK 7.86f
C12891 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK a_38960_n10028# 0.00117f
C12892 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 a_26349_n6010# 0.00613f
C12893 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_55315_n16684# 0.0157f
C12894 VDD99 a_32301_n15491# 3.14e-19
C12895 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 1.05e-19
C12896 CLK_div_108_new_mag_0.JK_FF_mag_1.Q a_53249_n6862# 0.00208f
C12897 CLK a_43993_n13477# 1.64e-20
C12898 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 4.44e-20
C12899 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_44953_5143# 0.00696f
C12900 CLK_div_93_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 6.02e-20
C12901 CLK a_32225_10099# 6.06e-21
C12902 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 a_24778_n9875# 0.00335f
C12903 CLK CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT 6.39e-19
C12904 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 0.00662f
C12905 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB 0.21f
C12906 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 4.09e-19
C12907 CLK_div_100_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_43719_n120# 9.16e-20
C12908 CLK CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 7.81e-19
C12909 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 a_53126_6240# 6.36e-19
C12910 mux_8x1_ibr_0.mux_2x1_ibr_0.I0 a_37999_n1822# 0.069f
C12911 VDD108 a_44321_n6273# 3.14e-19
C12912 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K 0.0823f
C12913 RST CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 0.0204f
C12914 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_54978_6284# 0.00118f
C12915 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 a_53844_5143# 3.6e-22
C12916 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_23019_5018# 9.1e-19
C12917 RST CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.131f
C12918 CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 a_55020_n2199# 0.0157f
C12919 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.00145f
C12920 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.119f
C12921 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 1.97e-19
C12922 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 7.07e-19
C12923 RST a_24778_n9875# 0.00189f
C12924 VDD105 dec3x8_ibr_mag_0.and_3_ibr_1.nand3_mag_ibr_0.OUT 1.25e-20
C12925 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_29116_398# 1.43e-19
C12926 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB a_29053_5018# 0.00695f
C12927 CLK_div_96_mag_0.JK_FF_mag_3.QB a_29307_n1855# 3.33e-19
C12928 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT 0.131f
C12929 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 2.29e-20
C12930 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 1.9e-21
C12931 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT 0.0349f
C12932 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN 0.129f
C12933 F1 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I1 0.0643f
C12934 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT a_47863_10154# 2.88e-20
C12935 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 5.32e-19
C12936 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 2.43e-19
C12937 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB 0.913f
C12938 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 1.22e-19
C12939 VDD93 a_33245_7558# 3.78e-19
C12940 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 7.11e-19
C12941 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 a_48023_n7840# 8.64e-19
C12942 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 6.46e-20
C12943 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.0496f
C12944 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 0.122f
C12945 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 m3_20882_n11188# 0.00275f
C12946 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.14f
C12947 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 2.13e-20
C12948 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 a_28663_n17626# 2.98e-20
C12949 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT 5.05e-20
C12950 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.IN2 4.26e-19
C12951 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 a_47341_1671# 0.011f
C12952 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT a_55179_7683# 0.00894f
C12953 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_54302_n1102# 0.011f
C12954 VDD100 a_43963_n1146# 0.00752f
C12955 RST CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 9.24e-20
C12956 VDD96 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 0.402f
C12957 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT 0.994f
C12958 CLK_div_96_mag_0.JK_FF_mag_5.QB a_21857_810# 0.0811f
C12959 VDD105 a_45570_10154# 0.00299f
C12960 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0622f
C12961 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB a_28657_n18723# 0.00392f
C12962 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_21736_n9884# 0.0202f
C12963 RST a_23179_5018# 0.00186f
C12964 a_48056_n5176# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.00964f
C12965 RST CLK_div_96_mag_0.JK_FF_mag_0.QB 0.229f
C12966 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT a_25478_6115# 0.0732f
C12967 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C12968 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_44846_10154# 2.88e-20
C12969 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 4.24e-20
C12970 CLK_div_96_mag_0.JK_FF_mag_4.Q a_23863_n287# 0.0101f
C12971 VDD99 a_29801_1733# 0.00114f
C12972 VDD110 a_45189_n15583# 3.14e-19
C12973 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00163f
C12974 VDD110 a_47190_n16726# 1.04e-19
C12975 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 0.397f
C12976 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 9.58e-20
C12977 CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 a_24391_n20290# 8.64e-19
C12978 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0622f
C12979 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.121f
C12980 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT 0.305f
C12981 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00169f
C12982 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 9.9e-19
C12983 VDD110 a_43993_n13477# 0.165f
C12984 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT 0.00187f
C12985 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN 3.46e-19
C12986 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 a_25535_354# 2.79e-20
C12987 RST a_36103_n10028# 0.00218f
C12988 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_54537_n6818# 0.00378f
C12989 CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 a_55067_297# 0.019f
C12990 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 1.16f
C12991 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.0995f
C12992 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 a_34896_n15539# 0.00119f
C12993 CLK_div_90_mag_0.CLK_div_10_mag_0.CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.235f
C12994 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 a_48422_n2199# 0.0036f
C12995 Vdiv100 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 0.00387f
C12996 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 a_50868_n16724# 0.0102f
C12997 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K a_22121_11196# 0.0811f
C12998 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB a_22559_n7106# 3.33e-19
C12999 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.235f
C13000 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 a_26052_n15491# 0.0697f
C13001 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN 0.111f
C13002 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB a_53221_2768# 0.00964f
C13003 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.0725f
C13004 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C13005 a_31128_n7028# CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 0.069f
C13006 RST a_45000_9057# 0.0014f
C13007 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 a_47723_574# 0.0105f
C13008 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 a_52139_n18696# 4.52e-20
C13009 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 3.6e-21
C13010 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.IN1 a_23139_n287# 0.0697f
C13011 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 0.0631f
C13012 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 0.109f
C13013 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_53168_n2243# 0.0731f
C13014 a_44315_n5176# CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0203f
C13015 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 a_49794_1671# 0.00118f
C13016 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT 0.103f
C13017 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.121f
C13018 VDD VDD90 0.356f
C13019 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_34308_n17626# 0.0733f
C13020 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.321f
C13021 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.0275f
C13022 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB 0.28f
C13023 a_49945_n6865# CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 2.99e-19
C13024 a_50768_2768# a_50928_2768# 0.0504f
C13025 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT 1.2e-19
C13026 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 4.53e-20
C13027 CLK_div_96_mag_0.JK_FF_mag_2.Q a_28583_n1899# 0.0101f
C13028 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K a_31445_n18723# 1.75e-19
C13029 VDD96 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT 0.995f
C13030 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN 0.0766f
C13031 CLK CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 9.71e-20
C13032 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 6.61e-20
C13033 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 5.36e-20
C13034 RST a_23948_n18723# 2.24e-19
C13035 CLK CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.271f
C13036 CLK_div_90_mag_0.CLK_div_10_mag_0.CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 9.71e-20
C13037 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB a_26196_5018# 0.00696f
C13038 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT 0.0286f
C13039 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 2.81e-20
C13040 VDD90 a_29241_7256# 6e-19
C13041 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 0.0595f
C13042 Vdiv110 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 0.00992f
C13043 a_31571_n16632# CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 5.54e-20
C13044 VDD110 a_49122_n18696# 3.56e-19
C13045 VDD100 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 1.07f
C13046 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 5.53e-19
C13047 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 1.14e-19
C13048 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00279f
C13049 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT 7.17e-19
C13050 VDD99 a_22551_n16006# 3.14e-19
C13051 VDD90 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K 0.497f
C13052 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 a_51005_n17599# 0.0102f
C13053 VDD93 a_36042_6265# 0.00175f
C13054 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 a_25420_n13385# 0.015f
C13055 CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 a_30760_n20290# 8.64e-19
C13056 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_26663_398# 0.011f
C13057 Vdiv108 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0212f
C13058 RST a_53785_2768# 0.00186f
C13059 RST a_26368_n2996# 0.0021f
C13060 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_54621_10154# 1.46e-19
C13061 CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_99_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 3.34e-19
C13062 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT a_48635_2768# 1.17e-20
C13063 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_4.IN2 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 0.321f
C13064 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 1.33e-19
C13065 RST a_53469_n15631# 7.84e-19
C13066 VDD99 a_24512_n18723# 3.14e-19
C13067 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT a_28580_n8735# 0.0202f
C13068 RST a_54027_n16728# 0.00199f
C13069 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB 0.414f
C13070 CLK_div_105_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_54414_6284# 5.94e-20
C13071 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 a_36588_n15495# 0.00372f
C13072 a_45927_6284# CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 4.52e-20
C13073 RST a_55020_n2199# 9.66e-19
C13074 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C13075 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 5.98e-20
C13076 CLK_div_108_new_mag_0.JK_FF_mag_0.QB a_53813_n6862# 0.00695f
C13077 dec3x8_ibr_mag_0.and_3_ibr_0.nand3_mag_ibr_0.OUT a_37328_6821# 3.58e-20
C13078 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB 0.00209f
C13079 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 9.08e-19
C13080 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C13081 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.198f
C13082 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_44069_5143# 0.0202f
C13083 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT Vdiv110 0.00836f
C13084 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 0.0635f
C13085 a_50103_5143# a_50263_5143# 0.0504f
C13086 a_26636_n8734# CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 4.52e-20
C13087 VDD100 a_53945_2768# 0.00123f
C13088 RST a_44888_1671# 0.0014f
C13089 VDD90 a_23025_6159# 3.14e-19
C13090 CLK a_22565_n6009# 0.00133f
C13091 CLK a_50103_5143# 0.00111f
C13092 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 a_24337_n6010# 0.0157f
C13093 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 a_48258_n10160# 1.27e-20
C13094 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB a_32009_n18723# 1.41e-20
C13095 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT 1.39e-19
C13096 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 a_33019_n16588# 0.0036f
C13097 RST CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.0152f
C13098 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 1.3f
C13099 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K a_47036_n15629# 0.00472f
C13100 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB 0.0838f
C13101 VDD110 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT 0.642f
C13102 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.OUT a_29871_n1855# 4.52e-20
C13103 CLK_div_108_new_mag_0.JK_FF_mag_1.QB CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 2.4e-20
C13104 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 a_35032_n17626# 2.58e-20
C13105 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 a_36588_n15495# 0.069f
C13106 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 0.00948f
C13107 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB a_24944_n8778# 1.07e-20
C13108 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0948f
C13109 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00254f
C13110 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0635f
C13111 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I1 a_37436_n1822# 0.00372f
C13112 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT 0.00481f
C13113 CLK a_54504_n10161# 0.00164f
C13114 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK a_50232_n7685# 3.27e-19
C13115 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00183f
C13116 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 4.75f
C13117 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 a_37436_880# 0.069f
C13118 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0622f
C13119 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_42083_n15712# 3.17e-19
C13120 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT 0.1f
C13121 a_51647_n10161# m3_20882_n11188# 0.00102f
C13122 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 7.24e-19
C13123 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 a_30209_7256# 0.0084f
C13124 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K 0.23f
C13125 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 a_25806_n17626# 5.98e-19
C13126 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT a_28335_6115# 0.0203f
C13127 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_27144_10099# 0.0203f
C13128 a_32015_n17626# a_32175_n17626# 0.0504f
C13129 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 6.26e-20
C13130 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 0.0295f
C13131 VDD108 a_51205_n7921# 5.92e-19
C13132 a_54504_n10161# a_54664_n10161# 0.0504f
C13133 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.00388f
C13134 RST CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 0.0196f
C13135 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK a_44413_n18696# 0.00939f
C13136 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 a_45618_2768# 0.00335f
C13137 VDD96 dec3x8_ibr_mag_0.and_3_ibr_1.nand3_mag_ibr_0.OUT 0.145f
C13138 Vdiv100 a_36873_280# 0.00152f
C13139 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0995f
C13140 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT 0.1f
C13141 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.00531f
C13142 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0377f
C13143 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_53785_2768# 8.64e-19
C13144 a_37168_6821# a_37328_6821# 0.0504f
C13145 VDD99 CLK_div_96_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.00271f
C13146 CLK_div_100_mag_0.CLK_div_10_mag_1.CLK CLK_div_100_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 0.0267f
C13147 VDD90 a_32640_6159# 3.14e-19
C13148 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 3.81e-19
C13149 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 0.273f
C13150 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT a_48148_n17599# 2.88e-20
C13151 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT 2.11e-20
C13152 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 a_38294_6265# 5.51e-19
C13153 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 1.53e-19
C13154 VDD105 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.442f
C13155 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB 2.59e-21
C13156 Vdiv110 mux_8x1_ibr_0.mux_2x1_ibr_0.I0 2.09e-19
C13157 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_53939_1671# 0.0202f
C13158 CLK a_44625_n15583# 3.8e-19
C13159 VDD dec3x8_ibr_mag_0.and_3_ibr_7.nand3_mag_ibr_0.OUT 0.671f
C13160 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.995f
C13161 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.338f
C13162 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 0.00488f
C13163 CLK a_47030_n16726# 0.00117f
C13164 RST a_46105_n18696# 6.14e-19
C13165 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT CLK_div_100_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.0654f
C13166 CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT 0.00132f
C13167 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT Vdiv93 3.84e-20
C13168 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.199f
C13169 VDD96 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 1.28f
C13170 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 a_49794_1671# 9.26e-19
C13171 CLK CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT 1.89e-21
C13172 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 a_26189_n6010# 0.006f
C13173 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C13174 VDD100 a_52839_n5# 3.14e-19
C13175 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_54751_n16684# 0.00859f
C13176 CLK_div_105_mag_0.CLK_div_10_mag_1.CLK CLK_div_105_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 0.0267f
C13177 CLK_div_108_new_mag_0.JK_FF_mag_1.Q a_53089_n6862# 0.00174f
C13178 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB a_44793_5143# 0.00695f
C13179 CLK a_31661_10099# 9.45e-19
C13180 CLK CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT 0.263f
C13181 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 0.209f
C13182 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN 0.00311f
C13183 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT CLK_div_96_mag_0.JK_FF_mag_3.Q 7.13e-20
C13184 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_51393_n6821# 0.0036f
C13185 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 a_48783_n13424# 0.0121f
C13186 mux_8x1_ibr_0.mux_2x1_ibr_0.I0 a_39124_280# 0.00293f
C13187 CLK_div_100_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN a_43559_n120# 5.39e-20
C13188 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.739f
C13189 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 a_51961_6284# 0.069f
C13190 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_33334_n18723# 4.52e-20
C13191 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.0854f
C13192 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.314f
C13193 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 a_53280_5143# 1.86e-20
C13194 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_54414_6284# 0.011f
C13195 VDD108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.397f
C13196 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_22455_5018# 0.0731f
C13197 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K 0.0823f
C13198 RST CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 0.301f
C13199 Vdiv110 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 3.1e-22
C13200 CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 a_54456_n2199# 0.00859f
C13201 RST CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 0.138f
C13202 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_108_new_mag_0.JK_FF_mag_1.Q 0.00335f
C13203 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K 4.04e-19
C13204 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 a_30164_n7017# 0.00347f
C13205 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_28552_354# 0.00119f
C13206 RST a_23748_n9840# 9.7e-19
C13207 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 a_22405_n6009# 8.64e-19
C13208 CLK_div_96_mag_0.JK_FF_mag_3.QB a_28743_n1899# 0.00392f
C13209 a_43757_n6273# CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 3.49e-20
C13210 VDD99 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.391f
C13211 a_29213_n7028# CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.069f
C13212 a_45075_n9063# a_45235_n9063# 0.0504f
C13213 RST CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.313f
C13214 CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_90_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.124f
C13215 VDD99 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 1.16f
C13216 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 1.16f
C13217 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT a_53129_n19793# 0.00138f
C13218 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT 0.053f
C13219 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00356f
C13220 Vdiv105 Vdiv90 0.00306f
C13221 m3_20882_n11188# VSS 12.8f $ **FLOATING
C13222 m1_42708_4265# VSS 0.371f $ **FLOATING
C13223 a_55357_n20487# VSS 0.0371f
C13224 a_55197_n20487# VSS 0.038f
C13225 CLK_div_110_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 VSS 0.337f
C13226 CLK_div_110_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS 0.669f
C13227 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT VSS 0.706f
C13228 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VSS 0.435f
C13229 a_53129_n19793# VSS 0.0679f
C13230 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT VSS 0.821f
C13231 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VSS 0.438f
C13232 a_52161_n19793# VSS 0.0679f
C13233 a_30760_n20290# VSS 0.0247f
C13234 CLK_div_110_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS 0.436f
C13235 a_51193_n19793# VSS 0.0676f
C13236 a_31733_n19822# VSS 0.0676f
C13237 CLK_div_99_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN VSS 0.435f
C13238 a_24391_n20290# VSS 0.0247f
C13239 CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 VSS 0.418f
C13240 CLK_div_99_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN VSS 0.6f
C13241 a_25364_n19822# VSS 0.0676f
C13242 CLK_div_99_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS 0.435f
C13243 CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 VSS 0.418f
C13244 CLK_div_99_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS 0.6f
C13245 a_55156_n18696# VSS 0.0676f
C13246 a_54592_n18696# VSS 0.0676f
C13247 a_54028_n18696# VSS 0.0676f
C13248 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.414f
C13249 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C13250 a_53464_n18696# VSS 0.0343f
C13251 a_53304_n18696# VSS 0.0881f
C13252 a_52139_n18696# VSS 0.0676f
C13253 a_51575_n18696# VSS 0.0676f
C13254 a_51011_n18696# VSS 0.0676f
C13255 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K VSS 0.633f
C13256 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VSS 0.414f
C13257 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VSS 0.509f
C13258 a_50447_n18696# VSS 0.0343f
C13259 a_50287_n18696# VSS 0.0881f
C13260 a_49122_n18696# VSS 0.0676f
C13261 a_48558_n18696# VSS 0.0676f
C13262 a_47994_n18696# VSS 0.0676f
C13263 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VSS 0.415f
C13264 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VSS 0.509f
C13265 a_47430_n18696# VSS 0.0343f
C13266 a_47270_n18696# VSS 0.0881f
C13267 a_46105_n18696# VSS 0.0676f
C13268 a_45541_n18696# VSS 0.0676f
C13269 a_44977_n18696# VSS 0.0676f
C13270 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.415f
C13271 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.509f
C13272 a_44413_n18696# VSS 0.0343f
C13273 a_44253_n18696# VSS 0.0881f
C13274 a_35186_n18723# VSS 0.0881f
C13275 a_35026_n18723# VSS 0.0343f
C13276 a_34462_n18723# VSS 0.0676f
C13277 a_33898_n18723# VSS 0.0676f
C13278 a_33334_n18723# VSS 0.0676f
C13279 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.509f
C13280 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.415f
C13281 a_32169_n18723# VSS 0.0881f
C13282 a_32009_n18723# VSS 0.0343f
C13283 a_31445_n18723# VSS 0.0676f
C13284 a_30881_n18723# VSS 0.0676f
C13285 a_30317_n18723# VSS 0.0676f
C13286 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C13287 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.415f
C13288 a_28817_n18723# VSS 0.0881f
C13289 a_28657_n18723# VSS 0.0343f
C13290 a_28093_n18723# VSS 0.0676f
C13291 a_27529_n18723# VSS 0.0676f
C13292 a_26965_n18723# VSS 0.0676f
C13293 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.509f
C13294 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.415f
C13295 a_25800_n18723# VSS 0.0881f
C13296 a_25640_n18723# VSS 0.0343f
C13297 a_25076_n18723# VSS 0.0676f
C13298 a_24512_n18723# VSS 0.0676f
C13299 a_23948_n18723# VSS 0.0676f
C13300 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C13301 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.415f
C13302 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K VSS 3.1f
C13303 a_55310_n17599# VSS 0.0675f
C13304 a_54746_n17599# VSS 0.0676f
C13305 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.415f
C13306 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.753f
C13307 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.807f
C13308 a_54182_n17599# VSS 0.0343f
C13309 a_54022_n17599# VSS 0.0881f
C13310 a_53458_n17599# VSS 0.0343f
C13311 a_53298_n17599# VSS 0.0881f
C13312 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB VSS 0.877f
C13313 a_52293_n17599# VSS 0.0675f
C13314 a_51729_n17599# VSS 0.0676f
C13315 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VSS 0.416f
C13316 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 VSS 0.693f
C13317 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VSS 0.808f
C13318 a_51165_n17599# VSS 0.0343f
C13319 a_51005_n17599# VSS 0.0881f
C13320 a_50441_n17599# VSS 0.0343f
C13321 a_50281_n17599# VSS 0.0881f
C13322 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB VSS 0.879f
C13323 a_49276_n17599# VSS 0.0675f
C13324 a_48712_n17599# VSS 0.0676f
C13325 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VSS 0.415f
C13326 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 VSS 0.696f
C13327 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VSS 0.809f
C13328 a_48148_n17599# VSS 0.0343f
C13329 a_47988_n17599# VSS 0.0881f
C13330 a_47424_n17599# VSS 0.0343f
C13331 a_47264_n17599# VSS 0.0881f
C13332 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB VSS 0.899f
C13333 a_46259_n17599# VSS 0.0675f
C13334 a_45695_n17599# VSS 0.0676f
C13335 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.416f
C13336 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.828f
C13337 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.81f
C13338 a_45131_n17599# VSS 0.0343f
C13339 a_44971_n17599# VSS 0.0881f
C13340 a_44407_n17599# VSS 0.0343f
C13341 a_44247_n17599# VSS 0.0881f
C13342 a_35192_n17626# VSS 0.0881f
C13343 a_35032_n17626# VSS 0.0343f
C13344 a_34468_n17626# VSS 0.0881f
C13345 a_34308_n17626# VSS 0.0343f
C13346 a_33744_n17626# VSS 0.0676f
C13347 a_33180_n17626# VSS 0.0675f
C13348 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB VSS 0.859f
C13349 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.811f
C13350 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.693f
C13351 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.418f
C13352 a_32175_n17626# VSS 0.0881f
C13353 a_32015_n17626# VSS 0.0343f
C13354 a_31451_n17626# VSS 0.0881f
C13355 a_31291_n17626# VSS 0.0343f
C13356 a_30727_n17626# VSS 0.0676f
C13357 a_30163_n17626# VSS 0.0675f
C13358 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K VSS 4.55f
C13359 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.811f
C13360 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.691f
C13361 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.417f
C13362 a_28823_n17626# VSS 0.0881f
C13363 a_28663_n17626# VSS 0.0343f
C13364 a_28099_n17626# VSS 0.0881f
C13365 a_27939_n17626# VSS 0.0343f
C13366 a_27375_n17626# VSS 0.0676f
C13367 a_26811_n17626# VSS 0.0675f
C13368 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB VSS 0.859f
C13369 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.81f
C13370 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.7f
C13371 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.417f
C13372 a_25806_n17626# VSS 0.0881f
C13373 a_25646_n17626# VSS 0.0343f
C13374 a_25082_n17626# VSS 0.0881f
C13375 a_24922_n17626# VSS 0.0343f
C13376 a_24358_n17626# VSS 0.0676f
C13377 a_23794_n17626# VSS 0.0675f
C13378 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K VSS 4.51f
C13379 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.81f
C13380 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.691f
C13381 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.417f
C13382 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.724f
C13383 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.519f
C13384 CLK_div_110_mag_0.CLK_div_10_mag_0.Q3 VSS 1.5f
C13385 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VSS 0.725f
C13386 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VSS 0.54f
C13387 CLK_div_110_mag_0.CLK_div_10_mag_0.Q2 VSS 2.23f
C13388 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VSS 0.726f
C13389 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VSS 0.539f
C13390 CLK_div_110_mag_0.CLK_div_10_mag_0.Q1 VSS 2.57f
C13391 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.724f
C13392 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.539f
C13393 CLK_div_110_mag_0.CLK_div_10_mag_0.Q0 VSS 3.35f
C13394 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.521f
C13395 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.726f
C13396 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0 VSS 2.54f
C13397 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.541f
C13398 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.727f
C13399 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.522f
C13400 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.726f
C13401 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0 VSS 2.3f
C13402 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.54f
C13403 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.726f
C13404 a_55315_n16684# VSS 0.0696f
C13405 a_54751_n16684# VSS 0.0698f
C13406 a_54187_n16728# VSS 0.0378f
C13407 a_54027_n16728# VSS 0.0916f
C13408 a_53463_n16728# VSS 0.0378f
C13409 a_53303_n16728# VSS 0.0917f
C13410 a_52156_n16680# VSS 0.069f
C13411 a_51592_n16680# VSS 0.0691f
C13412 a_51028_n16724# VSS 0.0367f
C13413 a_50868_n16724# VSS 0.0905f
C13414 a_50304_n16724# VSS 0.0368f
C13415 a_50144_n16724# VSS 0.0906f
C13416 a_49042_n16682# VSS 0.0693f
C13417 a_48478_n16682# VSS 0.0694f
C13418 a_47914_n16726# VSS 0.0372f
C13419 a_47754_n16726# VSS 0.0911f
C13420 a_47190_n16726# VSS 0.0373f
C13421 a_47030_n16726# VSS 0.0911f
C13422 a_45907_n16680# VSS 0.069f
C13423 a_45343_n16680# VSS 0.0691f
C13424 a_44779_n16724# VSS 0.0367f
C13425 a_44619_n16724# VSS 0.0905f
C13426 a_44055_n16724# VSS 0.0368f
C13427 a_43895_n16724# VSS 0.0906f
C13428 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 VSS 0.419f
C13429 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT VSS 0.551f
C13430 a_36742_n16592# VSS 0.0696f
C13431 a_36178_n16592# VSS 0.0698f
C13432 a_35614_n16636# VSS 0.0378f
C13433 a_35454_n16636# VSS 0.0916f
C13434 a_34890_n16636# VSS 0.0378f
C13435 a_34730_n16636# VSS 0.0917f
C13436 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 VSS 0.419f
C13437 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT VSS 0.549f
C13438 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.42f
C13439 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.551f
C13440 a_33583_n16588# VSS 0.069f
C13441 a_33019_n16588# VSS 0.0691f
C13442 a_32455_n16632# VSS 0.0367f
C13443 a_32295_n16632# VSS 0.0905f
C13444 a_31731_n16632# VSS 0.0368f
C13445 a_31571_n16632# VSS 0.0906f
C13446 a_30469_n16590# VSS 0.0693f
C13447 a_29905_n16590# VSS 0.0694f
C13448 a_29341_n16634# VSS 0.0372f
C13449 a_29181_n16634# VSS 0.0911f
C13450 a_28617_n16634# VSS 0.0373f
C13451 a_28457_n16634# VSS 0.0911f
C13452 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.418f
C13453 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.547f
C13454 a_41124_n16098# VSS 0.0716f
C13455 a_27334_n16588# VSS 0.069f
C13456 a_26770_n16588# VSS 0.0691f
C13457 a_26206_n16632# VSS 0.0367f
C13458 a_26046_n16632# VSS 0.0905f
C13459 a_25482_n16632# VSS 0.0368f
C13460 a_25322_n16632# VSS 0.0906f
C13461 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_4.IN2 VSS 0.421f
C13462 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_2.OUT VSS 0.553f
C13463 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_4.IN2 VSS 0.42f
C13464 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_2.OUT VSS 0.549f
C13465 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.42f
C13466 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.551f
C13467 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.419f
C13468 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.548f
C13469 a_55161_n15587# VSS 0.0744f
C13470 a_54597_n15587# VSS 0.0745f
C13471 a_54033_n15587# VSS 0.0744f
C13472 a_53469_n15631# VSS 0.047f
C13473 a_53309_n15631# VSS 0.101f
C13474 a_52002_n15583# VSS 0.0734f
C13475 a_51438_n15583# VSS 0.0735f
C13476 a_50874_n15583# VSS 0.0735f
C13477 a_50310_n15627# VSS 0.0449f
C13478 a_50150_n15627# VSS 0.0987f
C13479 a_48888_n15585# VSS 0.0739f
C13480 a_48324_n15585# VSS 0.074f
C13481 a_47760_n15585# VSS 0.0739f
C13482 a_47196_n15629# VSS 0.0459f
C13483 a_47036_n15629# VSS 0.0997f
C13484 a_45753_n15583# VSS 0.0737f
C13485 a_45189_n15583# VSS 0.0737f
C13486 a_44625_n15583# VSS 0.0737f
C13487 a_44061_n15627# VSS 0.0454f
C13488 a_43901_n15627# VSS 0.0992f
C13489 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 VSS 0.425f
C13490 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 VSS 0.906f
C13491 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 VSS 0.754f
C13492 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT VSS 0.83f
C13493 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT VSS 0.549f
C13494 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB VSS 0.954f
C13495 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN VSS 0.612f
C13496 a_42083_n15712# VSS 0.0247f
C13497 a_22551_n16006# VSS 0.0716f
C13498 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN VSS 0.45f
C13499 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 VSS 0.485f
C13500 a_36588_n15495# VSS 0.0744f
C13501 a_36024_n15495# VSS 0.0745f
C13502 a_35460_n15495# VSS 0.0744f
C13503 a_34896_n15539# VSS 0.047f
C13504 a_34736_n15539# VSS 0.101f
C13505 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 VSS 0.424f
C13506 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 VSS 0.86f
C13507 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 VSS 0.742f
C13508 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT VSS 0.827f
C13509 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT VSS 0.543f
C13510 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.424f
C13511 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.831f
C13512 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.743f
C13513 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.829f
C13514 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.546f
C13515 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB VSS 0.912f
C13516 a_33429_n15491# VSS 0.0734f
C13517 a_32865_n15491# VSS 0.0735f
C13518 a_32301_n15491# VSS 0.0735f
C13519 a_31737_n15535# VSS 0.0449f
C13520 a_31577_n15535# VSS 0.0987f
C13521 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.424f
C13522 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.844f
C13523 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.741f
C13524 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.826f
C13525 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.544f
C13526 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K VSS 1.92f
C13527 a_30315_n15493# VSS 0.0739f
C13528 a_29751_n15493# VSS 0.074f
C13529 a_29187_n15493# VSS 0.0739f
C13530 a_28623_n15537# VSS 0.0459f
C13531 a_28463_n15537# VSS 0.0997f
C13532 a_27180_n15491# VSS 0.0737f
C13533 a_26616_n15491# VSS 0.0737f
C13534 a_26052_n15491# VSS 0.0737f
C13535 a_25488_n15535# VSS 0.0454f
C13536 a_25328_n15535# VSS 0.0992f
C13537 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_1.IN2 VSS 0.425f
C13538 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand2_mag_3.IN1 VSS 0.908f
C13539 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.IN1 VSS 0.756f
C13540 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_1.OUT VSS 0.832f
C13541 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.nand3_mag_0.OUT VSS 0.549f
C13542 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.QB VSS 0.956f
C13543 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.GF_INV_MAG_1.IN VSS 0.612f
C13544 a_23510_n15620# VSS 0.0247f
C13545 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_0.GF_INV_MAG_0.IN VSS 0.45f
C13546 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN1 VSS 0.491f
C13547 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_1.IN2 VSS 0.424f
C13548 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand2_mag_3.IN1 VSS 0.86f
C13549 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.IN1 VSS 0.744f
C13550 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_1.OUT VSS 0.828f
C13551 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.nand3_mag_0.OUT VSS 0.543f
C13552 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.424f
C13553 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.832f
C13554 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.745f
C13555 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.83f
C13556 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.546f
C13557 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.QB VSS 0.912f
C13558 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.424f
C13559 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.844f
C13560 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.743f
C13561 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.827f
C13562 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.544f
C13563 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_0.K VSS 1.92f
C13564 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K VSS 3.1f
C13565 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 VSS 0.401f
C13566 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT VSS 0.585f
C13567 a_41284_n14596# VSS 0.0343f
C13568 a_41124_n14596# VSS 0.0881f
C13569 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN VSS 0.464f
C13570 a_42529_n14305# VSS 0.0676f
C13571 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K VSS 3.11f
C13572 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_0.IN2 VSS 0.403f
C13573 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_0.OUT VSS 0.585f
C13574 a_22711_n14504# VSS 0.0343f
C13575 a_22551_n14504# VSS 0.0881f
C13576 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_1.GF_INV_MAG_0.IN VSS 0.464f
C13577 a_23956_n14213# VSS 0.0676f
C13578 CLK_div_110_mag_0.CLK_div_10_mag_0.CLK VSS 11.2f
C13579 a_52385_n13362# VSS 0.0376f
C13580 a_52225_n13362# VSS 0.0391f
C13581 a_49488_n13383# VSS 0.0693f
C13582 a_48783_n13424# VSS 0.0362f
C13583 a_48623_n13424# VSS 0.0901f
C13584 a_41117_n13911# VSS 0.0678f
C13585 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT VSS 1.03f
C13586 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 VSS 0.555f
C13587 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K VSS 2.89f
C13588 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN VSS 0.676f
C13589 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT VSS 0.678f
C13590 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT VSS 1.93f
C13591 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN VSS 0.597f
C13592 a_43993_n13477# VSS 0.0247f
C13593 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K VSS 2.86f
C13594 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 VSS 18.6f
C13595 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 VSS 2.52f
C13596 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN VSS 0.589f
C13597 a_42521_n13474# VSS 0.0247f
C13598 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN VSS 0.453f
C13599 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q3 VSS 6.64f
C13600 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 VSS 0.532f
C13601 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN VSS 0.457f
C13602 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q1 VSS 6.62f
C13603 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS 0.701f
C13604 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q2 VSS 6.58f
C13605 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.Q0 VSS 5.91f
C13606 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 VSS 0.834f
C13607 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT VSS 0.741f
C13608 a_33812_n13270# VSS 0.0376f
C13609 a_33652_n13270# VSS 0.0391f
C13610 a_30915_n13291# VSS 0.0693f
C13611 a_30210_n13332# VSS 0.0362f
C13612 a_30050_n13332# VSS 0.0901f
C13613 a_22544_n13819# VSS 0.0678f
C13614 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.OUT VSS 1.03f
C13615 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nor_3_mag_0.IN3 VSS 0.555f
C13616 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_3.K VSS 2.9f
C13617 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_1.Inverter_delayed_mag_0.IN VSS 0.676f
C13618 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.GF_INV_MAG_1.OUT VSS 0.678f
C13619 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.OUT VSS 1.93f
C13620 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.GF_INV_MAG_1.IN VSS 0.597f
C13621 a_25420_n13385# VSS 0.0247f
C13622 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_2.K VSS 2.89f
C13623 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1 VSS 18.6f
C13624 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN2 VSS 2.52f
C13625 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.GF_INV_MAG_1.IN VSS 0.589f
C13626 a_23948_n13382# VSS 0.0247f
C13627 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_2.GF_INV_MAG_0.IN VSS 0.453f
C13628 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q3 VSS 6.53f
C13629 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_1.IN1 VSS 0.532f
C13630 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.GF_INV_MAG_0.IN VSS 0.457f
C13631 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q1 VSS 6.69f
C13632 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS 0.701f
C13633 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q2 VSS 6.76f
C13634 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.Q0 VSS 6.42f
C13635 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.and2_mag_3.IN1 VSS 0.834f
C13636 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.nand3_mag_1.OUT VSS 0.741f
C13637 a_54664_n10161# VSS 0.0881f
C13638 a_54504_n10161# VSS 0.0343f
C13639 a_53940_n10161# VSS 0.0881f
C13640 a_53780_n10161# VSS 0.0343f
C13641 a_53216_n10117# VSS 0.0676f
C13642 a_52652_n10117# VSS 0.0675f
C13643 a_51647_n10161# VSS 0.0881f
C13644 a_51487_n10161# VSS 0.0343f
C13645 a_50923_n10161# VSS 0.0881f
C13646 a_50763_n10161# VSS 0.0343f
C13647 a_50199_n10117# VSS 0.0676f
C13648 a_49635_n10117# VSS 0.0675f
C13649 a_48258_n10160# VSS 0.0881f
C13650 a_48098_n10160# VSS 0.0343f
C13651 a_47534_n10160# VSS 0.0881f
C13652 a_47374_n10160# VSS 0.0343f
C13653 a_46810_n10116# VSS 0.0676f
C13654 a_46246_n10116# VSS 0.0675f
C13655 a_45241_n10160# VSS 0.0881f
C13656 a_45081_n10160# VSS 0.0343f
C13657 a_44517_n10160# VSS 0.0881f
C13658 a_44357_n10160# VSS 0.0343f
C13659 a_43793_n10116# VSS 0.0676f
C13660 a_43229_n10116# VSS 0.0675f
C13661 a_40972_n9984# VSS 0.0675f
C13662 a_40408_n9984# VSS 0.0676f
C13663 a_39844_n10028# VSS 0.0343f
C13664 a_39684_n10028# VSS 0.0881f
C13665 a_39120_n10028# VSS 0.0343f
C13666 a_38960_n10028# VSS 0.0907f
C13667 a_37955_n9984# VSS 0.0675f
C13668 a_37391_n9984# VSS 0.0676f
C13669 a_36827_n10028# VSS 0.0343f
C13670 a_36667_n10028# VSS 0.0881f
C13671 a_36103_n10028# VSS 0.0343f
C13672 a_35943_n10028# VSS 0.0881f
C13673 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.521f
C13674 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.417f
C13675 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.541f
C13676 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.417f
C13677 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.521f
C13678 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.417f
C13679 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.541f
C13680 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.417f
C13681 a_29862_n9832# VSS 0.0675f
C13682 a_29298_n9832# VSS 0.0676f
C13683 a_28734_n9876# VSS 0.0343f
C13684 a_28574_n9876# VSS 0.0881f
C13685 a_28010_n9876# VSS 0.0343f
C13686 a_27850_n9876# VSS 0.0881f
C13687 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.417f
C13688 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.543f
C13689 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.417f
C13690 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.521f
C13691 a_26790_n9831# VSS 0.0675f
C13692 a_26226_n9831# VSS 0.0676f
C13693 a_25662_n9875# VSS 0.0343f
C13694 a_25502_n9875# VSS 0.0881f
C13695 a_24938_n9875# VSS 0.0343f
C13696 a_24778_n9875# VSS 0.0881f
C13697 a_23748_n9840# VSS 0.0686f
C13698 a_23184_n9840# VSS 0.0687f
C13699 a_22620_n9884# VSS 0.036f
C13700 a_22460_n9884# VSS 0.0898f
C13701 a_21896_n9884# VSS 0.036f
C13702 a_21736_n9884# VSS 0.0899f
C13703 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN VSS 0.677f
C13704 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN VSS 0.662f
C13705 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN VSS 0.662f
C13706 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN VSS 0.662f
C13707 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN VSS 0.666f
C13708 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN VSS 0.677f
C13709 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN VSS 0.762f
C13710 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 VSS 0.417f
C13711 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_2.OUT VSS 0.541f
C13712 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.417f
C13713 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.541f
C13714 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.419f
C13715 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.546f
C13716 a_54658_n9064# VSS 0.0881f
C13717 a_54498_n9064# VSS 0.0343f
C13718 a_53934_n9020# VSS 0.0676f
C13719 a_53370_n9020# VSS 0.0676f
C13720 a_52806_n9020# VSS 0.0676f
C13721 a_51641_n9064# VSS 0.0881f
C13722 a_51481_n9064# VSS 0.0343f
C13723 a_50917_n9020# VSS 0.0676f
C13724 a_50353_n9020# VSS 0.0676f
C13725 a_49789_n9020# VSS 0.0676f
C13726 a_48252_n9063# VSS 0.0881f
C13727 a_48092_n9063# VSS 0.0343f
C13728 a_47528_n9019# VSS 0.0676f
C13729 a_46964_n9019# VSS 0.0676f
C13730 a_46400_n9019# VSS 0.0676f
C13731 a_45235_n9063# VSS 0.0881f
C13732 a_45075_n9063# VSS 0.0343f
C13733 a_44511_n9019# VSS 0.0676f
C13734 a_43947_n9019# VSS 0.0676f
C13735 a_43383_n9019# VSS 0.0676f
C13736 a_40818_n8887# VSS 0.0676f
C13737 a_40254_n8887# VSS 0.0676f
C13738 a_39690_n8887# VSS 0.0676f
C13739 a_39126_n8931# VSS 0.0343f
C13740 a_38966_n8931# VSS 0.0884f
C13741 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.509f
C13742 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.811f
C13743 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.726f
C13744 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.693f
C13745 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.415f
C13746 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.QB VSS 0.859f
C13747 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C13748 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.811f
C13749 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.726f
C13750 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.692f
C13751 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.414f
C13752 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K VSS 4.41f
C13753 a_37801_n8887# VSS 0.0676f
C13754 a_37237_n8887# VSS 0.0676f
C13755 a_36673_n8887# VSS 0.0676f
C13756 a_36109_n8931# VSS 0.0343f
C13757 a_35949_n8931# VSS 0.0881f
C13758 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.508f
C13759 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.809f
C13760 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.724f
C13761 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.698f
C13762 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.415f
C13763 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB VSS 0.857f
C13764 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C13765 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.811f
C13766 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.726f
C13767 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.692f
C13768 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.415f
C13769 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K VSS 4.19f
C13770 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN VSS 0.707f
C13771 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN VSS 0.698f
C13772 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN VSS 0.698f
C13773 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN VSS 0.708f
C13774 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN VSS 0.681f
C13775 a_29708_n8735# VSS 0.0676f
C13776 a_29144_n8735# VSS 0.0676f
C13777 a_28580_n8735# VSS 0.0676f
C13778 a_28016_n8779# VSS 0.0343f
C13779 a_27856_n8779# VSS 0.0881f
C13780 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN VSS 0.761f
C13781 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN VSS 1.68f
C13782 CLK_div_93_mag_0.CLK_div_31_mag_0.Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN VSS 0.703f
C13783 a_26636_n8734# VSS 0.0676f
C13784 a_26072_n8734# VSS 0.0676f
C13785 a_25508_n8734# VSS 0.0676f
C13786 a_24944_n8778# VSS 0.0343f
C13787 a_24784_n8778# VSS 0.0881f
C13788 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.415f
C13789 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.692f
C13790 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.726f
C13791 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.811f
C13792 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C13793 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.415f
C13794 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.695f
C13795 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.726f
C13796 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.81f
C13797 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.509f
C13798 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB VSS 0.859f
C13799 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K VSS 4.55f
C13800 a_23594_n8743# VSS 0.0676f
C13801 a_23030_n8743# VSS 0.0676f
C13802 a_22466_n8743# VSS 0.0676f
C13803 a_21902_n8787# VSS 0.0343f
C13804 a_21742_n8787# VSS 0.0881f
C13805 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 VSS 0.413f
C13806 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 VSS 0.706f
C13807 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 VSS 0.724f
C13808 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_1.OUT VSS 0.809f
C13809 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.nand3_mag_0.OUT VSS 0.507f
C13810 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_4.QB VSS 0.929f
C13811 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.412f
C13812 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.691f
C13813 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.724f
C13814 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.809f
C13815 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.507f
C13816 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_1.QB VSS 0.886f
C13817 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.413f
C13818 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.739f
C13819 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.724f
C13820 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.814f
C13821 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.507f
C13822 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB VSS 1.61f
C13823 a_51205_n7921# VSS 0.0676f
C13824 a_50232_n7685# VSS 0.0247f
C13825 a_48023_n7840# VSS 0.0247f
C13826 a_44799_n7920# VSS 0.0676f
C13827 CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN VSS 0.598f
C13828 CLK_div_108_new_mag_0.CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN VSS 0.434f
C13829 CLK_div_108_new_mag_0.CLK_div_3_mag_2.or_2_mag_0.IN2 VSS 0.419f
C13830 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0 VSS 2.65f
C13831 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS 0.597f
C13832 CLK_div_108_new_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 VSS 0.416f
C13833 CLK_div_108_new_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS 0.433f
C13834 a_47050_n7372# VSS 0.0676f
C13835 a_43826_n7684# VSS 0.0247f
C13836 a_39402_n7788# VSS 0.0676f
C13837 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN VSS 0.601f
C13838 CLK_div_108_new_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN VSS 0.433f
C13839 CLK_div_108_new_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 VSS 0.416f
C13840 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0 VSS 2.73f
C13841 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS 0.601f
C13842 a_40375_n7552# VSS 0.0247f
C13843 CLK_div_93_mag_0.CLK_div_3_mag_0.Q0 VSS 1.7f
C13844 CLK_div_93_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 VSS 0.418f
C13845 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS 0.602f
C13846 a_32750_n7675# VSS 0.0247f
C13847 CLK_div_93_mag_0.CLK_div_31_mag_0.or_2_mag_0.IN1 VSS 1.34f
C13848 CLK_div_93_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS 0.435f
C13849 CLK_div_93_mag_0.CLK_div_3_mag_0.Q1 VSS 1.76f
C13850 CLK_div_93_mag_0.CLK_div_3_mag_0.CLK VSS 3.48f
C13851 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.GF_INV_MAG_0.IN VSS 0.413f
C13852 a_55101_n6818# VSS 0.0729f
C13853 a_54537_n6818# VSS 0.073f
C13854 a_53973_n6862# VSS 0.0439f
C13855 a_53813_n6862# VSS 0.0977f
C13856 a_53249_n6862# VSS 0.0439f
C13857 a_53089_n6862# VSS 0.0978f
C13858 a_51957_n6821# VSS 0.0736f
C13859 a_51393_n6821# VSS 0.0737f
C13860 a_50829_n6865# VSS 0.0454f
C13861 a_50669_n6865# VSS 0.0992f
C13862 a_50105_n6865# VSS 0.0454f
C13863 a_49945_n6865# VSS 0.0992f
C13864 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VSS 0.446f
C13865 a_31128_n7028# VSS 0.073f
C13866 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 VSS 0.4f
C13867 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VSS 0.451f
C13868 a_30164_n7017# VSS 0.0757f
C13869 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 VSS 0.397f
C13870 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VSS 0.443f
C13871 a_29213_n7028# VSS 0.073f
C13872 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 VSS 0.393f
C13873 CLK_div_93_mag_0.CLK_div_31_mag_0.nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS 0.445f
C13874 a_28267_n7033# VSS 0.072f
C13875 a_26343_n7107# VSS 0.0881f
C13876 a_26183_n7107# VSS 0.0343f
C13877 a_25619_n7107# VSS 0.0676f
C13878 a_25055_n7107# VSS 0.0676f
C13879 a_24491_n7107# VSS 0.0676f
C13880 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VSS 0.507f
C13881 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VSS 0.412f
C13882 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4 VSS 3.96f
C13883 a_23283_n7106# VSS 0.0881f
C13884 a_23123_n7106# VSS 0.0343f
C13885 a_22559_n7106# VSS 0.0676f
C13886 a_21995_n7106# VSS 0.0676f
C13887 a_21431_n7106# VSS 0.0676f
C13888 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VSS 0.506f
C13889 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VSS 0.413f
C13890 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.423f
C13891 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.57f
C13892 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.424f
C13893 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.57f
C13894 a_48466_n6273# VSS 0.0676f
C13895 a_47902_n6273# VSS 0.0676f
C13896 a_47338_n6273# VSS 0.0676f
C13897 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.415f
C13898 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C13899 a_46774_n6273# VSS 0.0343f
C13900 a_46614_n6273# VSS 0.0881f
C13901 a_45449_n6273# VSS 0.0676f
C13902 a_44885_n6273# VSS 0.0676f
C13903 a_44321_n6273# VSS 0.0676f
C13904 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.415f
C13905 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.508f
C13906 a_43757_n6273# VSS 0.0343f
C13907 a_43597_n6273# VSS 0.0881f
C13908 a_31129_n6271# VSS 0.073f
C13909 a_30165_n6282# VSS 0.0757f
C13910 a_29214_n6271# VSS 0.073f
C13911 a_54947_n5721# VSS 0.0676f
C13912 a_54383_n5721# VSS 0.0676f
C13913 a_53819_n5721# VSS 0.0676f
C13914 a_53255_n5765# VSS 0.0343f
C13915 a_53095_n5765# VSS 0.0881f
C13916 a_51803_n5724# VSS 0.0676f
C13917 a_51239_n5724# VSS 0.0676f
C13918 a_50675_n5724# VSS 0.0676f
C13919 a_50111_n5768# VSS 0.0343f
C13920 a_49951_n5768# VSS 0.0881f
C13921 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.VOUT VSS 2.77f
C13922 a_28268_n6266# VSS 0.0717f
C13923 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VSS 0.465f
C13924 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_3.IN2 VSS 0.4f
C13925 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VSS 0.451f
C13926 CLK_div_93_mag_0.CLK_div_31_mag_0.Q2 VSS 4.42f
C13927 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_2.IN2 VSS 0.398f
C13928 a_26349_n6010# VSS 0.0881f
C13929 a_26189_n6010# VSS 0.0343f
C13930 a_25625_n6010# VSS 0.0881f
C13931 a_25465_n6010# VSS 0.0343f
C13932 a_24901_n6010# VSS 0.0676f
C13933 a_24337_n6010# VSS 0.0675f
C13934 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.QB VSS 0.885f
C13935 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VSS 0.807f
C13936 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 VSS 0.699f
C13937 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VSS 0.416f
C13938 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VSS 0.445f
C13939 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3 VSS 6.07f
C13940 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_1.IN2 VSS 0.395f
C13941 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VSS 0.537f
C13942 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VSS 0.723f
C13943 a_23289_n6009# VSS 0.0881f
C13944 a_23129_n6009# VSS 0.0343f
C13945 a_22565_n6009# VSS 0.0881f
C13946 a_22405_n6009# VSS 0.0343f
C13947 a_21841_n6009# VSS 0.0676f
C13948 a_21277_n6009# VSS 0.0675f
C13949 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.QB VSS 0.923f
C13950 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VSS 0.807f
C13951 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 VSS 0.716f
C13952 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VSS 0.416f
C13953 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VSS 0.54f
C13954 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VSS 0.723f
C13955 CLK_div_93_mag_0.CLK_div_31_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS 0.448f
C13956 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1 VSS 7.25f
C13957 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0 VSS 3.73f
C13958 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.415f
C13959 CLK_div_108_new_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.829f
C13960 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.725f
C13961 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.84f
C13962 CLK_div_108_new_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C13963 CLK_div_108_new_mag_0.JK_FF_mag_0.QB VSS 0.873f
C13964 CLK_div_108_new_mag_0.JK_FF_mag_1.Q VSS 2.1f
C13965 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.415f
C13966 CLK_div_108_new_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.84f
C13967 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.723f
C13968 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.84f
C13969 CLK_div_108_new_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.509f
C13970 CLK_div_108_new_mag_0.JK_FF_mag_1.QB VSS 0.906f
C13971 CLK_div_108_new_mag_0.JK_FF_mag_1.CLK VSS 2.12f
C13972 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K VSS 4.34f
C13973 a_48620_n5176# VSS 0.0675f
C13974 a_48056_n5176# VSS 0.0676f
C13975 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.415f
C13976 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.69f
C13977 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.809f
C13978 a_47492_n5176# VSS 0.0343f
C13979 a_47332_n5176# VSS 0.0881f
C13980 a_46768_n5176# VSS 0.0343f
C13981 a_46608_n5176# VSS 0.0881f
C13982 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB VSS 0.857f
C13983 a_45603_n5176# VSS 0.0675f
C13984 a_45039_n5176# VSS 0.0676f
C13985 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.416f
C13986 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.697f
C13987 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.808f
C13988 a_44475_n5176# VSS 0.0343f
C13989 a_44315_n5176# VSS 0.0881f
C13990 a_43751_n5176# VSS 0.0343f
C13991 a_43591_n5176# VSS 0.0881f
C13992 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.724f
C13993 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.539f
C13994 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q0 VSS 1.64f
C13995 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.722f
C13996 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.519f
C13997 CLK_div_108_new_mag_0.CLK_div_3_mag_0.Q1 VSS 1.7f
C13998 a_30589_n2952# VSS 0.0765f
C13999 a_30025_n2952# VSS 0.0767f
C14000 a_29461_n2996# VSS 0.0522f
C14001 a_29301_n2996# VSS 0.106f
C14002 a_28737_n2996# VSS 0.0522f
C14003 a_28577_n2996# VSS 0.106f
C14004 a_27496_n2952# VSS 0.0765f
C14005 a_26932_n2952# VSS 0.0767f
C14006 a_26368_n2996# VSS 0.0522f
C14007 a_26208_n2996# VSS 0.106f
C14008 a_25644_n2996# VSS 0.0522f
C14009 a_25484_n2996# VSS 0.106f
C14010 a_24270_n2886# VSS 0.0675f
C14011 a_23706_n2886# VSS 0.0676f
C14012 a_23142_n2930# VSS 0.0343f
C14013 a_22982_n2930# VSS 0.0881f
C14014 a_22418_n2930# VSS 0.0343f
C14015 a_22258_n2930# VSS 0.0881f
C14016 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VSS 0.428f
C14017 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VSS 0.595f
C14018 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VSS 0.428f
C14019 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VSS 0.595f
C14020 a_55020_n2199# VSS 0.0675f
C14021 a_54456_n2199# VSS 0.0676f
C14022 a_53892_n2243# VSS 0.0343f
C14023 a_53732_n2243# VSS 0.0881f
C14024 a_53168_n2243# VSS 0.0343f
C14025 a_53008_n2243# VSS 0.0881f
C14026 a_52003_n2199# VSS 0.0675f
C14027 a_51439_n2199# VSS 0.0676f
C14028 a_50875_n2243# VSS 0.0343f
C14029 a_50715_n2243# VSS 0.0881f
C14030 a_50151_n2243# VSS 0.0343f
C14031 a_49991_n2243# VSS 0.0881f
C14032 a_48986_n2199# VSS 0.0675f
C14033 a_48422_n2199# VSS 0.0676f
C14034 a_47858_n2243# VSS 0.0343f
C14035 a_47698_n2243# VSS 0.0881f
C14036 a_47134_n2243# VSS 0.0343f
C14037 a_46974_n2243# VSS 0.0881f
C14038 a_45969_n2199# VSS 0.0675f
C14039 a_45405_n2199# VSS 0.0676f
C14040 a_44841_n2243# VSS 0.0343f
C14041 a_44681_n2243# VSS 0.0881f
C14042 a_44117_n2243# VSS 0.0343f
C14043 a_43957_n2243# VSS 0.0881f
C14044 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.416f
C14045 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.537f
C14046 a_37999_n1822# VSS 0.0676f
C14047 a_37436_n1822# VSS 0.0676f
C14048 a_36873_n1822# VSS 0.0676f
C14049 a_36310_n1822# VSS 0.0676f
C14050 a_35747_n1822# VSS 0.0676f
C14051 a_35184_n1822# VSS 0.0678f
C14052 a_30435_n1855# VSS 0.0676f
C14053 a_29871_n1855# VSS 0.0676f
C14054 a_29307_n1855# VSS 0.0676f
C14055 a_28743_n1899# VSS 0.0343f
C14056 a_28583_n1899# VSS 0.0881f
C14057 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_1.IN2 VSS 0.412f
C14058 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I1 VSS 0.416f
C14059 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_1.IN2 VSS 0.412f
C14060 Vdiv99 VSS 3.85f
C14061 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_1.IN2 VSS 0.43f
C14062 Vdiv93 VSS 9.87f
C14063 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.415f
C14064 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.519f
C14065 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VSS 0.415f
C14066 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VSS 0.539f
C14067 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VSS 0.415f
C14068 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VSS 0.539f
C14069 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.415f
C14070 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.539f
C14071 a_27342_n1855# VSS 0.0676f
C14072 a_26778_n1855# VSS 0.0676f
C14073 a_26214_n1855# VSS 0.0677f
C14074 a_25650_n1899# VSS 0.0349f
C14075 a_25490_n1899# VSS 0.0891f
C14076 a_24116_n1789# VSS 0.0685f
C14077 a_23552_n1789# VSS 0.068f
C14078 a_22988_n1789# VSS 0.0676f
C14079 a_22424_n1833# VSS 0.0343f
C14080 a_22264_n1833# VSS 0.0881f
C14081 a_54866_n1102# VSS 0.0676f
C14082 a_54302_n1102# VSS 0.0676f
C14083 a_53738_n1102# VSS 0.0676f
C14084 a_53174_n1146# VSS 0.0343f
C14085 a_53014_n1146# VSS 0.0881f
C14086 a_51849_n1102# VSS 0.0676f
C14087 a_51285_n1102# VSS 0.0676f
C14088 a_50721_n1102# VSS 0.0676f
C14089 a_50157_n1146# VSS 0.0343f
C14090 a_49997_n1146# VSS 0.0881f
C14091 a_48832_n1102# VSS 0.0676f
C14092 a_48268_n1102# VSS 0.0676f
C14093 a_47704_n1102# VSS 0.0676f
C14094 a_47140_n1146# VSS 0.0343f
C14095 a_46980_n1146# VSS 0.0881f
C14096 a_45815_n1102# VSS 0.0676f
C14097 a_45251_n1102# VSS 0.0676f
C14098 a_44687_n1102# VSS 0.0676f
C14099 a_44123_n1146# VSS 0.0343f
C14100 a_43963_n1146# VSS 0.0881f
C14101 a_37999_n1222# VSS 0.0676f
C14102 a_36873_n1222# VSS 0.0676f
C14103 a_35747_n1222# VSS 0.0676f
C14104 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VSS 0.414f
C14105 CLK_div_96_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 VSS 0.711f
C14106 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VSS 0.726f
C14107 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VSS 0.865f
C14108 CLK_div_96_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VSS 0.507f
C14109 CLK_div_96_mag_0.JK_FF_mag_3.QB VSS 0.907f
C14110 CLK_div_96_mag_0.JK_FF_mag_2.Q VSS 2.24f
C14111 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VSS 0.414f
C14112 CLK_div_96_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 VSS 0.774f
C14113 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VSS 0.727f
C14114 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VSS 0.866f
C14115 CLK_div_96_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VSS 0.514f
C14116 CLK_div_96_mag_0.JK_FF_mag_2.QB VSS 0.907f
C14117 CLK_div_96_mag_0.JK_FF_mag_0.Q VSS 2.39f
C14118 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.OUT VSS 0.597f
C14119 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.416f
C14120 CLK_div_96_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.742f
C14121 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.723f
C14122 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.805f
C14123 CLK_div_96_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.505f
C14124 CLK_div_96_mag_0.JK_FF_mag_0.QB VSS 0.894f
C14125 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.I0 VSS 0.765f
C14126 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_2.nand2_ibr_2.IN2 VSS 0.416f
C14127 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.OUT VSS 0.489f
C14128 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_1.nand2_ibr_2.IN2 VSS 0.417f
C14129 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.OUT VSS 0.429f
C14130 mux_8x1_ibr_0.mux_4x1_ibr_1.mux_2x1_ibr_0.nand2_ibr_2.IN2 VSS 0.436f
C14131 a_30398_n699# VSS 0.0675f
C14132 a_29834_n699# VSS 0.0676f
C14133 a_29270_n743# VSS 0.0343f
C14134 a_29110_n743# VSS 0.0881f
C14135 a_28546_n743# VSS 0.0343f
C14136 a_28386_n743# VSS 0.0881f
C14137 a_27381_n699# VSS 0.0675f
C14138 a_26817_n699# VSS 0.0676f
C14139 a_26253_n743# VSS 0.0344f
C14140 a_26093_n743# VSS 0.0883f
C14141 a_25529_n743# VSS 0.0352f
C14142 a_25369_n743# VSS 0.0893f
C14143 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.414f
C14144 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.753f
C14145 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.724f
C14146 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.807f
C14147 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C14148 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VSS 0.413f
C14149 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 VSS 0.692f
C14150 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VSS 0.724f
C14151 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VSS 0.808f
C14152 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VSS 0.509f
C14153 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB VSS 0.877f
C14154 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VSS 0.415f
C14155 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 VSS 0.695f
C14156 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VSS 0.724f
C14157 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VSS 0.806f
C14158 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VSS 0.506f
C14159 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB VSS 0.876f
C14160 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K VSS 3.14f
C14161 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.412f
C14162 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.767f
C14163 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.723f
C14164 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.806f
C14165 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.508f
C14166 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB VSS 0.888f
C14167 a_52839_n5# VSS 0.0679f
C14168 a_55067_297# VSS 0.0371f
C14169 a_54907_297# VSS 0.038f
C14170 a_51871_n5# VSS 0.0679f
C14171 a_50903_n5# VSS 0.0676f
C14172 CLK_div_100_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS 0.664f
C14173 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT VSS 0.701f
C14174 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K VSS 0.633f
C14175 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VSS 0.432f
C14176 CLK_div_100_mag_0.CLK_div_10_mag_0.Q0 VSS 3.36f
C14177 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VSS 0.438f
C14178 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS 0.433f
C14179 CLK_div_100_mag_0.CLK_div_10_mag_0.Q2 VSS 2.2f
C14180 CLK_div_100_mag_0.CLK_div_10_mag_0.Q1 VSS 2.59f
C14181 a_47723_574# VSS 0.0676f
C14182 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN VSS 0.433f
C14183 a_46755_574# VSS 0.0679f
C14184 a_43719_n120# VSS 0.038f
C14185 a_43559_n120# VSS 0.0371f
C14186 a_23863_n287# VSS 0.089f
C14187 a_23703_n287# VSS 0.0348f
C14188 a_23139_n287# VSS 0.0676f
C14189 a_22575_n287# VSS 0.0676f
C14190 a_22011_n287# VSS 0.0676f
C14191 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_0.OUT VSS 0.509f
C14192 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_1.IN2 VSS 0.41f
C14193 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.412f
C14194 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.537f
C14195 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.413f
C14196 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.524f
C14197 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN VSS 0.438f
C14198 a_45787_574# VSS 0.0679f
C14199 a_39124_280# VSS 0.0676f
C14200 mux_8x1_ibr_0.mux_2x1_ibr_0.I0 VSS 1.38f
C14201 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 VSS 0.422f
C14202 a_37999_280# VSS 0.0676f
C14203 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.IN2 VSS 0.414f
C14204 a_36873_280# VSS 0.0676f
C14205 Vdiv108 VSS 9.95f
C14206 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.IN2 VSS 0.417f
C14207 a_35747_280# VSS 0.0676f
C14208 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.IN2 VSS 0.436f
C14209 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN VSS 0.432f
C14210 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT VSS 0.701f
C14211 CLK_div_100_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS 0.664f
C14212 a_30244_398# VSS 0.0676f
C14213 a_29680_398# VSS 0.0676f
C14214 a_29116_398# VSS 0.0676f
C14215 a_28552_354# VSS 0.0343f
C14216 a_28392_354# VSS 0.0881f
C14217 CLK_div_100_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 VSS 0.335f
C14218 CLK_div_100_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT VSS 0.581f
C14219 Vdiv100 VSS 2.58f
C14220 CLK_div_100_mag_0.CLK_div_10_mag_0.Q3 VSS 1.78f
C14221 CLK_div_100_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT VSS 0.588f
C14222 CLK_div_100_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 VSS 0.335f
C14223 a_27227_398# VSS 0.0676f
C14224 a_26663_398# VSS 0.0676f
C14225 a_26099_398# VSS 0.0676f
C14226 a_25535_354# VSS 0.0343f
C14227 a_25375_354# VSS 0.0881f
C14228 a_39124_880# VSS 0.0676f
C14229 a_38561_880# VSS 0.0676f
C14230 a_37999_880# VSS 0.0676f
C14231 a_37436_880# VSS 0.0676f
C14232 a_36873_880# VSS 0.0676f
C14233 a_36310_880# VSS 0.0676f
C14234 a_35747_880# VSS 0.0676f
C14235 a_35184_880# VSS 0.0678f
C14236 a_23869_810# VSS 0.0949f
C14237 a_23709_810# VSS 0.041f
C14238 a_23145_810# VSS 0.0948f
C14239 a_22985_810# VSS 0.041f
C14240 a_22421_810# VSS 0.0715f
C14241 a_21857_810# VSS 0.0714f
C14242 CLK_div_96_mag_0.JK_FF_mag_5.QB VSS 0.894f
C14243 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.OUT VSS 0.826f
C14244 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_3.IN1 VSS 0.746f
C14245 CLK_div_96_mag_0.JK_FF_mag_5.nand2_mag_4.IN2 VSS 0.421f
C14246 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.415f
C14247 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.687f
C14248 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.721f
C14249 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.806f
C14250 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C14251 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.41f
C14252 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.699f
C14253 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.717f
C14254 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.802f
C14255 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.505f
C14256 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB VSS 0.852f
C14257 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K VSS 4.26f
C14258 CLK_div_96_mag_0.JK_FF_mag_5.Q VSS 3.04f
C14259 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_2.OUT VSS 0.56f
C14260 CLK_div_96_mag_0.JK_FF_mag_5.nand3_mag_1.IN1 VSS 0.722f
C14261 a_54663_1671# VSS 0.0881f
C14262 a_54503_1671# VSS 0.0343f
C14263 a_53939_1671# VSS 0.0676f
C14264 a_53375_1671# VSS 0.0676f
C14265 a_52811_1671# VSS 0.0676f
C14266 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.508f
C14267 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.412f
C14268 a_51646_1671# VSS 0.0881f
C14269 a_51486_1671# VSS 0.0343f
C14270 a_50922_1671# VSS 0.0676f
C14271 a_50358_1671# VSS 0.0676f
C14272 a_49794_1671# VSS 0.0676f
C14273 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT VSS 0.506f
C14274 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 VSS 0.415f
C14275 a_48629_1671# VSS 0.0881f
C14276 a_48469_1671# VSS 0.0343f
C14277 a_47905_1671# VSS 0.0676f
C14278 a_47341_1671# VSS 0.0676f
C14279 a_46777_1671# VSS 0.0676f
C14280 Vdiv VSS 7.83f
C14281 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I0 VSS 0.7f
C14282 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT VSS 0.623f
C14283 mux_8x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 VSS 0.412f
C14284 mux_8x1_ibr_0.mux_2x1_ibr_0.I1 VSS 0.416f
C14285 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_2.OUT VSS 0.488f
C14286 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.nand2_ibr_1.IN2 VSS 0.412f
C14287 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_2.I1 VSS 0.416f
C14288 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_2.OUT VSS 0.481f
C14289 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_1.nand2_ibr_1.IN2 VSS 0.412f
C14290 Vdiv110 VSS 15.3f
C14291 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_2.OUT VSS 0.429f
C14292 mux_8x1_ibr_0.mux_4x1_ibr_0.mux_2x1_ibr_0.nand2_ibr_1.IN2 VSS 0.432f
C14293 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT VSS 0.509f
C14294 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 VSS 0.413f
C14295 a_45612_1671# VSS 0.0881f
C14296 a_45452_1671# VSS 0.0343f
C14297 a_44888_1671# VSS 0.0676f
C14298 a_44324_1671# VSS 0.0676f
C14299 a_43760_1671# VSS 0.0676f
C14300 a_28828_1497# VSS 0.0676f
C14301 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C14302 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.414f
C14303 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K VSS 0.598f
C14304 Vdiv96 VSS 3.05f
C14305 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS 0.6f
C14306 a_29801_1733# VSS 0.0247f
C14307 CLK_div_96_mag_0.CLK_div_3_mag_0.Q0 VSS 1.73f
C14308 CLK_div_96_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 VSS 0.418f
C14309 CLK_div_96_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS 0.435f
C14310 CLK_div_96_mag_0.CLK_div_3_mag_0.Q1 VSS 1.72f
C14311 CLK_div_96_mag_0.JK_FF_mag_3.Q VSS 4.14f
C14312 a_26974_1919# VSS 0.0881f
C14313 a_26814_1919# VSS 0.0343f
C14314 a_26250_1919# VSS 0.0676f
C14315 a_25686_1919# VSS 0.0676f
C14316 a_25122_1919# VSS 0.0676f
C14317 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_0.OUT VSS 0.505f
C14318 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_1.IN2 VSS 0.41f
C14319 a_54669_2768# VSS 0.0881f
C14320 a_54509_2768# VSS 0.0343f
C14321 a_53945_2768# VSS 0.0881f
C14322 a_53785_2768# VSS 0.0343f
C14323 a_53221_2768# VSS 0.0676f
C14324 a_52657_2768# VSS 0.0675f
C14325 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB VSS 0.888f
C14326 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.806f
C14327 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.754f
C14328 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.415f
C14329 a_51652_2768# VSS 0.0881f
C14330 a_51492_2768# VSS 0.0343f
C14331 a_50928_2768# VSS 0.0881f
C14332 a_50768_2768# VSS 0.0343f
C14333 a_50204_2768# VSS 0.0676f
C14334 a_49640_2768# VSS 0.0675f
C14335 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB VSS 0.876f
C14336 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT VSS 0.806f
C14337 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 VSS 0.695f
C14338 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 VSS 0.415f
C14339 a_48635_2768# VSS 0.0881f
C14340 a_48475_2768# VSS 0.0343f
C14341 a_47911_2768# VSS 0.0881f
C14342 a_47751_2768# VSS 0.0343f
C14343 a_47187_2768# VSS 0.0676f
C14344 a_46623_2768# VSS 0.0675f
C14345 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB VSS 0.877f
C14346 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT VSS 0.808f
C14347 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 VSS 0.692f
C14348 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 VSS 0.415f
C14349 a_45618_2768# VSS 0.0881f
C14350 a_45458_2768# VSS 0.0343f
C14351 a_44894_2768# VSS 0.0881f
C14352 a_44734_2768# VSS 0.0343f
C14353 a_44170_2768# VSS 0.0676f
C14354 a_43606_2768# VSS 0.0675f
C14355 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K VSS 3.12f
C14356 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.807f
C14357 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.753f
C14358 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.415f
C14359 CLK_div_100_mag_0.CLK_div_10_mag_1.CLK VSS 1.62f
C14360 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.539f
C14361 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.723f
C14362 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT VSS 0.539f
C14363 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 VSS 0.724f
C14364 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1 VSS 2.99f
C14365 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT VSS 0.539f
C14366 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 VSS 0.724f
C14367 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0 VSS 3.52f
C14368 CLK_div_100_mag_0.CLK_div_10_mag_1.Q3 VSS 1.67f
C14369 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.519f
C14370 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.724f
C14371 a_26980_3016# VSS 0.0961f
C14372 a_26820_3016# VSS 0.0422f
C14373 a_26256_3016# VSS 0.096f
C14374 a_26096_3016# VSS 0.0422f
C14375 a_25532_3016# VSS 0.0721f
C14376 a_24968_3016# VSS 0.072f
C14377 CLK_div_96_mag_0.JK_FF_mag_4.QB VSS 0.899f
C14378 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.OUT VSS 0.83f
C14379 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_3.IN1 VSS 0.704f
C14380 CLK_div_96_mag_0.JK_FF_mag_4.nand2_mag_4.IN2 VSS 0.423f
C14381 CLK_div_96_mag_0.JK_FF_mag_4.Q VSS 3.6f
C14382 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_2.OUT VSS 0.564f
C14383 CLK_div_96_mag_0.JK_FF_mag_4.nand3_mag_1.IN1 VSS 0.722f
C14384 a_55132_5187# VSS 0.0675f
C14385 a_54568_5187# VSS 0.0676f
C14386 a_54004_5143# VSS 0.0343f
C14387 a_53844_5143# VSS 0.0881f
C14388 a_53280_5143# VSS 0.0343f
C14389 a_53120_5143# VSS 0.0881f
C14390 a_52115_5187# VSS 0.0675f
C14391 a_51551_5187# VSS 0.0676f
C14392 a_50987_5143# VSS 0.0343f
C14393 a_50827_5143# VSS 0.0881f
C14394 a_50263_5143# VSS 0.0343f
C14395 a_50103_5143# VSS 0.0881f
C14396 a_49098_5187# VSS 0.0675f
C14397 a_48534_5187# VSS 0.0676f
C14398 a_47970_5143# VSS 0.0343f
C14399 a_47810_5143# VSS 0.0881f
C14400 a_47246_5143# VSS 0.0343f
C14401 a_47086_5143# VSS 0.0881f
C14402 a_46081_5187# VSS 0.0675f
C14403 a_45517_5187# VSS 0.0676f
C14404 a_44953_5143# VSS 0.0343f
C14405 a_44793_5143# VSS 0.0881f
C14406 a_44229_5143# VSS 0.0343f
C14407 a_44069_5143# VSS 0.0881f
C14408 a_33358_5062# VSS 0.0675f
C14409 a_32794_5062# VSS 0.0676f
C14410 a_32230_5018# VSS 0.0343f
C14411 a_32070_5018# VSS 0.0881f
C14412 a_31506_5018# VSS 0.0343f
C14413 a_31346_5018# VSS 0.0881f
C14414 a_30341_5062# VSS 0.0675f
C14415 a_29777_5062# VSS 0.0676f
C14416 a_29213_5018# VSS 0.0343f
C14417 a_29053_5018# VSS 0.0881f
C14418 a_28489_5018# VSS 0.0343f
C14419 a_28329_5018# VSS 0.0881f
C14420 a_27324_5062# VSS 0.0675f
C14421 a_26760_5062# VSS 0.0676f
C14422 a_26196_5018# VSS 0.0343f
C14423 a_26036_5018# VSS 0.0881f
C14424 a_25472_5018# VSS 0.0343f
C14425 a_25312_5018# VSS 0.0881f
C14426 a_24307_5062# VSS 0.0675f
C14427 a_23743_5062# VSS 0.0676f
C14428 a_23179_5018# VSS 0.0343f
C14429 a_23019_5018# VSS 0.0881f
C14430 a_22455_5018# VSS 0.0343f
C14431 a_22295_5018# VSS 0.0881f
C14432 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.417f
C14433 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.521f
C14434 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VSS 0.416f
C14435 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VSS 0.541f
C14436 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VSS 0.416f
C14437 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VSS 0.541f
C14438 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.416f
C14439 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.541f
C14440 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.415f
C14441 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.519f
C14442 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_4.IN2 VSS 0.415f
C14443 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_2.OUT VSS 0.539f
C14444 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_4.IN2 VSS 0.415f
C14445 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_2.OUT VSS 0.539f
C14446 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.415f
C14447 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.541f
C14448 a_54978_6284# VSS 0.0676f
C14449 a_54414_6284# VSS 0.0676f
C14450 a_53850_6284# VSS 0.0676f
C14451 a_53286_6240# VSS 0.0343f
C14452 a_53126_6240# VSS 0.0881f
C14453 a_51961_6284# VSS 0.0676f
C14454 a_51397_6284# VSS 0.0676f
C14455 a_50833_6284# VSS 0.0676f
C14456 a_50269_6240# VSS 0.0343f
C14457 a_50109_6240# VSS 0.0881f
C14458 a_48944_6284# VSS 0.0676f
C14459 a_48380_6284# VSS 0.0676f
C14460 a_47816_6284# VSS 0.0676f
C14461 a_47252_6240# VSS 0.0343f
C14462 a_47092_6240# VSS 0.0881f
C14463 a_45927_6284# VSS 0.0676f
C14464 a_45363_6284# VSS 0.0676f
C14465 a_44799_6284# VSS 0.0676f
C14466 a_44235_6240# VSS 0.0343f
C14467 a_44075_6240# VSS 0.0881f
C14468 dec3x8_ibr_mag_0.and_3_ibr_7.nand3_mag_ibr_0.OUT VSS 0.506f
C14469 a_39580_6265# VSS 0.034f
C14470 a_39420_6265# VSS 0.0878f
C14471 dec3x8_ibr_mag_0.and_3_ibr_6.nand3_mag_ibr_0.OUT VSS 0.507f
C14472 a_38454_6265# VSS 0.034f
C14473 a_38294_6265# VSS 0.0878f
C14474 dec3x8_ibr_mag_0.and_3_ibr_5.nand3_mag_ibr_0.OUT VSS 0.506f
C14475 a_37328_6265# VSS 0.034f
C14476 a_37168_6265# VSS 0.0878f
C14477 dec3x8_ibr_mag_0.and_3_ibr_4.nand3_mag_ibr_0.OUT VSS 0.507f
C14478 a_36202_6265# VSS 0.034f
C14479 a_36042_6265# VSS 0.0878f
C14480 a_33204_6159# VSS 0.0676f
C14481 a_32640_6159# VSS 0.0676f
C14482 a_32076_6159# VSS 0.0676f
C14483 a_31512_6115# VSS 0.0343f
C14484 a_31352_6115# VSS 0.0881f
C14485 F0 VSS 13.9f
C14486 a_30187_6159# VSS 0.0676f
C14487 a_29623_6159# VSS 0.0676f
C14488 a_29059_6159# VSS 0.0676f
C14489 a_28495_6115# VSS 0.0343f
C14490 a_28335_6115# VSS 0.0881f
C14491 a_27170_6159# VSS 0.0676f
C14492 a_26606_6159# VSS 0.0676f
C14493 a_26042_6159# VSS 0.0676f
C14494 a_25478_6115# VSS 0.0343f
C14495 a_25318_6115# VSS 0.0881f
C14496 a_24153_6159# VSS 0.0676f
C14497 a_23589_6159# VSS 0.0676f
C14498 a_23025_6159# VSS 0.0676f
C14499 a_22461_6115# VSS 0.0343f
C14500 a_22301_6115# VSS 0.0881f
C14501 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.414f
C14502 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.755f
C14503 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.725f
C14504 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.808f
C14505 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C14506 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VSS 0.414f
C14507 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 VSS 0.693f
C14508 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VSS 0.726f
C14509 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VSS 0.809f
C14510 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VSS 0.509f
C14511 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB VSS 0.877f
C14512 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VSS 0.415f
C14513 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 VSS 0.696f
C14514 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VSS 0.725f
C14515 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VSS 0.81f
C14516 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VSS 0.509f
C14517 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB VSS 0.879f
C14518 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K VSS 3.14f
C14519 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.415f
C14520 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.91f
C14521 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.726f
C14522 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.811f
C14523 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.511f
C14524 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB VSS 0.899f
C14525 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.414f
C14526 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.753f
C14527 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.724f
C14528 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.807f
C14529 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C14530 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_1.IN2 VSS 0.413f
C14531 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand2_mag_3.IN1 VSS 0.692f
C14532 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.IN1 VSS 0.724f
C14533 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_1.OUT VSS 0.808f
C14534 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.nand3_mag_0.OUT VSS 0.509f
C14535 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_3.QB VSS 0.877f
C14536 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_1.IN2 VSS 0.415f
C14537 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand2_mag_3.IN1 VSS 0.695f
C14538 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.IN1 VSS 0.724f
C14539 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_1.OUT VSS 0.806f
C14540 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.nand3_mag_0.OUT VSS 0.506f
C14541 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.QB VSS 0.876f
C14542 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K VSS 3.14f
C14543 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.412f
C14544 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.76f
C14545 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.723f
C14546 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.806f
C14547 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.508f
C14548 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_1.QB VSS 0.888f
C14549 a_39580_6821# VSS 0.034f
C14550 a_39420_6821# VSS 0.0878f
C14551 a_38454_6821# VSS 0.034f
C14552 a_38294_6821# VSS 0.0878f
C14553 a_52951_7381# VSS 0.0679f
C14554 a_55179_7683# VSS 0.0371f
C14555 a_55019_7683# VSS 0.038f
C14556 a_51983_7381# VSS 0.0679f
C14557 a_51015_7381# VSS 0.0676f
C14558 CLK_div_105_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS 0.664f
C14559 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT VSS 0.701f
C14560 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K VSS 0.633f
C14561 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VSS 0.432f
C14562 CLK_div_105_mag_0.CLK_div_10_mag_0.Q0 VSS 3.36f
C14563 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VSS 0.438f
C14564 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS 0.433f
C14565 CLK_div_105_mag_0.CLK_div_10_mag_0.Q2 VSS 2.2f
C14566 CLK_div_105_mag_0.CLK_div_10_mag_0.Q1 VSS 2.59f
C14567 a_47835_7960# VSS 0.0676f
C14568 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.GF_INV_MAG_0.IN VSS 0.433f
C14569 a_46867_7960# VSS 0.0679f
C14570 a_43831_7266# VSS 0.038f
C14571 a_43671_7266# VSS 0.0371f
C14572 a_37328_6821# VSS 0.034f
C14573 a_37168_6821# VSS 0.0878f
C14574 dec3x8_ibr_mag_0.and_3_ibr_3.nand3_mag_ibr_0.OUT VSS 0.517f
C14575 a_36202_6821# VSS 0.034f
C14576 a_36042_6821# VSS 0.0878f
C14577 dec3x8_ibr_mag_0.and_3_ibr_2.nand3_mag_ibr_0.OUT VSS 0.501f
C14578 dec3x8_ibr_mag_0.and_3_ibr_1.nand3_mag_ibr_0.OUT VSS 0.501f
C14579 F1 VSS 8.07f
C14580 dec3x8_ibr_mag_0.and_3_ibr_0.nand3_mag_ibr_0.OUT VSS 0.501f
C14581 dec3x8_ibr_mag_0.and_3_ibr_3.IN1 VSS 1.49f
C14582 dec3x8_ibr_mag_0.and_3_ibr_6.IN3 VSS 1.9f
C14583 dec3x8_ibr_mag_0.and_3_ibr_5.IN3 VSS 1.92f
C14584 F2 VSS 8.63f
C14585 a_31177_7256# VSS 0.0679f
C14586 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_2.GF_INV_MAG_0.IN VSS 0.438f
C14587 a_45899_7960# VSS 0.0679f
C14588 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.GF_INV_MAG_0.IN VSS 0.432f
C14589 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_1.OUT VSS 0.701f
C14590 CLK_div_105_mag_0.CLK_div_10_mag_1.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS 0.664f
C14591 CLK_div_105_mag_0.CLK_div_10_mag_1.nor_3_mag_0.IN3 VSS 0.335f
C14592 CLK_div_105_mag_0.CLK_div_10_mag_1.and2_mag_0.OUT VSS 0.58f
C14593 Vdiv90 VSS 3.16f
C14594 a_33405_7558# VSS 0.0371f
C14595 a_33245_7558# VSS 0.038f
C14596 a_30209_7256# VSS 0.0679f
C14597 a_29241_7256# VSS 0.0676f
C14598 CLK_div_90_mag_0.CLK_div_10_mag_0.Buffer_delayed_mag_0.Inverter_delayed_mag_0.IN VSS 0.669f
C14599 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.OUT VSS 0.706f
C14600 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_0.K VSS 0.633f
C14601 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_1.GF_INV_MAG_0.IN VSS 0.435f
C14602 CLK_div_90_mag_0.CLK_div_10_mag_0.Q0 VSS 3.5f
C14603 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_2.GF_INV_MAG_0.IN VSS 0.438f
C14604 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS 0.435f
C14605 CLK_div_90_mag_0.CLK_div_10_mag_0.Q2 VSS 2.22f
C14606 CLK_div_90_mag_0.CLK_div_10_mag_0.Q1 VSS 2.63f
C14607 Vdiv105 VSS 8.67f
C14608 CLK_div_90_mag_0.CLK_div_10_mag_0.Q3 VSS 1.64f
C14609 CLK_div_90_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT VSS 0.737f
C14610 CLK_div_90_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 VSS 0.337f
C14611 CLK_div_105_mag_0.CLK_div_10_mag_0.Q3 VSS 1.92f
C14612 CLK_div_105_mag_0.CLK_div_10_mag_0.and2_mag_0.OUT VSS 0.599f
C14613 CLK_div_105_mag_0.CLK_div_10_mag_0.nor_3_mag_0.IN3 VSS 0.335f
C14614 a_54775_9057# VSS 0.0881f
C14615 a_54615_9057# VSS 0.0343f
C14616 a_54051_9057# VSS 0.0676f
C14617 a_53487_9057# VSS 0.0676f
C14618 a_52923_9057# VSS 0.0676f
C14619 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.508f
C14620 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.412f
C14621 a_51758_9057# VSS 0.0881f
C14622 a_51598_9057# VSS 0.0343f
C14623 a_51034_9057# VSS 0.0676f
C14624 a_50470_9057# VSS 0.0676f
C14625 a_49906_9057# VSS 0.0676f
C14626 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_0.OUT VSS 0.506f
C14627 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_1.IN2 VSS 0.415f
C14628 a_48741_9057# VSS 0.0881f
C14629 a_48581_9057# VSS 0.0343f
C14630 a_48017_9057# VSS 0.0676f
C14631 a_47453_9057# VSS 0.0676f
C14632 a_46889_9057# VSS 0.0676f
C14633 a_29087_8532# VSS 0.0247f
C14634 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_0.OUT VSS 0.509f
C14635 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_1.IN2 VSS 0.413f
C14636 a_45724_9057# VSS 0.0881f
C14637 a_45564_9057# VSS 0.0343f
C14638 a_45000_9057# VSS 0.0676f
C14639 a_44436_9057# VSS 0.0676f
C14640 a_43872_9057# VSS 0.0676f
C14641 a_30060_9000# VSS 0.0676f
C14642 CLK_div_90_mag_0.CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN VSS 0.434f
C14643 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C14644 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.414f
C14645 a_22718_8532# VSS 0.0259f
C14646 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.K VSS 0.598f
C14647 CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.IN2 VSS 0.416f
C14648 CLK_div_90_mag_0.CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN VSS 0.6f
C14649 a_23691_9000# VSS 0.0676f
C14650 CLK_div_90_mag_0.CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS 0.436f
C14651 CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.IN2 VSS 0.42f
C14652 CLK_div_90_mag_0.CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS 0.606f
C14653 CLK_div_90_mag_0.CLK_div_10_mag_0.CLK VSS 2.59f
C14654 a_54781_10154# VSS 0.0881f
C14655 a_54621_10154# VSS 0.0343f
C14656 a_54057_10154# VSS 0.0881f
C14657 a_53897_10154# VSS 0.0343f
C14658 a_53333_10154# VSS 0.0676f
C14659 a_52769_10154# VSS 0.0675f
C14660 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.QB VSS 0.888f
C14661 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.806f
C14662 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.757f
C14663 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.415f
C14664 a_51764_10154# VSS 0.0881f
C14665 a_51604_10154# VSS 0.0343f
C14666 a_51040_10154# VSS 0.0881f
C14667 a_50880_10154# VSS 0.0343f
C14668 a_50316_10154# VSS 0.0676f
C14669 a_49752_10154# VSS 0.0675f
C14670 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.QB VSS 0.876f
C14671 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.OUT VSS 0.806f
C14672 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_3.IN1 VSS 0.695f
C14673 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand2_mag_4.IN2 VSS 0.415f
C14674 a_48747_10154# VSS 0.0881f
C14675 a_48587_10154# VSS 0.0343f
C14676 a_48023_10154# VSS 0.0881f
C14677 a_47863_10154# VSS 0.0343f
C14678 a_47299_10154# VSS 0.0676f
C14679 a_46735_10154# VSS 0.0675f
C14680 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.QB VSS 0.877f
C14681 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.OUT VSS 0.808f
C14682 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_3.IN1 VSS 0.692f
C14683 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand2_mag_4.IN2 VSS 0.415f
C14684 a_45730_10154# VSS 0.0881f
C14685 a_45570_10154# VSS 0.0343f
C14686 a_45006_10154# VSS 0.0881f
C14687 a_44846_10154# VSS 0.0343f
C14688 a_44282_10154# VSS 0.0676f
C14689 a_43718_10154# VSS 0.0675f
C14690 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K VSS 3.12f
C14691 a_33513_10099# VSS 0.0881f
C14692 a_33353_10099# VSS 0.0343f
C14693 a_32789_10099# VSS 0.0676f
C14694 a_32225_10099# VSS 0.0676f
C14695 a_31661_10099# VSS 0.0676f
C14696 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.509f
C14697 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.415f
C14698 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.807f
C14699 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.753f
C14700 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.415f
C14701 a_30496_10099# VSS 0.0881f
C14702 a_30336_10099# VSS 0.0343f
C14703 a_29772_10099# VSS 0.0676f
C14704 a_29208_10099# VSS 0.0676f
C14705 a_28644_10099# VSS 0.0676f
C14706 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C14707 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.415f
C14708 a_27144_10099# VSS 0.0881f
C14709 a_26984_10099# VSS 0.0343f
C14710 a_26420_10099# VSS 0.0676f
C14711 a_25856_10099# VSS 0.0676f
C14712 a_25292_10099# VSS 0.0676f
C14713 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.509f
C14714 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.415f
C14715 a_24127_10099# VSS 0.0881f
C14716 a_23967_10099# VSS 0.0343f
C14717 a_23403_10099# VSS 0.0676f
C14718 a_22839_10099# VSS 0.0676f
C14719 a_22275_10099# VSS 0.0676f
C14720 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C14721 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.415f
C14722 CLK_div_105_mag_0.CLK_div_10_mag_1.CLK VSS 1.63f
C14723 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.539f
C14724 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.723f
C14725 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_2.OUT VSS 0.539f
C14726 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.nand3_mag_1.IN1 VSS 0.724f
C14727 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1 VSS 2.99f
C14728 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_2.OUT VSS 0.539f
C14729 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_3.nand3_mag_1.IN1 VSS 0.724f
C14730 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0 VSS 3.52f
C14731 CLK_div_105_mag_0.CLK_div_10_mag_1.Q3 VSS 1.79f
C14732 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.519f
C14733 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.724f
C14734 a_33519_11196# VSS 0.0881f
C14735 a_33359_11196# VSS 0.0343f
C14736 a_32795_11196# VSS 0.0881f
C14737 a_32635_11196# VSS 0.0343f
C14738 a_32071_11196# VSS 0.0676f
C14739 a_31507_11196# VSS 0.0675f
C14740 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.QB VSS 0.859f
C14741 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.81f
C14742 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.695f
C14743 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.417f
C14744 a_30502_11196# VSS 0.0881f
C14745 a_30342_11196# VSS 0.0343f
C14746 a_29778_11196# VSS 0.0881f
C14747 a_29618_11196# VSS 0.0343f
C14748 a_29054_11196# VSS 0.0676f
C14749 a_28490_11196# VSS 0.0675f
C14750 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K VSS 4.54f
C14751 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.81f
C14752 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.691f
C14753 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.416f
C14754 a_27150_11196# VSS 0.0881f
C14755 a_26990_11196# VSS 0.0343f
C14756 a_26426_11196# VSS 0.0881f
C14757 a_26266_11196# VSS 0.0343f
C14758 a_25702_11196# VSS 0.0676f
C14759 a_25138_11196# VSS 0.0675f
C14760 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.QB VSS 0.859f
C14761 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.81f
C14762 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.7f
C14763 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.417f
C14764 a_24133_11196# VSS 0.0881f
C14765 a_23973_11196# VSS 0.0343f
C14766 a_23409_11196# VSS 0.0881f
C14767 a_23249_11196# VSS 0.0343f
C14768 a_22685_11196# VSS 0.0676f
C14769 a_22121_11196# VSS 0.0675f
C14770 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K VSS 4.55f
C14771 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.81f
C14772 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.691f
C14773 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.416f
C14774 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.521f
C14775 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.725f
C14776 CLK VSS 96.2f
C14777 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0 VSS 2.64f
C14778 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.54f
C14779 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.725f
C14780 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.521f
C14781 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.725f
C14782 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0 VSS 2.77f
C14783 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.54f
C14784 RST VSS 96.7f
C14785 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.725f
C14786 VDD110 VSS 0.171p
C14787 VDD99 VSS 0.191p
C14788 VDD93 VSS 0.152p
C14789 VDD108 VSS 0.146p
C14790 VDD100 VSS 0.138p
C14791 VDD96 VSS 0.106p
C14792 VDD105 VSS 0.136p
C14793 VDD90 VSS 0.147p
C14794 VDD VSS 72.4f
C14795 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t3 VSS 0.0207f
C14796 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t5 VSS 0.0271f
C14797 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n0 VSS 0.0537f
C14798 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t4 VSS 0.0273f
C14799 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t2 VSS 0.0207f
C14800 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n1 VSS 0.0537f
C14801 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n2 VSS 0.675f
C14802 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n3 VSS 0.0327f
C14803 Vdiv90.t4 VSS 0.0116f
C14804 Vdiv90.t5 VSS 0.0146f
C14805 Vdiv90.n0 VSS 0.0345f
C14806 Vdiv90.n1 VSS 0.00688f
C14807 Vdiv90.n2 VSS 0.00422f
C14808 Vdiv90.n3 VSS 0.0022f
C14809 Vdiv90.n4 VSS 0.00309f
C14810 Vdiv90.n5 VSS 0.0887f
C14811 Vdiv90.t3 VSS 0.00295f
C14812 Vdiv90.n6 VSS 0.00295f
C14813 Vdiv90.n7 VSS 0.0141f
C14814 Vdiv90.n8 VSS 0.00674f
C14815 Vdiv90.n9 VSS 0.0714f
C14816 Vdiv90.n10 VSS 0.103f
C14817 Vdiv90.n11 VSS 0.549f
C14818 Vdiv90.n12 VSS 0.349f
C14819 Vdiv90.n13 VSS 0.0126f
C14820 Vdiv90.n14 VSS 9.94e-19
C14821 Vdiv90.n15 VSS 0.00597f
C14822 Vdiv90.n16 VSS 0.00365f
C14823 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n0 VSS 2.2f
C14824 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n1 VSS 0.159f
C14825 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t6 VSS 0.0515f
C14826 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t5 VSS 0.0808f
C14827 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n2 VSS 0.143f
C14828 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t8 VSS 0.0739f
C14829 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t7 VSS 0.0576f
C14830 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n3 VSS 0.147f
C14831 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t4 VSS 0.046f
C14832 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t3 VSS 0.0576f
C14833 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n4 VSS 0.148f
C14834 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n5 VSS 1.23f
C14835 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t0 VSS 0.0359f
C14836 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n6 VSS 0.0359f
C14837 CLK_div_108_new_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n7 VSS 0.0766f
C14838 F2.n0 VSS 0.116f
C14839 F2.n1 VSS 0.0117f
C14840 F2.t6 VSS 0.0237f
C14841 F2.t8 VSS 0.0185f
C14842 F2.n2 VSS 0.0471f
C14843 F2.n3 VSS 0.00659f
C14844 F2.n4 VSS 0.00332f
C14845 F2.n5 VSS 0.0296f
C14846 F2.n6 VSS 0.00885f
C14847 F2.n7 VSS 0.00494f
C14848 F2.n8 VSS 1.88e-19
C14849 F2.t11 VSS 0.0255f
C14850 F2.t9 VSS 0.0162f
C14851 F2.n9 VSS 0.0154f
C14852 F2.n10 VSS 0.0308f
C14853 F2.n11 VSS 3.77e-19
C14854 F2.n12 VSS 0.00245f
C14855 F2.n13 VSS 0.115f
C14856 F2.n14 VSS 0.00292f
C14857 F2.n15 VSS 0.00661f
C14858 F2.t7 VSS 0.0182f
C14859 F2.t5 VSS 0.024f
C14860 F2.n16 VSS 0.0469f
C14861 F2.n17 VSS 0.0123f
C14862 F2.n18 VSS 0.0217f
C14863 F2.n19 VSS 0.131f
C14864 F2.n20 VSS 0.165f
C14865 F2.n21 VSS 0.112f
C14866 F2.n22 VSS 2.16e-19
C14867 F2.t10 VSS 0.0163f
C14868 F2.n23 VSS 0.016f
C14869 F2.t12 VSS 0.0254f
C14870 F2.n24 VSS 0.0303f
C14871 F2.n25 VSS 6.48e-19
C14872 F2.n26 VSS 0.00302f
C14873 F2.n27 VSS 0.006f
C14874 F2.n28 VSS 0.00944f
C14875 F2.n29 VSS 0.212f
C14876 F2.t1 VSS 0.0196f
C14877 F2.n30 VSS 0.0198f
C14878 F2.t3 VSS 0.00319f
C14879 F2.n31 VSS 0.0121f
C14880 F2.n32 VSS 0.00695f
C14881 F2.n33 VSS 2.45e-19
C14882 F2.n34 VSS 0.138f
C14883 F2.t2 VSS 0.0147f
C14884 F2.t0 VSS 0.0185f
C14885 F2.n35 VSS 0.0437f
C14886 F2.n36 VSS 0.0229f
C14887 F2.n37 VSS 0.00448f
C14888 F2.n38 VSS 5.89e-19
C14889 F2.t4 VSS 0.00537f
C14890 F2.t13 VSS 0.0214f
C14891 F2.n39 VSS 0.0348f
C14892 F2.n40 VSS 8.93e-19
C14893 F2.n41 VSS 0.0847f
C14894 F2.n42 VSS 1.16f
C14895 F2.n43 VSS 2.81f
C14896 F1.n0 VSS 0.156f
C14897 F1.t17 VSS 0.00619f
C14898 F1.n1 VSS 0.0155f
C14899 F1.t16 VSS 0.0282f
C14900 F1.n2 VSS 0.0322f
C14901 F1.n3 VSS 7.45e-19
C14902 F1.n4 VSS 0.00164f
C14903 F1.n5 VSS 0.0132f
C14904 F1.n6 VSS 0.00858f
C14905 F1.t9 VSS 0.0219f
C14906 F1.n7 VSS 0.0193f
C14907 F1.t11 VSS 0.0341f
C14908 F1.n8 VSS 0.0418f
C14909 F1.n9 VSS 7.75e-19
C14910 F1.n10 VSS 0.00362f
C14911 F1.n11 VSS 0.125f
C14912 F1.n12 VSS 0.131f
C14913 F1.n13 VSS 7.51e-19
C14914 F1.t10 VSS 0.0342f
C14915 F1.t6 VSS 0.0225f
C14916 F1.n14 VSS 0.0604f
C14917 F1.n15 VSS 1.36e-19
C14918 F1.n16 VSS 0.00403f
C14919 F1.n17 VSS 0.00564f
C14920 F1.n18 VSS 0.00755f
C14921 F1.n19 VSS 0.238f
C14922 F1.t3 VSS 0.0225f
C14923 F1.t7 VSS 0.0342f
C14924 F1.n20 VSS 0.0604f
C14925 F1.n21 VSS 0.00236f
C14926 F1.n22 VSS 0.0968f
C14927 F1.n23 VSS 0.168f
C14928 F1.n24 VSS 0.00372f
C14929 F1.n25 VSS 0.00276f
C14930 F1.n26 VSS 7.53e-19
C14931 F1.n27 VSS 0.00301f
C14932 F1.t2 VSS 0.0215f
C14933 F1.n28 VSS 0.0198f
C14934 F1.t5 VSS 0.0341f
C14935 F1.n29 VSS 0.0417f
C14936 F1.n30 VSS 5.02e-19
C14937 F1.n31 VSS 8.78e-19
C14938 F1.n32 VSS 0.00905f
C14939 F1.n33 VSS 4.24e-19
C14940 F1.n34 VSS 0.00509f
C14941 F1.n35 VSS 0.00226f
C14942 F1.n36 VSS 0.0115f
C14943 F1.n37 VSS 0.00397f
C14944 F1.n38 VSS 0.0658f
C14945 F1.n39 VSS 0.639f
C14946 F1.n40 VSS 0.238f
C14947 F1.n41 VSS 0.0112f
C14948 F1.n42 VSS 0.134f
C14949 F1.n43 VSS 0.00805f
C14950 F1.t13 VSS 0.0196f
C14951 F1.t8 VSS 0.0246f
C14952 F1.n44 VSS 0.0582f
C14953 F1.n45 VSS 0.0211f
C14954 F1.n46 VSS 0.0137f
C14955 F1.n47 VSS 0.00597f
C14956 F1.t1 VSS 0.0285f
C14957 F1.t12 VSS 0.00716f
C14958 F1.n48 VSS 0.0464f
C14959 F1.n49 VSS 0.0159f
C14960 F1.t14 VSS 0.0196f
C14961 F1.t4 VSS 0.0246f
C14962 F1.n50 VSS 0.0582f
C14963 F1.n51 VSS 0.0211f
C14964 F1.n52 VSS 0.00827f
C14965 F1.n53 VSS 0.125f
C14966 F1.n54 VSS 0.118f
C14967 F1.n55 VSS 0.00597f
C14968 F1.n56 VSS 0.179f
C14969 F1.n57 VSS 0.18f
C14970 F1.t15 VSS 0.00716f
C14971 F1.t0 VSS 0.0285f
C14972 F1.n58 VSS 0.0464f
C14973 F1.n59 VSS 0.0159f
C14974 F1.n60 VSS 0.113f
C14975 F1.n61 VSS 1.33f
C14976 F1.n62 VSS 4.09f
C14977 Vdiv93.t3 VSS 0.00555f
C14978 Vdiv93.t2 VSS 0.0102f
C14979 Vdiv93.n0 VSS 0.0191f
C14980 Vdiv93.n1 VSS 0.0122f
C14981 Vdiv93.n2 VSS 0.00366f
C14982 Vdiv93.n3 VSS 0.0413f
C14983 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n0 VSS 0.511f
C14984 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n1 VSS 0.322f
C14985 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n2 VSS 0.0205f
C14986 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n3 VSS 0.0485f
C14987 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n4 VSS 0.0485f
C14988 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t0 VSS 0.0562f
C14989 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t1 VSS 0.0169f
C14990 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n5 VSS 0.194f
C14991 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t13 VSS 0.033f
C14992 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t9 VSS 0.0501f
C14993 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n6 VSS 0.0885f
C14994 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t5 VSS 0.033f
C14995 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t2 VSS 0.0501f
C14996 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n7 VSS 0.0885f
C14997 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t6 VSS 0.0465f
C14998 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t10 VSS 0.0259f
C14999 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n8 VSS 0.0884f
C15000 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n9 VSS 0.283f
C15001 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t3 VSS 0.033f
C15002 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t8 VSS 0.0501f
C15003 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n10 VSS 0.0885f
C15004 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t15 VSS 0.033f
C15005 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t11 VSS 0.0501f
C15006 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n11 VSS 0.0885f
C15007 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t14 VSS 0.0414f
C15008 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t7 VSS 0.0106f
C15009 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n12 VSS 0.0686f
C15010 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n13 VSS 0.66f
C15011 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n14 VSS 0.66f
C15012 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t4 VSS 0.0414f
C15013 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.t12 VSS 0.0106f
C15014 CLK_div_108_new_mag_0.CLK_div_3_mag_1.CLK.n15 VSS 0.0686f
C15015 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.n0 VSS 2.09f
C15016 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.t0 VSS 0.0341f
C15017 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.n1 VSS 0.0341f
C15018 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.n2 VSS 0.0805f
C15019 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.t2 VSS 0.0546f
C15020 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.t3 VSS 0.0704f
C15021 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.n3 VSS 0.139f
C15022 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.t4 VSS 0.0437f
C15023 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.t7 VSS 0.0545f
C15024 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.n4 VSS 0.141f
C15025 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.t5 VSS 0.0768f
C15026 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.t6 VSS 0.0489f
C15027 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.n5 VSS 0.136f
C15028 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.n6 VSS 1.17f
C15029 CLK_div_108_new_mag_0.CLK_div_3_mag_2.JK_FF_mag_1.K.n7 VSS 0.264f
C15030 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.t2 VSS 0.0246f
C15031 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.t0 VSS 0.0203f
C15032 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.n0 VSS 0.0203f
C15033 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.n1 VSS 0.0557f
C15034 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.t5 VSS 0.0632f
C15035 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.t7 VSS 0.0195f
C15036 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.n2 VSS 0.0665f
C15037 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.t8 VSS 0.0298f
C15038 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.t4 VSS 0.0452f
C15039 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.n3 VSS 0.0802f
C15040 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.t3 VSS 0.0259f
C15041 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.t6 VSS 0.0324f
C15042 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.n4 VSS 0.0753f
C15043 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.n5 VSS 0.597f
C15044 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q0.n6 VSS 0.441f
C15045 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n0 VSS 0.196f
C15046 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n1 VSS 0.191f
C15047 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n2 VSS 0.00491f
C15048 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n3 VSS 0.0761f
C15049 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n4 VSS 0.0132f
C15050 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n5 VSS 0.119f
C15051 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n6 VSS 0.0879f
C15052 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n7 VSS 0.0167f
C15053 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n8 VSS 0.0244f
C15054 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t1 VSS 0.0233f
C15055 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t2 VSS 0.0192f
C15056 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n9 VSS 0.0192f
C15057 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n10 VSS 0.0462f
C15058 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n11 VSS 0.144f
C15059 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t5 VSS 0.0428f
C15060 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t4 VSS 0.0282f
C15061 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n12 VSS 0.076f
C15062 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n13 VSS 0.298f
C15063 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t7 VSS 0.0307f
C15064 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t6 VSS 0.0246f
C15065 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n14 VSS 0.0713f
C15066 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n15 VSS 0.0442f
C15067 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n16 VSS 0.567f
C15068 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t13 VSS 0.0428f
C15069 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t8 VSS 0.0282f
C15070 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n17 VSS 0.0756f
C15071 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t11 VSS 0.0428f
C15072 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t9 VSS 0.0282f
C15073 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n18 VSS 0.0757f
C15074 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t3 VSS 0.0307f
C15075 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t16 VSS 0.0246f
C15076 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n19 VSS 0.0695f
C15077 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t15 VSS 0.0219f
C15078 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t12 VSS 0.0401f
C15079 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n20 VSS 0.0755f
C15080 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n21 VSS 0.66f
C15081 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t10 VSS 0.0353f
C15082 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.t14 VSS 0.00913f
C15083 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n22 VSS 0.0585f
C15084 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n23 VSS 0.0619f
C15085 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n24 VSS 0.144f
C15086 CLK_div_100_mag_0.CLK_div_10_mag_1.Q1.n25 VSS 0.0182f
C15087 CLK_div_96_mag_0.JK_FF_mag_4.Q.n0 VSS 0.225f
C15088 CLK_div_96_mag_0.JK_FF_mag_4.Q.t1 VSS 0.0155f
C15089 CLK_div_96_mag_0.JK_FF_mag_4.Q.t0 VSS 0.0128f
C15090 CLK_div_96_mag_0.JK_FF_mag_4.Q.n1 VSS 0.0128f
C15091 CLK_div_96_mag_0.JK_FF_mag_4.Q.n2 VSS 0.0307f
C15092 CLK_div_96_mag_0.JK_FF_mag_4.Q.t8 VSS 0.0285f
C15093 CLK_div_96_mag_0.JK_FF_mag_4.Q.t7 VSS 0.0187f
C15094 CLK_div_96_mag_0.JK_FF_mag_4.Q.n3 VSS 0.0505f
C15095 CLK_div_96_mag_0.JK_FF_mag_4.Q.t6 VSS 0.0204f
C15096 CLK_div_96_mag_0.JK_FF_mag_4.Q.t5 VSS 0.0163f
C15097 CLK_div_96_mag_0.JK_FF_mag_4.Q.n4 VSS 0.0474f
C15098 CLK_div_96_mag_0.JK_FF_mag_4.Q.n5 VSS 0.378f
C15099 CLK_div_96_mag_0.JK_FF_mag_4.Q.t12 VSS 0.0285f
C15100 CLK_div_96_mag_0.JK_FF_mag_4.Q.t11 VSS 0.0187f
C15101 CLK_div_96_mag_0.JK_FF_mag_4.Q.n6 VSS 0.0503f
C15102 CLK_div_96_mag_0.JK_FF_mag_4.Q.t3 VSS 0.0285f
C15103 CLK_div_96_mag_0.JK_FF_mag_4.Q.t4 VSS 0.0187f
C15104 CLK_div_96_mag_0.JK_FF_mag_4.Q.n7 VSS 0.0503f
C15105 CLK_div_96_mag_0.JK_FF_mag_4.Q.t10 VSS 0.0235f
C15106 CLK_div_96_mag_0.JK_FF_mag_4.Q.t9 VSS 0.00607f
C15107 CLK_div_96_mag_0.JK_FF_mag_4.Q.n8 VSS 0.039f
C15108 CLK_div_96_mag_0.JK_FF_mag_4.Q.n9 VSS 0.39f
C15109 Vdiv108.t5 VSS 0.00207f
C15110 Vdiv108.t8 VSS 0.0026f
C15111 Vdiv108.n0 VSS 0.0063f
C15112 Vdiv108.n1 VSS 0.00192f
C15113 Vdiv108.n2 VSS 0.00197f
C15114 Vdiv108.t0 VSS 0.00162f
C15115 Vdiv108.n3 VSS 0.00162f
C15116 Vdiv108.n4 VSS 0.00445f
C15117 Vdiv108.n5 VSS 0.0144f
C15118 Vdiv108.n6 VSS 0.0015f
C15119 Vdiv108.t3 VSS 0.00207f
C15120 Vdiv108.t7 VSS 0.0026f
C15121 Vdiv108.n7 VSS 0.00601f
C15122 Vdiv108.n8 VSS 0.00375f
C15123 Vdiv108.t6 VSS 0.00238f
C15124 Vdiv108.t4 VSS 0.00361f
C15125 Vdiv108.n9 VSS 0.00642f
C15126 Vdiv108.n10 VSS 0.0252f
C15127 Vdiv108.n11 VSS 0.0469f
C15128 Vdiv108.n12 VSS 0.0182f
C15129 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n0 VSS 0.317f
C15130 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.t1 VSS 0.0207f
C15131 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.t2 VSS 0.0171f
C15132 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n1 VSS 0.0171f
C15133 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n2 VSS 0.047f
C15134 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.t7 VSS 0.0273f
C15135 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.t9 VSS 0.0352f
C15136 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n3 VSS 0.0697f
C15137 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.t10 VSS 0.0218f
C15138 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.t6 VSS 0.0273f
C15139 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n4 VSS 0.0618f
C15140 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.t5 VSS 0.0251f
C15141 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.t3 VSS 0.0381f
C15142 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n5 VSS 0.0676f
C15143 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.t8 VSS 0.0218f
C15144 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.t4 VSS 0.0273f
C15145 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n6 VSS 0.0634f
C15146 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n7 VSS 0.499f
C15147 CLK_div_108_new_mag_0.CLK_div_3_mag_2.Q1.n8 VSS 0.207f
C15148 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t5 VSS 0.154f
C15149 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t7 VSS 0.0457f
C15150 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n0 VSS 0.158f
C15151 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t4 VSS 0.0621f
C15152 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t8 VSS 0.0779f
C15153 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n1 VSS 0.184f
C15154 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t6 VSS 0.109f
C15155 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t3 VSS 0.0696f
C15156 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n2 VSS 0.193f
C15157 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n3 VSS 1.79f
C15158 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n4 VSS 0.0486f
C15159 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t1 VSS 0.163f
C15160 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n5 VSS 0.377f
C15161 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n0 VSS 0.52f
C15162 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n1 VSS 0.328f
C15163 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n2 VSS 0.0208f
C15164 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n3 VSS 0.0494f
C15165 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n4 VSS 0.0494f
C15166 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t0 VSS 0.0172f
C15167 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t1 VSS 0.0571f
C15168 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n5 VSS 0.198f
C15169 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t15 VSS 0.0109f
C15170 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t7 VSS 0.042f
C15171 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n6 VSS 0.0697f
C15172 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t4 VSS 0.0509f
C15173 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t11 VSS 0.0335f
C15174 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n7 VSS 0.09f
C15175 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t6 VSS 0.0509f
C15176 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t12 VSS 0.0335f
C15177 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n8 VSS 0.09f
C15178 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t9 VSS 0.0509f
C15179 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t14 VSS 0.0335f
C15180 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n9 VSS 0.09f
C15181 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t8 VSS 0.0264f
C15182 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t5 VSS 0.0472f
C15183 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n10 VSS 0.0899f
C15184 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n11 VSS 0.288f
C15185 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t2 VSS 0.0509f
C15186 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t10 VSS 0.0335f
C15187 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n12 VSS 0.09f
C15188 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t3 VSS 0.042f
C15189 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.t13 VSS 0.0109f
C15190 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n13 VSS 0.0697f
C15191 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n14 VSS 0.67f
C15192 CLK_div_99_mag_0.CLK_div_3_mag_0.CLK.n15 VSS 0.671f
C15193 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n0 VSS 2.13f
C15194 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t1 VSS 0.0354f
C15195 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n1 VSS 0.0354f
C15196 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n2 VSS 0.0755f
C15197 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t5 VSS 0.0797f
C15198 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t2 VSS 0.0507f
C15199 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n3 VSS 0.141f
C15200 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t7 VSS 0.0568f
C15201 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t3 VSS 0.0729f
C15202 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n4 VSS 0.145f
C15203 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t4 VSS 0.0566f
C15204 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t6 VSS 0.0453f
C15205 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n5 VSS 0.134f
C15206 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n6 VSS 1.21f
C15207 CLK_div_90_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n7 VSS 0.221f
C15208 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n0 VSS 2.15f
C15209 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n1 VSS 0.208f
C15210 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t8 VSS 0.0724f
C15211 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t6 VSS 0.0562f
C15212 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n2 VSS 0.143f
C15213 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t3 VSS 0.0449f
C15214 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t7 VSS 0.0563f
C15215 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n3 VSS 0.145f
C15216 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t4 VSS 0.079f
C15217 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t5 VSS 0.0503f
C15218 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n4 VSS 0.14f
C15219 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n5 VSS 1.2f
C15220 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t0 VSS 0.0351f
C15221 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n6 VSS 0.0351f
C15222 CLK_div_93_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n7 VSS 0.0828f
C15223 Vdiv110.n0 VSS 0.00199f
C15224 Vdiv110.n1 VSS 0.00104f
C15225 Vdiv110.n2 VSS 9.7e-19
C15226 Vdiv110.t4 VSS 0.00399f
C15227 Vdiv110.t5 VSS 0.00218f
C15228 Vdiv110.n3 VSS 0.00749f
C15229 Vdiv110.n4 VSS 6.46e-19
C15230 Vdiv110.n5 VSS 4.96e-19
C15231 Vdiv110.n6 VSS 5.03e-19
C15232 Vdiv110.n7 VSS 1.57f
C15233 Vdiv110.t0 VSS 6.2e-19
C15234 Vdiv110.n8 VSS 6.2e-19
C15235 Vdiv110.n9 VSS 0.00297f
C15236 Vdiv110.n10 VSS 0.00141f
C15237 Vdiv110.n11 VSS 0.0151f
C15238 Vdiv110.n12 VSS 0.0186f
C15239 Vdiv110.n13 VSS 0.0214f
C15240 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.t1 VSS 0.021f
C15241 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.t0 VSS 0.0173f
C15242 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n0 VSS 0.0173f
C15243 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n1 VSS 0.0415f
C15244 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.t9 VSS 0.0276f
C15245 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.t8 VSS 0.0221f
C15246 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n2 VSS 0.0625f
C15247 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.t5 VSS 0.0277f
C15248 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.t7 VSS 0.0355f
C15249 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n3 VSS 0.0706f
C15250 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n4 VSS 0.321f
C15251 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.t3 VSS 0.0385f
C15252 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.t10 VSS 0.0254f
C15253 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n5 VSS 0.0684f
C15254 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.t6 VSS 0.0276f
C15255 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.t4 VSS 0.0221f
C15256 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n6 VSS 0.0642f
C15257 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n7 VSS 0.505f
C15258 CLK_div_90_mag_0.CLK_div_3_mag_1.Q1.n8 VSS 0.209f
C15259 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.t2 VSS 0.021f
C15260 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.t0 VSS 0.0173f
C15261 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n0 VSS 0.0173f
C15262 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n1 VSS 0.0415f
C15263 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.t10 VSS 0.0276f
C15264 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.t9 VSS 0.0221f
C15265 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n2 VSS 0.0625f
C15266 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.t5 VSS 0.0277f
C15267 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.t8 VSS 0.0355f
C15268 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n3 VSS 0.0706f
C15269 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n4 VSS 0.321f
C15270 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.t7 VSS 0.0385f
C15271 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.t3 VSS 0.0254f
C15272 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n5 VSS 0.0684f
C15273 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.t4 VSS 0.0276f
C15274 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.t6 VSS 0.0221f
C15275 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n6 VSS 0.0642f
C15276 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n7 VSS 0.505f
C15277 CLK_div_99_mag_0.CLK_div_3_mag_0.Q1.n8 VSS 0.209f
C15278 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t3 VSS 0.154f
C15279 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t6 VSS 0.0457f
C15280 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n0 VSS 0.158f
C15281 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t8 VSS 0.0621f
C15282 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t5 VSS 0.0779f
C15283 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n1 VSS 0.184f
C15284 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t4 VSS 0.109f
C15285 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t7 VSS 0.0696f
C15286 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n2 VSS 0.193f
C15287 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.n3 VSS 1.79f
C15288 CLK_div_110_mag_0.CLK_DIV_11_mag_new_0.or_2_mag_3.IN1.t0 VSS 0.589f
C15289 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t2 VSS 0.0207f
C15290 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t4 VSS 0.0271f
C15291 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n0 VSS 0.0537f
C15292 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t5 VSS 0.0273f
C15293 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.t3 VSS 0.0207f
C15294 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n1 VSS 0.0537f
C15295 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n2 VSS 0.675f
C15296 CLK_div_99_mag_0.CLK_DIV_11_mag_new_0.JK_FF_mag_1.K.n3 VSS 0.0327f
C15297 CLK_div_96_mag_0.JK_FF_mag_5.Q.n0 VSS 0.25f
C15298 CLK_div_96_mag_0.JK_FF_mag_5.Q.t0 VSS 0.0172f
C15299 CLK_div_96_mag_0.JK_FF_mag_5.Q.t2 VSS 0.0142f
C15300 CLK_div_96_mag_0.JK_FF_mag_5.Q.n1 VSS 0.0142f
C15301 CLK_div_96_mag_0.JK_FF_mag_5.Q.n2 VSS 0.0341f
C15302 CLK_div_96_mag_0.JK_FF_mag_5.Q.t3 VSS 0.0208f
C15303 CLK_div_96_mag_0.JK_FF_mag_5.Q.t11 VSS 0.0316f
C15304 CLK_div_96_mag_0.JK_FF_mag_5.Q.n3 VSS 0.0559f
C15305 CLK_div_96_mag_0.JK_FF_mag_5.Q.t12 VSS 0.0208f
C15306 CLK_div_96_mag_0.JK_FF_mag_5.Q.t10 VSS 0.0316f
C15307 CLK_div_96_mag_0.JK_FF_mag_5.Q.n4 VSS 0.0559f
C15308 CLK_div_96_mag_0.JK_FF_mag_5.Q.t7 VSS 0.00668f
C15309 CLK_div_96_mag_0.JK_FF_mag_5.Q.t4 VSS 0.0261f
C15310 CLK_div_96_mag_0.JK_FF_mag_5.Q.n5 VSS 0.0433f
C15311 CLK_div_96_mag_0.JK_FF_mag_5.Q.t9 VSS 0.0316f
C15312 CLK_div_96_mag_0.JK_FF_mag_5.Q.t8 VSS 0.0208f
C15313 CLK_div_96_mag_0.JK_FF_mag_5.Q.n6 VSS 0.0562f
C15314 CLK_div_96_mag_0.JK_FF_mag_5.Q.t6 VSS 0.0227f
C15315 CLK_div_96_mag_0.JK_FF_mag_5.Q.t5 VSS 0.0182f
C15316 CLK_div_96_mag_0.JK_FF_mag_5.Q.n7 VSS 0.0527f
C15317 CLK_div_96_mag_0.JK_FF_mag_5.Q.n8 VSS 0.419f
C15318 CLK_div_96_mag_0.JK_FF_mag_5.Q.n9 VSS 0.295f
C15319 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t1 VSS 0.0149f
C15320 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n0 VSS 0.0149f
C15321 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n1 VSS 0.0318f
C15322 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t3 VSS 0.0238f
C15323 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t2 VSS 0.0308f
C15324 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n2 VSS 0.0609f
C15325 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t7 VSS 0.0335f
C15326 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t6 VSS 0.0214f
C15327 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n3 VSS 0.0593f
C15328 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n4 VSS 1.14f
C15329 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t5 VSS 0.0238f
C15330 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t4 VSS 0.0191f
C15331 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n5 VSS 0.0566f
C15332 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n6 VSS 0.381f
C15333 CLK_div_105_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n7 VSS 0.0932f
C15334 Vdiv105.t4 VSS 0.00875f
C15335 Vdiv105.t5 VSS 0.00478f
C15336 Vdiv105.n0 VSS 0.0165f
C15337 Vdiv105.t0 VSS 0.00136f
C15338 Vdiv105.n1 VSS 0.00136f
C15339 Vdiv105.n2 VSS 0.00652f
C15340 Vdiv105.t1 VSS 0.00311f
C15341 Vdiv105.n3 VSS 0.0331f
C15342 Vdiv105.n4 VSS 0.00473f
C15343 Vdiv105.t2 VSS 0.0392f
C15344 Vdiv105.n5 VSS 0.138f
C15345 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n0 VSS 2.07f
C15346 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t0 VSS 0.0344f
C15347 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n1 VSS 0.0344f
C15348 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n2 VSS 0.0734f
C15349 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t6 VSS 0.0774f
C15350 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t3 VSS 0.0493f
C15351 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n3 VSS 0.137f
C15352 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t4 VSS 0.0552f
C15353 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t7 VSS 0.0708f
C15354 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n4 VSS 0.141f
C15355 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t5 VSS 0.055f
C15356 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t2 VSS 0.044f
C15357 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n5 VSS 0.131f
C15358 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n6 VSS 1.18f
C15359 CLK_div_99_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n7 VSS 0.215f
C15360 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n0 VSS 0.0877f
C15361 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t5 VSS 0.0189f
C15362 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t6 VSS 0.0237f
C15363 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n1 VSS 0.0561f
C15364 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t4 VSS 0.0333f
C15365 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t3 VSS 0.0212f
C15366 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n2 VSS 0.0588f
C15367 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t7 VSS 0.0306f
C15368 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t8 VSS 0.0235f
C15369 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n3 VSS 0.0604f
C15370 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n4 VSS 1.13f
C15371 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n5 VSS 0.378f
C15372 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t1 VSS 0.0148f
C15373 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n6 VSS 0.0148f
C15374 CLK_div_105_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n7 VSS 0.0349f
C15375 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.t2 VSS 0.025f
C15376 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.t0 VSS 0.0206f
C15377 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.n0 VSS 0.0206f
C15378 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.n1 VSS 0.0494f
C15379 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.t8 VSS 0.0459f
C15380 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.t4 VSS 0.0302f
C15381 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.n2 VSS 0.0814f
C15382 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.t7 VSS 0.0329f
C15383 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.t3 VSS 0.0263f
C15384 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.n3 VSS 0.0764f
C15385 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.n4 VSS 0.606f
C15386 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.t6 VSS 0.0641f
C15387 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.t5 VSS 0.0199f
C15388 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.n5 VSS 0.0675f
C15389 CLK_div_99_mag_0.CLK_div_3_mag_1.Q0.n6 VSS 0.447f
C15390 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.t0 VSS 0.025f
C15391 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.t2 VSS 0.0206f
C15392 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.n0 VSS 0.0206f
C15393 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.n1 VSS 0.0494f
C15394 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.t6 VSS 0.0459f
C15395 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.t4 VSS 0.0302f
C15396 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.n2 VSS 0.0814f
C15397 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.t7 VSS 0.0329f
C15398 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.t5 VSS 0.0263f
C15399 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.n3 VSS 0.0764f
C15400 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.n4 VSS 0.606f
C15401 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.t3 VSS 0.0641f
C15402 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.t8 VSS 0.0199f
C15403 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.n5 VSS 0.0675f
C15404 CLK_div_90_mag_0.CLK_div_3_mag_1.Q0.n6 VSS 0.447f
C15405 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t2 VSS 0.02f
C15406 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t0 VSS 0.0165f
C15407 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n0 VSS 0.0165f
C15408 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n1 VSS 0.0396f
C15409 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t10 VSS 0.0367f
C15410 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t9 VSS 0.0242f
C15411 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n2 VSS 0.0652f
C15412 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t8 VSS 0.0263f
C15413 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t7 VSS 0.0211f
C15414 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n3 VSS 0.0612f
C15415 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n4 VSS 0.486f
C15416 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t11 VSS 0.019f
C15417 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t6 VSS 0.034f
C15418 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n5 VSS 0.0648f
C15419 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t5 VSS 0.0263f
C15420 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t3 VSS 0.0211f
C15421 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n6 VSS 0.0612f
C15422 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n7 VSS 0.325f
C15423 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t4 VSS 0.0263f
C15424 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.t12 VSS 0.0211f
C15425 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n8 VSS 0.0612f
C15426 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n9 VSS 0.308f
C15427 CLK_div_100_mag_0.CLK_div_10_mag_1.Q2.n10 VSS 0.15f
C15428 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n0 VSS 2.12f
C15429 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t0 VSS 0.0346f
C15430 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n1 VSS 0.0346f
C15431 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n2 VSS 0.0817f
C15432 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t7 VSS 0.0554f
C15433 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t2 VSS 0.0714f
C15434 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n3 VSS 0.141f
C15435 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t6 VSS 0.0443f
C15436 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t3 VSS 0.0553f
C15437 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n4 VSS 0.143f
C15438 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t4 VSS 0.0779f
C15439 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t5 VSS 0.0496f
C15440 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n5 VSS 0.138f
C15441 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n6 VSS 1.18f
C15442 CLK_div_108_new_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n7 VSS 0.268f
C15443 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n0 VSS 0.109f
C15444 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n1 VSS 0.0183f
C15445 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t0 VSS 0.0256f
C15446 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t2 VSS 0.0211f
C15447 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n2 VSS 0.0211f
C15448 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n3 VSS 0.0508f
C15449 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n4 VSS 0.158f
C15450 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n5 VSS 0.0296f
C15451 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t13 VSS 0.0388f
C15452 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t12 VSS 0.0101f
C15453 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n6 VSS 0.0644f
C15454 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n7 VSS 0.00386f
C15455 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n8 VSS 0.0154f
C15456 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t5 VSS 0.0471f
C15457 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t9 VSS 0.031f
C15458 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n9 VSS 0.0832f
C15459 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n10 VSS 0.0109f
C15460 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n11 VSS 0.00782f
C15461 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n12 VSS 0.0039f
C15462 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n13 VSS 0.156f
C15463 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t15 VSS 0.0471f
C15464 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t4 VSS 0.031f
C15465 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n14 VSS 0.0832f
C15466 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n15 VSS 0.0109f
C15467 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n16 VSS 0.00782f
C15468 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n17 VSS 0.154f
C15469 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n18 VSS 0.0951f
C15470 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n19 VSS 0.1f
C15471 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t10 VSS 0.0471f
C15472 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t14 VSS 0.031f
C15473 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n20 VSS 0.0836f
C15474 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n21 VSS 0.0283f
C15475 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t11 VSS 0.0441f
C15476 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t8 VSS 0.0241f
C15477 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n22 VSS 0.0838f
C15478 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t3 VSS 0.0241f
C15479 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t7 VSS 0.0441f
C15480 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n23 VSS 0.0838f
C15481 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n24 VSS 0.479f
C15482 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n25 VSS 0.725f
C15483 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t16 VSS 0.0338f
C15484 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.t6 VSS 0.027f
C15485 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n26 VSS 0.0785f
C15486 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n27 VSS 0.0487f
C15487 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n28 VSS 0.5f
C15488 CLK_div_93_mag_0.CLK_div_31_mag_0.Q0.n29 VSS 0.02f
C15489 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n0 VSS 2.15f
C15490 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n1 VSS 0.208f
C15491 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t6 VSS 0.0724f
C15492 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t7 VSS 0.0562f
C15493 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n2 VSS 0.143f
C15494 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t8 VSS 0.0449f
C15495 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t3 VSS 0.0563f
C15496 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n3 VSS 0.145f
C15497 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t5 VSS 0.079f
C15498 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t4 VSS 0.0503f
C15499 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n4 VSS 0.14f
C15500 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n5 VSS 1.2f
C15501 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t2 VSS 0.0351f
C15502 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n6 VSS 0.0351f
C15503 CLK_div_96_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n7 VSS 0.0828f
C15504 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n0 VSS 0.826f
C15505 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n1 VSS 0.0344f
C15506 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n2 VSS 0.254f
C15507 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n3 VSS 0.0151f
C15508 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n4 VSS 0.241f
C15509 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n5 VSS 0.0151f
C15510 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n6 VSS 0.15f
C15511 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n7 VSS 0.103f
C15512 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n8 VSS 0.103f
C15513 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n9 VSS 0.035f
C15514 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t1 VSS 0.0201f
C15515 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t2 VSS 0.0165f
C15516 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n10 VSS 0.0165f
C15517 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n11 VSS 0.0397f
C15518 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n12 VSS 0.124f
C15519 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t18 VSS 0.0368f
C15520 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t11 VSS 0.0243f
C15521 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n13 VSS 0.0654f
C15522 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n14 VSS 0.257f
C15523 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t13 VSS 0.0264f
C15524 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t5 VSS 0.0211f
C15525 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n15 VSS 0.0614f
C15526 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n16 VSS 0.0381f
C15527 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n17 VSS 0.488f
C15528 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t9 VSS 0.0368f
C15529 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t8 VSS 0.0243f
C15530 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n18 VSS 0.0651f
C15531 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t7 VSS 0.0368f
C15532 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t6 VSS 0.0243f
C15533 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n19 VSS 0.0651f
C15534 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t3 VSS 0.0304f
C15535 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t10 VSS 0.00786f
C15536 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n20 VSS 0.0504f
C15537 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t14 VSS 0.0368f
C15538 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t4 VSS 0.0243f
C15539 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n21 VSS 0.0651f
C15540 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t16 VSS 0.0368f
C15541 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t15 VSS 0.0243f
C15542 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n22 VSS 0.0651f
C15543 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n23 VSS 0.11f
C15544 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t19 VSS 0.0342f
C15545 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t20 VSS 0.0189f
C15546 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n24 VSS 0.0652f
C15547 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n25 VSS 0.869f
C15548 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t12 VSS 0.0304f
C15549 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.t17 VSS 0.00786f
C15550 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n26 VSS 0.0504f
C15551 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n27 VSS 0.124f
C15552 CLK_div_105_mag_0.CLK_div_10_mag_1.Q0.n28 VSS 0.0156f
C15553 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.t0 VSS 0.0246f
C15554 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.t2 VSS 0.0203f
C15555 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.n0 VSS 0.0203f
C15556 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.n1 VSS 0.0557f
C15557 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.t8 VSS 0.0632f
C15558 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.t5 VSS 0.0195f
C15559 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.n2 VSS 0.0665f
C15560 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.t7 VSS 0.0298f
C15561 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.t3 VSS 0.0452f
C15562 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.n3 VSS 0.0802f
C15563 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.t4 VSS 0.0259f
C15564 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.t6 VSS 0.0324f
C15565 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.n4 VSS 0.0753f
C15566 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.n5 VSS 0.597f
C15567 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q0.n6 VSS 0.441f
C15568 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n0 VSS 0.196f
C15569 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n1 VSS 0.191f
C15570 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n2 VSS 0.00491f
C15571 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n3 VSS 0.0761f
C15572 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n4 VSS 0.0132f
C15573 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n5 VSS 0.119f
C15574 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n6 VSS 0.0879f
C15575 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n7 VSS 0.0167f
C15576 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n8 VSS 0.0244f
C15577 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t1 VSS 0.0233f
C15578 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t2 VSS 0.0192f
C15579 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n9 VSS 0.0192f
C15580 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n10 VSS 0.0462f
C15581 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n11 VSS 0.144f
C15582 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t9 VSS 0.0428f
C15583 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t10 VSS 0.0282f
C15584 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n12 VSS 0.076f
C15585 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n13 VSS 0.298f
C15586 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t8 VSS 0.0307f
C15587 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t11 VSS 0.0246f
C15588 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n14 VSS 0.0713f
C15589 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n15 VSS 0.0442f
C15590 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n16 VSS 0.567f
C15591 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t14 VSS 0.0428f
C15592 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t12 VSS 0.0282f
C15593 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n17 VSS 0.0756f
C15594 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t15 VSS 0.0428f
C15595 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t16 VSS 0.0282f
C15596 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n18 VSS 0.0757f
C15597 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t5 VSS 0.0307f
C15598 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t4 VSS 0.0246f
C15599 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n19 VSS 0.0695f
C15600 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t7 VSS 0.0219f
C15601 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t6 VSS 0.0401f
C15602 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n20 VSS 0.0755f
C15603 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n21 VSS 0.66f
C15604 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t13 VSS 0.0353f
C15605 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.t3 VSS 0.00913f
C15606 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n22 VSS 0.0585f
C15607 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n23 VSS 0.0619f
C15608 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n24 VSS 0.144f
C15609 CLK_div_105_mag_0.CLK_div_10_mag_1.Q1.n25 VSS 0.0182f
C15610 CLK.n0 VSS 0.207f
C15611 CLK.n1 VSS 7.41e-19
C15612 CLK.t65 VSS 0.00294f
C15613 CLK.t76 VSS 0.00447f
C15614 CLK.n2 VSS 0.00789f
C15615 CLK.n3 VSS 0.00102f
C15616 CLK.n4 VSS 3.7e-19
C15617 CLK.n5 VSS 0.00144f
C15618 CLK.n6 VSS 0.0146f
C15619 CLK.n7 VSS 0.0148f
C15620 CLK.n8 VSS 7.41e-19
C15621 CLK.t78 VSS 0.00294f
C15622 CLK.t92 VSS 0.00447f
C15623 CLK.n9 VSS 0.00789f
C15624 CLK.n10 VSS 0.00102f
C15625 CLK.n11 VSS 3.66e-19
C15626 CLK.n12 VSS 0.00903f
C15627 CLK.n13 VSS 0.0096f
C15628 CLK.n14 VSS 0.00141f
C15629 CLK.n15 VSS 6.51e-19
C15630 CLK.n16 VSS 3.98e-19
C15631 CLK.n17 VSS 0.00318f
C15632 CLK.t42 VSS 0.00364f
C15633 CLK.n18 VSS 0.00413f
C15634 CLK.t51 VSS 8.84e-19
C15635 CLK.n19 VSS 0.00209f
C15636 CLK.n20 VSS 2.6e-19
C15637 CLK.n21 VSS 4.16e-19
C15638 CLK.n22 VSS 1.04e-19
C15639 CLK.n23 VSS 0.00709f
C15640 CLK.n24 VSS 0.0538f
C15641 CLK.n25 VSS 0.00128f
C15642 CLK.t6 VSS 0.00369f
C15643 CLK.t93 VSS 9.43e-19
C15644 CLK.n26 VSS 0.00611f
C15645 CLK.n27 VSS 0.0013f
C15646 CLK.n28 VSS 0.00231f
C15647 CLK.n29 VSS 4.51e-19
C15648 CLK.n30 VSS 4e-19
C15649 CLK.n31 VSS 7.41e-19
C15650 CLK.t83 VSS 0.00294f
C15651 CLK.t70 VSS 0.00447f
C15652 CLK.n32 VSS 0.00789f
C15653 CLK.n33 VSS 0.00102f
C15654 CLK.n34 VSS 3.72e-19
C15655 CLK.n35 VSS 0.00162f
C15656 CLK.n36 VSS 0.00713f
C15657 CLK.n37 VSS 0.0143f
C15658 CLK.n38 VSS 2.13e-19
C15659 CLK.n39 VSS 7.41e-19
C15660 CLK.t30 VSS 0.00294f
C15661 CLK.t29 VSS 0.00447f
C15662 CLK.n40 VSS 0.00789f
C15663 CLK.n41 VSS 0.00102f
C15664 CLK.n42 VSS 3.63e-19
C15665 CLK.n43 VSS 4.8e-19
C15666 CLK.n44 VSS 1.75e-19
C15667 CLK.n45 VSS 0.0156f
C15668 CLK.n46 VSS 0.0864f
C15669 CLK.n47 VSS 0.293f
C15670 CLK.n48 VSS 4.06f
C15671 CLK.n49 VSS 4.51e-19
C15672 CLK.t89 VSS 9.53e-19
C15673 CLK.t64 VSS 0.00368f
C15674 CLK.n50 VSS 0.00611f
C15675 CLK.n51 VSS 0.0013f
C15676 CLK.n52 VSS 3.66e-19
C15677 CLK.n53 VSS 0.00146f
C15678 CLK.t41 VSS 0.00447f
C15679 CLK.t18 VSS 0.00294f
C15680 CLK.n54 VSS 0.00789f
C15681 CLK.n55 VSS 0.00103f
C15682 CLK.n56 VSS 7.41e-19
C15683 CLK.n57 VSS 3.7e-19
C15684 CLK.n58 VSS 0.0148f
C15685 CLK.t91 VSS 0.00447f
C15686 CLK.t33 VSS 0.00294f
C15687 CLK.n59 VSS 0.00789f
C15688 CLK.n60 VSS 0.00103f
C15689 CLK.n61 VSS 7.41e-19
C15690 CLK.n62 VSS 0.0146f
C15691 CLK.n63 VSS 0.00854f
C15692 CLK.n64 VSS 3.66e-19
C15693 CLK.n65 VSS 0.00146f
C15694 CLK.t14 VSS 0.00447f
C15695 CLK.t82 VSS 0.00294f
C15696 CLK.n66 VSS 0.00789f
C15697 CLK.n67 VSS 0.00103f
C15698 CLK.n68 VSS 7.41e-19
C15699 CLK.n69 VSS 3.7e-19
C15700 CLK.n70 VSS 0.0138f
C15701 CLK.t54 VSS 0.00232f
C15702 CLK.t47 VSS 0.00414f
C15703 CLK.n71 VSS 0.00788f
C15704 CLK.n72 VSS 0.0253f
C15705 CLK.n73 VSS 0.0304f
C15706 CLK.t27 VSS 0.00447f
C15707 CLK.t71 VSS 0.00294f
C15708 CLK.n74 VSS 0.00789f
C15709 CLK.n75 VSS 0.00103f
C15710 CLK.n76 VSS 7.41e-19
C15711 CLK.n77 VSS 0.00114f
C15712 CLK.n78 VSS 0.00854f
C15713 CLK.n79 VSS 0.00159f
C15714 CLK.n80 VSS 0.00265f
C15715 CLK.t77 VSS 0.00368f
C15716 CLK.t45 VSS 9.53e-19
C15717 CLK.n81 VSS 0.00611f
C15718 CLK.n82 VSS 0.0013f
C15719 CLK.n83 VSS 4.51e-19
C15720 CLK.n84 VSS 9.65e-19
C15721 CLK.n85 VSS 0.0564f
C15722 CLK.n86 VSS 0.0565f
C15723 CLK.n87 VSS 9.65e-19
C15724 CLK.n88 VSS 0.00159f
C15725 CLK.n89 VSS 0.00125f
C15726 CLK.n90 VSS 1.75f
C15727 CLK.n91 VSS 4.51e-19
C15728 CLK.n92 VSS 3.66e-19
C15729 CLK.n93 VSS 0.00146f
C15730 CLK.t25 VSS 0.00447f
C15731 CLK.t20 VSS 0.00294f
C15732 CLK.n94 VSS 0.00789f
C15733 CLK.n95 VSS 0.00103f
C15734 CLK.n96 VSS 7.41e-19
C15735 CLK.n97 VSS 3.7e-19
C15736 CLK.n98 VSS 0.0148f
C15737 CLK.t87 VSS 0.00447f
C15738 CLK.t15 VSS 0.00294f
C15739 CLK.n99 VSS 0.00789f
C15740 CLK.n100 VSS 0.00103f
C15741 CLK.n101 VSS 7.41e-19
C15742 CLK.n102 VSS 0.0146f
C15743 CLK.n103 VSS 0.00933f
C15744 CLK.n104 VSS 0.00926f
C15745 CLK.t67 VSS 0.00368f
C15746 CLK.t74 VSS 9.53e-19
C15747 CLK.n105 VSS 0.00611f
C15748 CLK.n106 VSS 0.0013f
C15749 CLK.n107 VSS 0.00131f
C15750 CLK.n108 VSS 0.00265f
C15751 CLK.n109 VSS 2.3f
C15752 CLK.t7 VSS 0.00256f
C15753 CLK.t79 VSS 0.00321f
C15754 CLK.n110 VSS 0.0076f
C15755 CLK.n111 VSS 0.0552f
C15756 CLK.n112 VSS 0.103f
C15757 CLK.n113 VSS 0.039f
C15758 CLK.n114 VSS 7.7e-19
C15759 CLK.t81 VSS 0.00368f
C15760 CLK.t66 VSS 9.53e-19
C15761 CLK.n115 VSS 0.00611f
C15762 CLK.n116 VSS 0.0013f
C15763 CLK.n117 VSS 4.51e-19
C15764 CLK.t50 VSS 0.00447f
C15765 CLK.t84 VSS 0.00294f
C15766 CLK.n118 VSS 0.00789f
C15767 CLK.n119 VSS 0.00103f
C15768 CLK.n120 VSS 7.41e-19
C15769 CLK.n121 VSS 3.66e-19
C15770 CLK.n122 VSS 7.41e-19
C15771 CLK.n123 VSS 3.7e-19
C15772 CLK.t88 VSS 0.00447f
C15773 CLK.t17 VSS 0.00294f
C15774 CLK.n124 VSS 0.00789f
C15775 CLK.n125 VSS 0.00103f
C15776 CLK.n126 VSS 0.00146f
C15777 CLK.n127 VSS 0.0148f
C15778 CLK.n128 VSS 0.0146f
C15779 CLK.n129 VSS 0.0093f
C15780 CLK.n130 VSS 0.00939f
C15781 CLK.n131 VSS 0.00188f
C15782 CLK.n132 VSS 0.00148f
C15783 CLK.n133 VSS 9.51e-19
C15784 CLK.n134 VSS 0.00203f
C15785 CLK.n135 VSS 0.00249f
C15786 CLK.n136 VSS 0.00206f
C15787 CLK.n137 VSS 0.00101f
C15788 CLK.n138 VSS 7.6e-19
C15789 CLK.n139 VSS 0.00141f
C15790 CLK.n140 VSS 0.0287f
C15791 CLK.n141 VSS 0.174f
C15792 CLK.n142 VSS 0.317f
C15793 CLK.n143 VSS 4.51e-19
C15794 CLK.n144 VSS 3.7e-19
C15795 CLK.t28 VSS 0.00294f
C15796 CLK.t32 VSS 0.00447f
C15797 CLK.n145 VSS 0.00789f
C15798 CLK.n146 VSS 0.00103f
C15799 CLK.n147 VSS 7.41e-19
C15800 CLK.n148 VSS 0.00144f
C15801 CLK.n149 VSS 0.0146f
C15802 CLK.n150 VSS 0.0148f
C15803 CLK.t72 VSS 0.00294f
C15804 CLK.t60 VSS 0.00447f
C15805 CLK.n151 VSS 0.00789f
C15806 CLK.n152 VSS 0.00103f
C15807 CLK.n153 VSS 7.41e-19
C15808 CLK.n154 VSS 3.66e-19
C15809 CLK.n155 VSS 0.00854f
C15810 CLK.t35 VSS 0.00231f
C15811 CLK.t63 VSS 0.00415f
C15812 CLK.n156 VSS 0.00789f
C15813 CLK.n157 VSS 0.0253f
C15814 CLK.n158 VSS 3.7e-19
C15815 CLK.t31 VSS 0.00294f
C15816 CLK.t62 VSS 0.00447f
C15817 CLK.n159 VSS 0.00789f
C15818 CLK.n160 VSS 0.00103f
C15819 CLK.n161 VSS 7.41e-19
C15820 CLK.n162 VSS 0.00144f
C15821 CLK.n163 VSS 0.0136f
C15822 CLK.n164 VSS 0.0306f
C15823 CLK.n165 VSS 0.00114f
C15824 CLK.t9 VSS 0.00294f
C15825 CLK.t0 VSS 0.00447f
C15826 CLK.n166 VSS 0.00789f
C15827 CLK.n167 VSS 0.00103f
C15828 CLK.n168 VSS 7.41e-19
C15829 CLK.n169 VSS 3.66e-19
C15830 CLK.n170 VSS 0.00854f
C15831 CLK.n171 VSS 0.00155f
C15832 CLK.n172 VSS 0.00265f
C15833 CLK.t19 VSS 0.00369f
C15834 CLK.t73 VSS 9.43e-19
C15835 CLK.n173 VSS 0.00611f
C15836 CLK.n174 VSS 0.0013f
C15837 CLK.n175 VSS 4.51e-19
C15838 CLK.n176 VSS 9.85e-19
C15839 CLK.n177 VSS 0.0564f
C15840 CLK.n178 VSS 0.0565f
C15841 CLK.n179 VSS 9.85e-19
C15842 CLK.t46 VSS 0.00369f
C15843 CLK.t11 VSS 9.43e-19
C15844 CLK.n180 VSS 0.00611f
C15845 CLK.n181 VSS 0.0013f
C15846 CLK.n182 VSS 0.00155f
C15847 CLK.n183 VSS 0.00125f
C15848 CLK.n184 VSS 11.6f
C15849 CLK.n185 VSS 4.51e-19
C15850 CLK.n186 VSS 3.7e-19
C15851 CLK.n187 VSS 7.41e-19
C15852 CLK.t3 VSS 0.00294f
C15853 CLK.t53 VSS 0.00447f
C15854 CLK.n188 VSS 0.00789f
C15855 CLK.n189 VSS 0.00102f
C15856 CLK.n190 VSS 0.00144f
C15857 CLK.n191 VSS 0.0146f
C15858 CLK.n192 VSS 0.0148f
C15859 CLK.n193 VSS 7.41e-19
C15860 CLK.t49 VSS 0.00294f
C15861 CLK.t16 VSS 0.00447f
C15862 CLK.n194 VSS 0.00789f
C15863 CLK.n195 VSS 0.00102f
C15864 CLK.n196 VSS 3.66e-19
C15865 CLK.n197 VSS 0.00935f
C15866 CLK.n198 VSS 0.00927f
C15867 CLK.n199 VSS 4.51e-19
C15868 CLK.n200 VSS 3.7e-19
C15869 CLK.n201 VSS 7.41e-19
C15870 CLK.t37 VSS 0.00294f
C15871 CLK.t5 VSS 0.00447f
C15872 CLK.n202 VSS 0.00789f
C15873 CLK.n203 VSS 0.00102f
C15874 CLK.n204 VSS 0.00144f
C15875 CLK.n205 VSS 0.0146f
C15876 CLK.n206 VSS 0.0148f
C15877 CLK.n207 VSS 7.41e-19
C15878 CLK.t61 VSS 0.00294f
C15879 CLK.t24 VSS 0.00447f
C15880 CLK.n208 VSS 0.00789f
C15881 CLK.n209 VSS 0.00102f
C15882 CLK.n210 VSS 3.66e-19
C15883 CLK.n211 VSS 0.00935f
C15884 CLK.n212 VSS 0.00927f
C15885 CLK.t59 VSS 0.00369f
C15886 CLK.t26 VSS 9.43e-19
C15887 CLK.n213 VSS 0.00611f
C15888 CLK.n214 VSS 0.0013f
C15889 CLK.n215 VSS 0.00128f
C15890 CLK.n216 VSS 0.00265f
C15891 CLK.n217 VSS 4.51e-19
C15892 CLK.n218 VSS 3.7e-19
C15893 CLK.n219 VSS 7.41e-19
C15894 CLK.t34 VSS 0.00294f
C15895 CLK.t4 VSS 0.00447f
C15896 CLK.n220 VSS 0.00789f
C15897 CLK.n221 VSS 0.00102f
C15898 CLK.n222 VSS 0.00144f
C15899 CLK.n223 VSS 0.0146f
C15900 CLK.n224 VSS 0.0148f
C15901 CLK.n225 VSS 7.41e-19
C15902 CLK.t58 VSS 0.00294f
C15903 CLK.t48 VSS 0.00447f
C15904 CLK.n226 VSS 0.00789f
C15905 CLK.n227 VSS 0.00102f
C15906 CLK.n228 VSS 3.66e-19
C15907 CLK.n229 VSS 0.00935f
C15908 CLK.n230 VSS 0.00927f
C15909 CLK.t56 VSS 0.00369f
C15910 CLK.t23 VSS 9.43e-19
C15911 CLK.n231 VSS 0.00611f
C15912 CLK.n232 VSS 0.0013f
C15913 CLK.n233 VSS 0.00128f
C15914 CLK.n234 VSS 0.00265f
C15915 CLK.n235 VSS 0.00238f
C15916 CLK.n236 VSS 4e-19
C15917 CLK.t52 VSS 0.00294f
C15918 CLK.t22 VSS 0.00447f
C15919 CLK.n237 VSS 0.00792f
C15920 CLK.n238 VSS 0.00119f
C15921 CLK.n239 VSS 4.86e-19
C15922 CLK.n240 VSS 0.0399f
C15923 CLK.n241 VSS 4.51e-19
C15924 CLK.n242 VSS 3.7e-19
C15925 CLK.n243 VSS 7.41e-19
C15926 CLK.t86 VSS 0.00294f
C15927 CLK.t40 VSS 0.00447f
C15928 CLK.n244 VSS 0.00789f
C15929 CLK.n245 VSS 0.00102f
C15930 CLK.n246 VSS 0.00144f
C15931 CLK.n247 VSS 0.0146f
C15932 CLK.n248 VSS 0.0148f
C15933 CLK.n249 VSS 7.41e-19
C15934 CLK.t10 VSS 0.00294f
C15935 CLK.t68 VSS 0.00447f
C15936 CLK.n250 VSS 0.00789f
C15937 CLK.n251 VSS 0.00102f
C15938 CLK.n252 VSS 3.66e-19
C15939 CLK.n253 VSS 0.00935f
C15940 CLK.n254 VSS 0.00927f
C15941 CLK.t39 VSS 9.43e-19
C15942 CLK.t80 VSS 0.00369f
C15943 CLK.n255 VSS 0.00611f
C15944 CLK.n256 VSS 0.0013f
C15945 CLK.n257 VSS 0.00128f
C15946 CLK.n258 VSS 0.00265f
C15947 CLK.n259 VSS 0.0622f
C15948 CLK.n260 VSS 0.367f
C15949 CLK.n261 VSS 0.351f
C15950 CLK.t43 VSS 9.43e-19
C15951 CLK.t85 VSS 0.00369f
C15952 CLK.n262 VSS 0.00611f
C15953 CLK.n263 VSS 0.0013f
C15954 CLK.n264 VSS 0.0611f
C15955 CLK.n265 VSS 0.00265f
C15956 CLK.n266 VSS 0.0645f
C15957 CLK.n267 VSS 0.0153f
C15958 CLK.n268 VSS 0.388f
C15959 CLK.n269 VSS 6.21f
C15960 CLK.n270 VSS 4.51e-19
C15961 CLK.n271 VSS 3.66e-19
C15962 CLK.n272 VSS 0.00146f
C15963 CLK.t75 VSS 0.00447f
C15964 CLK.t13 VSS 0.00294f
C15965 CLK.n273 VSS 0.00789f
C15966 CLK.n274 VSS 0.00103f
C15967 CLK.n275 VSS 7.41e-19
C15968 CLK.n276 VSS 3.7e-19
C15969 CLK.n277 VSS 0.0148f
C15970 CLK.t90 VSS 0.00447f
C15971 CLK.t21 VSS 0.00294f
C15972 CLK.n278 VSS 0.00789f
C15973 CLK.n279 VSS 0.00103f
C15974 CLK.n280 VSS 7.41e-19
C15975 CLK.n281 VSS 0.0146f
C15976 CLK.n282 VSS 0.00854f
C15977 CLK.n283 VSS 3.66e-19
C15978 CLK.n284 VSS 0.00146f
C15979 CLK.t57 VSS 0.00447f
C15980 CLK.t2 VSS 0.00294f
C15981 CLK.n285 VSS 0.00789f
C15982 CLK.n286 VSS 0.00103f
C15983 CLK.n287 VSS 7.41e-19
C15984 CLK.n288 VSS 3.7e-19
C15985 CLK.n289 VSS 0.0138f
C15986 CLK.t44 VSS 0.00232f
C15987 CLK.t36 VSS 0.00414f
C15988 CLK.n290 VSS 0.00788f
C15989 CLK.n291 VSS 0.0253f
C15990 CLK.n292 VSS 0.0304f
C15991 CLK.t69 VSS 0.00447f
C15992 CLK.t8 VSS 0.00294f
C15993 CLK.n293 VSS 0.00789f
C15994 CLK.n294 VSS 0.00103f
C15995 CLK.n295 VSS 7.41e-19
C15996 CLK.n296 VSS 0.00114f
C15997 CLK.n297 VSS 0.00854f
C15998 CLK.n298 VSS 0.00159f
C15999 CLK.n299 VSS 0.00265f
C16000 CLK.t38 VSS 0.00368f
C16001 CLK.t1 VSS 9.53e-19
C16002 CLK.n300 VSS 0.00611f
C16003 CLK.n301 VSS 0.0013f
C16004 CLK.n302 VSS 4.51e-19
C16005 CLK.n303 VSS 9.65e-19
C16006 CLK.n304 VSS 0.0564f
C16007 CLK.n305 VSS 0.0565f
C16008 CLK.n306 VSS 9.65e-19
C16009 CLK.t55 VSS 0.00368f
C16010 CLK.t12 VSS 9.53e-19
C16011 CLK.n307 VSS 0.00611f
C16012 CLK.n308 VSS 0.0013f
C16013 CLK.n309 VSS 0.00159f
C16014 CLK.n310 VSS 0.00125f
C16015 CLK.n311 VSS 6.8f
C16016 CLK.n312 VSS 7.99f
C16017 CLK.n313 VSS 3.58f
C16018 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.t2 VSS 0.025f
C16019 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.t0 VSS 0.0206f
C16020 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.n0 VSS 0.0206f
C16021 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.n1 VSS 0.0494f
C16022 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.t3 VSS 0.0459f
C16023 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.t6 VSS 0.0302f
C16024 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.n2 VSS 0.0814f
C16025 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.t5 VSS 0.0329f
C16026 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.t8 VSS 0.0263f
C16027 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.n3 VSS 0.0764f
C16028 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.n4 VSS 0.606f
C16029 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.t7 VSS 0.0641f
C16030 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.t4 VSS 0.0199f
C16031 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.n5 VSS 0.0675f
C16032 CLK_div_99_mag_0.CLK_div_3_mag_0.Q0.n6 VSS 0.447f
C16033 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n0 VSS 2.13f
C16034 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t0 VSS 0.0354f
C16035 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n1 VSS 0.0354f
C16036 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n2 VSS 0.0755f
C16037 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t2 VSS 0.0797f
C16038 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t5 VSS 0.0507f
C16039 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n3 VSS 0.141f
C16040 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t3 VSS 0.0568f
C16041 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t6 VSS 0.0729f
C16042 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n4 VSS 0.145f
C16043 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t4 VSS 0.0566f
C16044 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.t7 VSS 0.0453f
C16045 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n5 VSS 0.134f
C16046 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n6 VSS 1.21f
C16047 CLK_div_99_mag_0.CLK_div_3_mag_1.JK_FF_mag_1.K.n7 VSS 0.221f
C16048 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t2 VSS 0.02f
C16049 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t0 VSS 0.0165f
C16050 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n0 VSS 0.0165f
C16051 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n1 VSS 0.0396f
C16052 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t9 VSS 0.0367f
C16053 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t3 VSS 0.0242f
C16054 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n2 VSS 0.0652f
C16055 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t4 VSS 0.0263f
C16056 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t10 VSS 0.0211f
C16057 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n3 VSS 0.0612f
C16058 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n4 VSS 0.486f
C16059 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t6 VSS 0.019f
C16060 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t5 VSS 0.034f
C16061 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n5 VSS 0.0648f
C16062 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t8 VSS 0.0263f
C16063 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t7 VSS 0.0211f
C16064 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n6 VSS 0.0612f
C16065 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n7 VSS 0.325f
C16066 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t12 VSS 0.0263f
C16067 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.t11 VSS 0.0211f
C16068 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n8 VSS 0.0612f
C16069 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n9 VSS 0.308f
C16070 CLK_div_105_mag_0.CLK_div_10_mag_1.Q2.n10 VSS 0.15f
C16071 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n0 VSS 0.521f
C16072 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n1 VSS 0.0208f
C16073 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n2 VSS 0.337f
C16074 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n3 VSS 0.0208f
C16075 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n4 VSS 0.141f
C16076 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n5 VSS 0.131f
C16077 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n6 VSS 0.0495f
C16078 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n7 VSS 0.0495f
C16079 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t0 VSS 0.0571f
C16080 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t1 VSS 0.0172f
C16081 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n8 VSS 0.198f
C16082 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t13 VSS 0.0509f
C16083 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t15 VSS 0.0335f
C16084 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n9 VSS 0.09f
C16085 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t9 VSS 0.0509f
C16086 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t12 VSS 0.0335f
C16087 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n10 VSS 0.09f
C16088 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t6 VSS 0.0509f
C16089 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t7 VSS 0.0335f
C16090 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n11 VSS 0.09f
C16091 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t11 VSS 0.0472f
C16092 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t8 VSS 0.0264f
C16093 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n12 VSS 0.0899f
C16094 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n13 VSS 0.288f
C16095 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t3 VSS 0.0509f
C16096 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t4 VSS 0.0335f
C16097 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n14 VSS 0.09f
C16098 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t2 VSS 0.042f
C16099 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t10 VSS 0.0109f
C16100 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n15 VSS 0.0697f
C16101 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n16 VSS 0.671f
C16102 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n17 VSS 0.67f
C16103 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t14 VSS 0.042f
C16104 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.t5 VSS 0.0109f
C16105 CLK_div_108_new_mag_0.CLK_div_3_mag_0.CLK.n18 VSS 0.0697f
C16106 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n0 VSS 0.317f
C16107 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.t2 VSS 0.0207f
C16108 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.t0 VSS 0.0171f
C16109 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n1 VSS 0.0171f
C16110 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n2 VSS 0.047f
C16111 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.t8 VSS 0.0273f
C16112 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.t10 VSS 0.0352f
C16113 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n3 VSS 0.0697f
C16114 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.t7 VSS 0.0218f
C16115 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.t3 VSS 0.0273f
C16116 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n4 VSS 0.0618f
C16117 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.t4 VSS 0.0251f
C16118 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.t5 VSS 0.0381f
C16119 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n5 VSS 0.0676f
C16120 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.t6 VSS 0.0218f
C16121 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.t9 VSS 0.0273f
C16122 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n6 VSS 0.0634f
C16123 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n7 VSS 0.499f
C16124 CLK_div_108_new_mag_0.CLK_div_3_mag_1.Q1.n8 VSS 0.207f
C16125 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t0 VSS 0.0149f
C16126 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n0 VSS 0.0149f
C16127 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n1 VSS 0.0318f
C16128 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t2 VSS 0.0238f
C16129 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t6 VSS 0.0308f
C16130 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n2 VSS 0.0609f
C16131 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t7 VSS 0.0335f
C16132 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t5 VSS 0.0214f
C16133 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n3 VSS 0.0593f
C16134 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n4 VSS 1.14f
C16135 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t4 VSS 0.0238f
C16136 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.t3 VSS 0.0191f
C16137 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n5 VSS 0.0566f
C16138 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n6 VSS 0.381f
C16139 CLK_div_100_mag_0.CLK_div_10_mag_1.JK_FF_mag_2.K.n7 VSS 0.0932f
C16140 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.n0 VSS 0.123f
C16141 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.t4 VSS 0.0265f
C16142 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.t3 VSS 0.0332f
C16143 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.n1 VSS 0.0786f
C16144 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.t6 VSS 0.0297f
C16145 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.t5 VSS 0.0466f
C16146 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.n2 VSS 0.0825f
C16147 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.n3 VSS 0.763f
C16148 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.t0 VSS 0.0207f
C16149 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.n4 VSS 0.0207f
C16150 CLK_div_93_mag_0.CLK_div_31_mag_0.JK_FF_mag_0.QB.n5 VSS 0.0489f
C16151 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.t1 VSS 0.021f
C16152 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.t0 VSS 0.0173f
C16153 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n0 VSS 0.0173f
C16154 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n1 VSS 0.0415f
C16155 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.t7 VSS 0.0276f
C16156 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.t5 VSS 0.0221f
C16157 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n2 VSS 0.0625f
C16158 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.t6 VSS 0.0277f
C16159 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.t10 VSS 0.0355f
C16160 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n3 VSS 0.0706f
C16161 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n4 VSS 0.321f
C16162 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.t4 VSS 0.0385f
C16163 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.t9 VSS 0.0254f
C16164 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n5 VSS 0.0684f
C16165 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.t3 VSS 0.0276f
C16166 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.t8 VSS 0.0221f
C16167 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n6 VSS 0.0642f
C16168 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n7 VSS 0.505f
C16169 CLK_div_99_mag_0.CLK_div_3_mag_1.Q1.n8 VSS 0.209f
C16170 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n0 VSS 0.0877f
C16171 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t7 VSS 0.0189f
C16172 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t6 VSS 0.0237f
C16173 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n1 VSS 0.0561f
C16174 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t8 VSS 0.0333f
C16175 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t5 VSS 0.0212f
C16176 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n2 VSS 0.0588f
C16177 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t3 VSS 0.0306f
C16178 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t4 VSS 0.0235f
C16179 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n3 VSS 0.0604f
C16180 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n4 VSS 1.13f
C16181 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n5 VSS 0.378f
C16182 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t1 VSS 0.0148f
C16183 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n6 VSS 0.0148f
C16184 CLK_div_100_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n7 VSS 0.0349f
C16185 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.t1 VSS 0.021f
C16186 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.t2 VSS 0.0173f
C16187 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n0 VSS 0.0173f
C16188 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n1 VSS 0.0415f
C16189 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.t9 VSS 0.0276f
C16190 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.t8 VSS 0.0221f
C16191 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n2 VSS 0.0625f
C16192 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.t5 VSS 0.0277f
C16193 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.t3 VSS 0.0355f
C16194 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n3 VSS 0.0706f
C16195 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n4 VSS 0.321f
C16196 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.t6 VSS 0.0385f
C16197 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.t10 VSS 0.0254f
C16198 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n5 VSS 0.0684f
C16199 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.t7 VSS 0.0276f
C16200 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.t4 VSS 0.0221f
C16201 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n6 VSS 0.0642f
C16202 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n7 VSS 0.505f
C16203 CLK_div_90_mag_0.CLK_div_3_mag_0.Q1.n8 VSS 0.209f
C16204 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n0 VSS 0.52f
C16205 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n1 VSS 0.328f
C16206 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n2 VSS 0.0208f
C16207 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n3 VSS 0.0494f
C16208 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n4 VSS 0.0494f
C16209 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t1 VSS 0.0172f
C16210 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t0 VSS 0.0571f
C16211 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n5 VSS 0.198f
C16212 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t4 VSS 0.0109f
C16213 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t13 VSS 0.042f
C16214 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n6 VSS 0.0697f
C16215 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t9 VSS 0.0509f
C16216 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t7 VSS 0.0335f
C16217 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n7 VSS 0.09f
C16218 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t2 VSS 0.0509f
C16219 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t14 VSS 0.0335f
C16220 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n8 VSS 0.09f
C16221 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t5 VSS 0.0509f
C16222 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t15 VSS 0.0335f
C16223 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n9 VSS 0.09f
C16224 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t12 VSS 0.0264f
C16225 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t10 VSS 0.0472f
C16226 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n10 VSS 0.0899f
C16227 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n11 VSS 0.288f
C16228 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t8 VSS 0.0509f
C16229 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t6 VSS 0.0335f
C16230 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n12 VSS 0.09f
C16231 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t3 VSS 0.042f
C16232 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.t11 VSS 0.0109f
C16233 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n13 VSS 0.0697f
C16234 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n14 VSS 0.67f
C16235 CLK_div_90_mag_0.CLK_div_3_mag_0.CLK.n15 VSS 0.671f
C16236 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n0 VSS 0.0639f
C16237 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t6 VSS 0.0298f
C16238 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t5 VSS 0.023f
C16239 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n1 VSS 0.059f
C16240 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t8 VSS 0.0207f
C16241 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t7 VSS 0.0324f
C16242 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n2 VSS 0.0574f
C16243 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n3 VSS 1.11f
C16244 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t4 VSS 0.0185f
C16245 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t3 VSS 0.0231f
C16246 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n4 VSS 0.0547f
C16247 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n5 VSS 0.368f
C16248 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t1 VSS 0.0144f
C16249 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n6 VSS 0.0144f
C16250 CLK_div_110_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n7 VSS 0.0308f
C16251 VDD105.t214 VSS 0.00577f
C16252 VDD105.t25 VSS 0.0697f
C16253 VDD105.n0 VSS 0.00577f
C16254 VDD105.t465 VSS 0.00577f
C16255 VDD105.t156 VSS 0.0396f
C16256 VDD105.n1 VSS 0.00577f
C16257 VDD105.n2 VSS 0.00575f
C16258 VDD105.t98 VSS 0.00577f
C16259 VDD105.t295 VSS 0.0697f
C16260 VDD105.n3 VSS 0.00577f
C16261 VDD105.t391 VSS 0.00237f
C16262 VDD105.n4 VSS 0.00237f
C16263 VDD105.n5 VSS 0.00518f
C16264 VDD105.n6 VSS 0.00577f
C16265 VDD105.n7 VSS 0.0337f
C16266 VDD105.t53 VSS 0.0695f
C16267 VDD105.n8 VSS 0.00619f
C16268 VDD105.t248 VSS 0.00237f
C16269 VDD105.n9 VSS 0.00237f
C16270 VDD105.n10 VSS 0.00518f
C16271 VDD105.n11 VSS 0.0329f
C16272 VDD105.n12 VSS 0.0445f
C16273 VDD105.n13 VSS 0.0358f
C16274 VDD105.t247 VSS 0.0393f
C16275 VDD105.t89 VSS 0.0849f
C16276 VDD105.t262 VSS 0.0697f
C16277 VDD105.t289 VSS 0.0849f
C16278 VDD105.t390 VSS 0.0393f
C16279 VDD105.n14 VSS 0.0358f
C16280 VDD105.n15 VSS 0.0179f
C16281 VDD105.n16 VSS 0.0329f
C16282 VDD105.n17 VSS 0.0336f
C16283 VDD105.t226 VSS 0.00577f
C16284 VDD105.n18 VSS 0.00577f
C16285 VDD105.n19 VSS 0.0265f
C16286 VDD105.n20 VSS 0.0286f
C16287 VDD105.n21 VSS 0.02f
C16288 VDD105.n22 VSS 0.0358f
C16289 VDD105.t225 VSS 0.076f
C16290 VDD105.t227 VSS 0.0697f
C16291 VDD105.t97 VSS 0.075f
C16292 VDD105.n23 VSS 0.0358f
C16293 VDD105.n24 VSS 0.02f
C16294 VDD105.n25 VSS 0.051f
C16295 VDD105.t105 VSS 0.00577f
C16296 VDD105.t292 VSS 0.0697f
C16297 VDD105.n26 VSS 0.00577f
C16298 VDD105.t299 VSS 0.00577f
C16299 VDD105.t60 VSS 0.0396f
C16300 VDD105.n27 VSS 0.00577f
C16301 VDD105.n28 VSS 0.0273f
C16302 VDD105.t243 VSS 0.00237f
C16303 VDD105.n29 VSS 0.00237f
C16304 VDD105.n30 VSS 0.00518f
C16305 VDD105.n31 VSS 0.00577f
C16306 VDD105.t234 VSS 0.0695f
C16307 VDD105.n32 VSS 0.0358f
C16308 VDD105.t96 VSS 0.00577f
C16309 VDD105.n33 VSS 0.00575f
C16310 VDD105.t95 VSS 0.0453f
C16311 VDD105.t322 VSS 0.0513f
C16312 VDD105.n34 VSS 0.0838f
C16313 VDD105.n35 VSS 0.00577f
C16314 VDD105.t92 VSS 0.0396f
C16315 VDD105.n36 VSS 0.0358f
C16316 VDD105.t233 VSS 0.00577f
C16317 VDD105.n37 VSS 0.00575f
C16318 VDD105.t232 VSS 0.0453f
C16319 VDD105.t362 VSS 0.0513f
C16320 VDD105.n38 VSS 0.0838f
C16321 VDD105.n39 VSS 0.00577f
C16322 VDD105.t460 VSS 0.0396f
C16323 VDD105.n40 VSS 0.0358f
C16324 VDD105.t100 VSS 0.00577f
C16325 VDD105.n41 VSS 0.00575f
C16326 VDD105.t99 VSS 0.0453f
C16327 VDD105.n42 VSS 0.0532f
C16328 VDD105.t150 VSS 0.0819f
C16329 VDD105.t108 VSS 0.0478f
C16330 VDD105.n43 VSS 0.0813f
C16331 VDD105.n44 VSS 0.00575f
C16332 VDD105.t111 VSS 0.0738f
C16333 VDD105.n45 VSS 0.0444f
C16334 VDD105.t436 VSS 0.00237f
C16335 VDD105.n46 VSS 0.00237f
C16336 VDD105.n47 VSS 0.0052f
C16337 VDD105.n48 VSS 0.0182f
C16338 VDD105.n49 VSS 0.176f
C16339 VDD105.t164 VSS 0.0459f
C16340 VDD105.n50 VSS 0.00577f
C16341 VDD105.t283 VSS 0.00577f
C16342 VDD105.n51 VSS 0.00577f
C16343 VDD105.n52 VSS 0.0286f
C16344 VDD105.t437 VSS 0.0606f
C16345 VDD105.n53 VSS 0.00577f
C16346 VDD105.t429 VSS 0.00575f
C16347 VDD105.t194 VSS 0.00577f
C16348 VDD105.n54 VSS 0.0272f
C16349 VDD105.t193 VSS 0.0314f
C16350 VDD105.t180 VSS 0.041f
C16351 VDD105.n55 VSS 0.00577f
C16352 VDD105.t181 VSS 0.00577f
C16353 VDD105.n56 VSS 0.00577f
C16354 VDD105.n57 VSS 0.0286f
C16355 VDD105.t218 VSS 0.0606f
C16356 VDD105.n58 VSS 0.00577f
C16357 VDD105.t149 VSS 0.00575f
C16358 VDD105.t58 VSS 0.00577f
C16359 VDD105.n59 VSS 0.0272f
C16360 VDD105.t57 VSS 0.0314f
C16361 VDD105.t118 VSS 0.041f
C16362 VDD105.n60 VSS 0.00577f
C16363 VDD105.t119 VSS 0.00577f
C16364 VDD105.n61 VSS 0.00577f
C16365 VDD105.n62 VSS 0.0286f
C16366 VDD105.t80 VSS 0.0606f
C16367 VDD105.n63 VSS 0.00577f
C16368 VDD105.t413 VSS 0.00575f
C16369 VDD105.t3 VSS 0.00577f
C16370 VDD105.n64 VSS 0.0272f
C16371 VDD105.t412 VSS 0.0509f
C16372 VDD105.t430 VSS 0.0395f
C16373 VDD105.t189 VSS 0.00237f
C16374 VDD105.n65 VSS 0.00237f
C16375 VDD105.n66 VSS 0.00518f
C16376 VDD105.t301 VSS 0.00577f
C16377 VDD105.n67 VSS 0.00577f
C16378 VDD105.n68 VSS 0.0286f
C16379 VDD105.t200 VSS 0.0762f
C16380 VDD105.n69 VSS 0.00577f
C16381 VDD105.t321 VSS 0.00577f
C16382 VDD105.n70 VSS 0.00577f
C16383 VDD105.n71 VSS 0.00577f
C16384 VDD105.t365 VSS 0.0751f
C16385 VDD105.n72 VSS 0.0358f
C16386 VDD105.t207 VSS 0.00577f
C16387 VDD105.n73 VSS 0.00577f
C16388 VDD105.t206 VSS 0.0696f
C16389 VDD105.t203 VSS 0.0762f
C16390 VDD105.n74 VSS 0.0358f
C16391 VDD105.t332 VSS 0.00577f
C16392 VDD105.t350 VSS 0.00237f
C16393 VDD105.n75 VSS 0.00237f
C16394 VDD105.n76 VSS 0.00518f
C16395 VDD105.t331 VSS 0.0696f
C16396 VDD105.t349 VSS 0.0849f
C16397 VDD105.t392 VSS 0.0395f
C16398 VDD105.n77 VSS 0.0358f
C16399 VDD105.t278 VSS 0.00577f
C16400 VDD105.t369 VSS 0.00237f
C16401 VDD105.n78 VSS 0.00237f
C16402 VDD105.n79 VSS 0.00518f
C16403 VDD105.t277 VSS 0.0696f
C16404 VDD105.t368 VSS 0.0849f
C16405 VDD105.t414 VSS 0.0395f
C16406 VDD105.t71 VSS 0.0694f
C16407 VDD105.n80 VSS 0.0358f
C16408 VDD105.t72 VSS 0.00539f
C16409 VDD105.t70 VSS 0.00495f
C16410 VDD105.t479 VSS 0.00375f
C16411 VDD105.n81 VSS 0.00967f
C16412 VDD105.n82 VSS 0.00172f
C16413 VDD105.t49 VSS 0.00495f
C16414 VDD105.t490 VSS 0.00375f
C16415 VDD105.n83 VSS 0.00967f
C16416 VDD105.n84 VSS 0.00227f
C16417 VDD105.n85 VSS 0.00117f
C16418 VDD105.n86 VSS 5.93e-19
C16419 VDD105.n87 VSS 0.00529f
C16420 VDD105.n88 VSS 5.7e-19
C16421 VDD105.t38 VSS 0.00481f
C16422 VDD105.n89 VSS 0.00475f
C16423 VDD105.t493 VSS 0.00374f
C16424 VDD105.n90 VSS 0.0016f
C16425 VDD105.n91 VSS 0.00507f
C16426 VDD105.n92 VSS 0.00175f
C16427 VDD105.n93 VSS 0.00144f
C16428 VDD105.t35 VSS 0.00492f
C16429 VDD105.t476 VSS 0.00376f
C16430 VDD105.n94 VSS 0.0097f
C16431 VDD105.n95 VSS 0.00182f
C16432 VDD105.n96 VSS 0.00154f
C16433 VDD105.n97 VSS 5.93e-19
C16434 VDD105.n98 VSS 0.0187f
C16435 VDD105.n99 VSS 0.0725f
C16436 VDD105.n100 VSS 0.106f
C16437 VDD105.t481 VSS 0.00383f
C16438 VDD105.t63 VSS 0.00486f
C16439 VDD105.n101 VSS 0.00968f
C16440 VDD105.n102 VSS 0.00353f
C16441 VDD105.n103 VSS 0.00144f
C16442 VDD105.t485 VSS 0.00376f
C16443 VDD105.t56 VSS 0.00492f
C16444 VDD105.n104 VSS 0.0097f
C16445 VDD105.n105 VSS 0.00189f
C16446 VDD105.n106 VSS 0.00149f
C16447 VDD105.n107 VSS 5.93e-19
C16448 VDD105.n108 VSS 0.0187f
C16449 VDD105.n109 VSS 0.0244f
C16450 VDD105.n110 VSS 0.117f
C16451 VDD105.n111 VSS 0.0494f
C16452 VDD105.n112 VSS 5.6e-19
C16453 VDD105.n113 VSS 0.00464f
C16454 VDD105.n114 VSS 0.0134f
C16455 VDD105.n115 VSS 0.0329f
C16456 VDD105.n116 VSS 0.0329f
C16457 VDD105.n117 VSS 0.0337f
C16458 VDD105.n118 VSS 0.0179f
C16459 VDD105.n119 VSS 0.0329f
C16460 VDD105.n120 VSS 0.0336f
C16461 VDD105.n121 VSS 0.0199f
C16462 VDD105.n122 VSS 0.0286f
C16463 VDD105.n123 VSS 0.0266f
C16464 VDD105.n124 VSS 0.0199f
C16465 VDD105.n125 VSS 0.0544f
C16466 VDD105.n126 VSS 0.0618f
C16467 VDD105.t190 VSS 0.0751f
C16468 VDD105.t320 VSS 0.0696f
C16469 VDD105.n127 VSS 0.0358f
C16470 VDD105.n128 VSS 0.0199f
C16471 VDD105.n129 VSS 0.0266f
C16472 VDD105.n130 VSS 0.0286f
C16473 VDD105.t352 VSS 0.00577f
C16474 VDD105.n131 VSS 0.0266f
C16475 VDD105.n132 VSS 0.0199f
C16476 VDD105.n133 VSS 0.0358f
C16477 VDD105.t351 VSS 0.0696f
C16478 VDD105.t328 VSS 0.0762f
C16479 VDD105.t188 VSS 0.0849f
C16480 VDD105.t300 VSS 0.0696f
C16481 VDD105.n134 VSS 0.0358f
C16482 VDD105.n135 VSS 0.0199f
C16483 VDD105.n136 VSS 0.0252f
C16484 VDD105.n137 VSS 0.0236f
C16485 VDD105.n138 VSS 0.0179f
C16486 VDD105.n139 VSS 0.0358f
C16487 VDD105.t2 VSS 0.0395f
C16488 VDD105.n140 VSS 0.0536f
C16489 VDD105.n141 VSS 0.0181f
C16490 VDD105.n142 VSS 0.00577f
C16491 VDD105.t374 VSS 0.0751f
C16492 VDD105.n143 VSS 0.0358f
C16493 VDD105.t107 VSS 0.00577f
C16494 VDD105.n144 VSS 0.00577f
C16495 VDD105.t106 VSS 0.0696f
C16496 VDD105.t353 VSS 0.0762f
C16497 VDD105.n145 VSS 0.0358f
C16498 VDD105.t24 VSS 0.00577f
C16499 VDD105.t121 VSS 0.00237f
C16500 VDD105.n146 VSS 0.00237f
C16501 VDD105.n147 VSS 0.00518f
C16502 VDD105.t23 VSS 0.0696f
C16503 VDD105.t120 VSS 0.0849f
C16504 VDD105.t387 VSS 0.0395f
C16505 VDD105.n148 VSS 0.0358f
C16506 VDD105.t14 VSS 0.00577f
C16507 VDD105.t378 VSS 0.00237f
C16508 VDD105.n149 VSS 0.00237f
C16509 VDD105.n150 VSS 0.00518f
C16510 VDD105.t13 VSS 0.0696f
C16511 VDD105.t377 VSS 0.0849f
C16512 VDD105.t132 VSS 0.0395f
C16513 VDD105.t64 VSS 0.0694f
C16514 VDD105.n151 VSS 0.0358f
C16515 VDD105.t65 VSS 0.00619f
C16516 VDD105.n152 VSS 0.0444f
C16517 VDD105.n153 VSS 0.0329f
C16518 VDD105.n154 VSS 0.0337f
C16519 VDD105.n155 VSS 0.0179f
C16520 VDD105.n156 VSS 0.0329f
C16521 VDD105.n157 VSS 0.0336f
C16522 VDD105.n158 VSS 0.0199f
C16523 VDD105.n159 VSS 0.0286f
C16524 VDD105.n160 VSS 0.0266f
C16525 VDD105.n161 VSS 0.0199f
C16526 VDD105.n162 VSS 0.0511f
C16527 VDD105.n163 VSS 0.0408f
C16528 VDD105.n164 VSS 0.0293f
C16529 VDD105.t16 VSS 0.00577f
C16530 VDD105.n165 VSS 0.0266f
C16531 VDD105.n166 VSS 0.0199f
C16532 VDD105.n167 VSS 0.0309f
C16533 VDD105.t15 VSS 0.0553f
C16534 VDD105.t356 VSS 0.0606f
C16535 VDD105.n168 VSS 0.0309f
C16536 VDD105.n169 VSS 0.0199f
C16537 VDD105.n170 VSS 0.0266f
C16538 VDD105.n171 VSS 0.0286f
C16539 VDD105.n172 VSS 0.0199f
C16540 VDD105.t84 VSS 0.00237f
C16541 VDD105.n173 VSS 0.00237f
C16542 VDD105.n174 VSS 0.00518f
C16543 VDD105.t147 VSS 0.00577f
C16544 VDD105.n175 VSS 0.00577f
C16545 VDD105.n176 VSS 0.0283f
C16546 VDD105.t12 VSS 0.00575f
C16547 VDD105.n177 VSS 0.0203f
C16548 VDD105.t11 VSS 0.0512f
C16549 VDD105.t135 VSS 0.0455f
C16550 VDD105.n178 VSS 0.00577f
C16551 VDD105.t1 VSS 0.00575f
C16552 VDD105.t434 VSS 0.00577f
C16553 VDD105.n179 VSS 0.0269f
C16554 VDD105.t0 VSS 0.0512f
C16555 VDD105.t384 VSS 0.0455f
C16556 VDD105.n180 VSS 0.00577f
C16557 VDD105.t86 VSS 0.00575f
C16558 VDD105.t319 VSS 0.00585f
C16559 VDD105.n181 VSS 0.0313f
C16560 VDD105.t195 VSS 0.0738f
C16561 VDD105.t196 VSS 0.00575f
C16562 VDD105.n182 VSS 0.0259f
C16563 VDD105.t46 VSS 0.054f
C16564 VDD105.t88 VSS 0.0224f
C16565 VDD105.n183 VSS 0.00577f
C16566 VDD105.n184 VSS 0.00602f
C16567 VDD105.t304 VSS 0.19f
C16568 VDD105.t463 VSS 0.068f
C16569 VDD105.t87 VSS 0.0847f
C16570 VDD105.n185 VSS 0.0731f
C16571 VDD105.n186 VSS 0.00996f
C16572 VDD105.n187 VSS 0.0253f
C16573 VDD105.n188 VSS 0.0271f
C16574 VDD105.n189 VSS 0.0167f
C16575 VDD105.n190 VSS 0.0563f
C16576 VDD105.t128 VSS 0.076f
C16577 VDD105.n191 VSS 0.00577f
C16578 VDD105.t303 VSS 0.00237f
C16579 VDD105.n192 VSS 0.00237f
C16580 VDD105.n193 VSS 0.0052f
C16581 VDD105.n194 VSS 0.0182f
C16582 VDD105.n195 VSS 0.0252f
C16583 VDD105.t129 VSS 0.00577f
C16584 VDD105.n196 VSS 0.00577f
C16585 VDD105.t268 VSS 0.0697f
C16586 VDD105.n197 VSS 0.0358f
C16587 VDD105.t373 VSS 0.00577f
C16588 VDD105.n198 VSS 0.00577f
C16589 VDD105.t372 VSS 0.076f
C16590 VDD105.t271 VSS 0.0697f
C16591 VDD105.t175 VSS 0.075f
C16592 VDD105.n199 VSS 0.0358f
C16593 VDD105.t176 VSS 0.00577f
C16594 VDD105.n200 VSS 0.00575f
C16595 VDD105.t455 VSS 0.051f
C16596 VDD105.n201 VSS 0.0536f
C16597 VDD105.n202 VSS 0.00577f
C16598 VDD105.t210 VSS 0.0396f
C16599 VDD105.n203 VSS 0.0358f
C16600 VDD105.t449 VSS 0.00237f
C16601 VDD105.n204 VSS 0.00237f
C16602 VDD105.n205 VSS 0.00518f
C16603 VDD105.n206 VSS 0.00577f
C16604 VDD105.t448 VSS 0.0393f
C16605 VDD105.t249 VSS 0.0849f
C16606 VDD105.t279 VSS 0.0697f
C16607 VDD105.n207 VSS 0.0358f
C16608 VDD105.t261 VSS 0.00577f
C16609 VDD105.n208 VSS 0.00577f
C16610 VDD105.t260 VSS 0.076f
C16611 VDD105.t312 VSS 0.0697f
C16612 VDD105.n209 VSS 0.0358f
C16613 VDD105.t117 VSS 0.00577f
C16614 VDD105.n210 VSS 0.00577f
C16615 VDD105.t116 VSS 0.076f
C16616 VDD105.t315 VSS 0.0697f
C16617 VDD105.t252 VSS 0.075f
C16618 VDD105.n211 VSS 0.0358f
C16619 VDD105.t253 VSS 0.00577f
C16620 VDD105.n212 VSS 0.00575f
C16621 VDD105.t244 VSS 0.051f
C16622 VDD105.n213 VSS 0.0536f
C16623 VDD105.n214 VSS 0.0181f
C16624 VDD105.t241 VSS 0.00577f
C16625 VDD105.t257 VSS 0.0697f
C16626 VDD105.n215 VSS 0.00577f
C16627 VDD105.t396 VSS 0.00237f
C16628 VDD105.n216 VSS 0.00237f
C16629 VDD105.n217 VSS 0.00518f
C16630 VDD105.n218 VSS 0.00577f
C16631 VDD105.n219 VSS 0.0337f
C16632 VDD105.t67 VSS 0.0695f
C16633 VDD105.n220 VSS 0.00619f
C16634 VDD105.t451 VSS 0.00237f
C16635 VDD105.n221 VSS 0.00237f
C16636 VDD105.n222 VSS 0.00518f
C16637 VDD105.n223 VSS 0.0329f
C16638 VDD105.n224 VSS 0.0445f
C16639 VDD105.n225 VSS 0.0358f
C16640 VDD105.t450 VSS 0.0393f
C16641 VDD105.t237 VSS 0.0849f
C16642 VDD105.t325 VSS 0.0697f
C16643 VDD105.t309 VSS 0.0849f
C16644 VDD105.t395 VSS 0.0393f
C16645 VDD105.n226 VSS 0.0358f
C16646 VDD105.n227 VSS 0.0179f
C16647 VDD105.n228 VSS 0.0329f
C16648 VDD105.n229 VSS 0.0336f
C16649 VDD105.t115 VSS 0.00577f
C16650 VDD105.n230 VSS 0.00577f
C16651 VDD105.n231 VSS 0.0265f
C16652 VDD105.n232 VSS 0.0286f
C16653 VDD105.n233 VSS 0.02f
C16654 VDD105.n234 VSS 0.0358f
C16655 VDD105.t114 VSS 0.076f
C16656 VDD105.t254 VSS 0.0697f
C16657 VDD105.t240 VSS 0.075f
C16658 VDD105.n235 VSS 0.0358f
C16659 VDD105.n236 VSS 0.02f
C16660 VDD105.n237 VSS 0.051f
C16661 VDD105.n238 VSS 0.0407f
C16662 VDD105.n239 VSS 0.0293f
C16663 VDD105.n240 VSS 0.02f
C16664 VDD105.n241 VSS 0.0265f
C16665 VDD105.n242 VSS 0.0286f
C16666 VDD105.n243 VSS 0.02f
C16667 VDD105.n244 VSS 0.0265f
C16668 VDD105.n245 VSS 0.0286f
C16669 VDD105.n246 VSS 0.02f
C16670 VDD105.n247 VSS 0.0252f
C16671 VDD105.n248 VSS 0.0236f
C16672 VDD105.n249 VSS 0.0179f
C16673 VDD105.n250 VSS 0.0273f
C16674 VDD105.n251 VSS 0.0177f
C16675 VDD105.t447 VSS 0.00577f
C16676 VDD105.t125 VSS 0.0697f
C16677 VDD105.n252 VSS 0.00577f
C16678 VDD105.t398 VSS 0.00237f
C16679 VDD105.n253 VSS 0.00237f
C16680 VDD105.n254 VSS 0.00518f
C16681 VDD105.n255 VSS 0.00577f
C16682 VDD105.n256 VSS 0.0337f
C16683 VDD105.t74 VSS 0.0695f
C16684 VDD105.n257 VSS 0.00619f
C16685 VDD105.t308 VSS 0.00237f
C16686 VDD105.n258 VSS 0.00237f
C16687 VDD105.n259 VSS 0.00518f
C16688 VDD105.n260 VSS 0.0329f
C16689 VDD105.n261 VSS 0.0445f
C16690 VDD105.n262 VSS 0.0358f
C16691 VDD105.t307 VSS 0.0393f
C16692 VDD105.t452 VSS 0.0849f
C16693 VDD105.t274 VSS 0.0697f
C16694 VDD105.t265 VSS 0.0849f
C16695 VDD105.t397 VSS 0.0393f
C16696 VDD105.n263 VSS 0.0358f
C16697 VDD105.n264 VSS 0.0179f
C16698 VDD105.n265 VSS 0.0329f
C16699 VDD105.n266 VSS 0.0336f
C16700 VDD105.t371 VSS 0.00577f
C16701 VDD105.n267 VSS 0.00577f
C16702 VDD105.n268 VSS 0.0265f
C16703 VDD105.n269 VSS 0.0286f
C16704 VDD105.n270 VSS 0.02f
C16705 VDD105.n271 VSS 0.0358f
C16706 VDD105.t370 VSS 0.076f
C16707 VDD105.t122 VSS 0.0697f
C16708 VDD105.t446 VSS 0.075f
C16709 VDD105.n272 VSS 0.0358f
C16710 VDD105.n273 VSS 0.02f
C16711 VDD105.n274 VSS 0.051f
C16712 VDD105.n275 VSS 0.0362f
C16713 VDD105.n276 VSS 0.0293f
C16714 VDD105.n277 VSS 0.02f
C16715 VDD105.n278 VSS 0.0265f
C16716 VDD105.n279 VSS 0.0286f
C16717 VDD105.n280 VSS 0.02f
C16718 VDD105.n281 VSS 0.0265f
C16719 VDD105.n282 VSS 0.0286f
C16720 VDD105.n283 VSS 0.02f
C16721 VDD105.n284 VSS 0.0358f
C16722 VDD105.t359 VSS 0.0697f
C16723 VDD105.t177 VSS 0.0849f
C16724 VDD105.t302 VSS 0.0366f
C16725 VDD105.n285 VSS 0.0559f
C16726 VDD105.n286 VSS 0.0444f
C16727 VDD105.n287 VSS 0.0273f
C16728 VDD105.n288 VSS 0.019f
C16729 VDD105.n289 VSS 0.0813f
C16730 VDD105.t318 VSS 0.048f
C16731 VDD105.t85 VSS 0.0815f
C16732 VDD105.n290 VSS 0.0532f
C16733 VDD105.n291 VSS 0.0203f
C16734 VDD105.n292 VSS 0.0283f
C16735 VDD105.n293 VSS 0.0202f
C16736 VDD105.n294 VSS 0.0358f
C16737 VDD105.t433 VSS 0.0395f
C16738 VDD105.n295 VSS 0.0838f
C16739 VDD105.n296 VSS 0.0203f
C16740 VDD105.n297 VSS 0.0283f
C16741 VDD105.t380 VSS 0.00577f
C16742 VDD105.n298 VSS 0.0269f
C16743 VDD105.n299 VSS 0.0202f
C16744 VDD105.n300 VSS 0.0358f
C16745 VDD105.t379 VSS 0.0395f
C16746 VDD105.n301 VSS 0.0838f
C16747 VDD105.t381 VSS 0.0455f
C16748 VDD105.t146 VSS 0.0694f
C16749 VDD105.n302 VSS 0.0358f
C16750 VDD105.n303 VSS 0.0202f
C16751 VDD105.n304 VSS 0.0519f
C16752 VDD105.t408 VSS 0.00577f
C16753 VDD105.n305 VSS 0.0189f
C16754 VDD105.n306 VSS 0.029f
C16755 VDD105.n307 VSS 0.0236f
C16756 VDD105.n308 VSS 0.0179f
C16757 VDD105.n309 VSS 0.0309f
C16758 VDD105.t143 VSS 0.0314f
C16759 VDD105.t83 VSS 0.0676f
C16760 VDD105.t407 VSS 0.0553f
C16761 VDD105.n310 VSS 0.0309f
C16762 VDD105.t20 VSS 0.0266f
C16763 VDD105.n311 VSS 0.16f
C16764 VDD105.n312 VSS 0.0884f
C16765 VDD105.t148 VSS 0.0636f
C16766 VDD105.n313 VSS 0.0181f
C16767 VDD105.n314 VSS 0.00577f
C16768 VDD105.t138 VSS 0.0751f
C16769 VDD105.n315 VSS 0.0358f
C16770 VDD105.t342 VSS 0.00577f
C16771 VDD105.n316 VSS 0.00577f
C16772 VDD105.t341 VSS 0.0696f
C16773 VDD105.t338 VSS 0.0762f
C16774 VDD105.n317 VSS 0.0358f
C16775 VDD105.t8 VSS 0.00577f
C16776 VDD105.t183 VSS 0.00237f
C16777 VDD105.n318 VSS 0.00237f
C16778 VDD105.n319 VSS 0.00518f
C16779 VDD105.t7 VSS 0.0696f
C16780 VDD105.t182 VSS 0.0849f
C16781 VDD105.t402 VSS 0.0395f
C16782 VDD105.n320 VSS 0.0358f
C16783 VDD105.t209 VSS 0.00577f
C16784 VDD105.t142 VSS 0.00237f
C16785 VDD105.n321 VSS 0.00237f
C16786 VDD105.n322 VSS 0.00518f
C16787 VDD105.t208 VSS 0.0696f
C16788 VDD105.t141 VSS 0.0849f
C16789 VDD105.t423 VSS 0.0395f
C16790 VDD105.t50 VSS 0.0694f
C16791 VDD105.n323 VSS 0.0358f
C16792 VDD105.t51 VSS 0.00619f
C16793 VDD105.n324 VSS 0.0444f
C16794 VDD105.n325 VSS 0.0329f
C16795 VDD105.n326 VSS 0.0337f
C16796 VDD105.n327 VSS 0.0179f
C16797 VDD105.n328 VSS 0.0329f
C16798 VDD105.n329 VSS 0.0336f
C16799 VDD105.n330 VSS 0.0199f
C16800 VDD105.n331 VSS 0.0286f
C16801 VDD105.n332 VSS 0.0266f
C16802 VDD105.n333 VSS 0.0199f
C16803 VDD105.n334 VSS 0.0511f
C16804 VDD105.n335 VSS 0.0408f
C16805 VDD105.n336 VSS 0.0293f
C16806 VDD105.t10 VSS 0.00577f
C16807 VDD105.n337 VSS 0.0266f
C16808 VDD105.n338 VSS 0.0199f
C16809 VDD105.n339 VSS 0.0309f
C16810 VDD105.t9 VSS 0.0553f
C16811 VDD105.t335 VSS 0.0606f
C16812 VDD105.n340 VSS 0.0309f
C16813 VDD105.n341 VSS 0.0199f
C16814 VDD105.n342 VSS 0.0266f
C16815 VDD105.n343 VSS 0.0286f
C16816 VDD105.n344 VSS 0.0199f
C16817 VDD105.t222 VSS 0.00237f
C16818 VDD105.n345 VSS 0.00237f
C16819 VDD105.n346 VSS 0.00518f
C16820 VDD105.t185 VSS 0.00577f
C16821 VDD105.n347 VSS 0.0252f
C16822 VDD105.n348 VSS 0.0236f
C16823 VDD105.n349 VSS 0.0179f
C16824 VDD105.n350 VSS 0.0309f
C16825 VDD105.t420 VSS 0.0314f
C16826 VDD105.t221 VSS 0.0676f
C16827 VDD105.t184 VSS 0.0553f
C16828 VDD105.n351 VSS 0.0309f
C16829 VDD105.t4 VSS 0.0266f
C16830 VDD105.n352 VSS 0.16f
C16831 VDD105.n353 VSS 0.0884f
C16832 VDD105.t428 VSS 0.0636f
C16833 VDD105.n354 VSS 0.0177f
C16834 VDD105.n355 VSS 0.00577f
C16835 VDD105.t417 VSS 0.0751f
C16836 VDD105.n356 VSS 0.0358f
C16837 VDD105.t231 VSS 0.00577f
C16838 VDD105.n357 VSS 0.00577f
C16839 VDD105.t230 VSS 0.0696f
C16840 VDD105.t170 VSS 0.0762f
C16841 VDD105.n358 VSS 0.0358f
C16842 VDD105.t163 VSS 0.00577f
C16843 VDD105.t285 VSS 0.00237f
C16844 VDD105.n359 VSS 0.00237f
C16845 VDD105.n360 VSS 0.00518f
C16846 VDD105.t162 VSS 0.0696f
C16847 VDD105.t284 VSS 0.0849f
C16848 VDD105.t399 VSS 0.0395f
C16849 VDD105.n361 VSS 0.0358f
C16850 VDD105.t187 VSS 0.00577f
C16851 VDD105.t427 VSS 0.00237f
C16852 VDD105.n362 VSS 0.00237f
C16853 VDD105.n363 VSS 0.00518f
C16854 VDD105.t186 VSS 0.0696f
C16855 VDD105.t426 VSS 0.0849f
C16856 VDD105.t470 VSS 0.0395f
C16857 VDD105.t39 VSS 0.0694f
C16858 VDD105.n364 VSS 0.0358f
C16859 VDD105.t40 VSS 0.00619f
C16860 VDD105.n365 VSS 0.0444f
C16861 VDD105.n366 VSS 0.0329f
C16862 VDD105.n367 VSS 0.0337f
C16863 VDD105.n368 VSS 0.0179f
C16864 VDD105.n369 VSS 0.0329f
C16865 VDD105.n370 VSS 0.0336f
C16866 VDD105.n371 VSS 0.0199f
C16867 VDD105.n372 VSS 0.0286f
C16868 VDD105.n373 VSS 0.0266f
C16869 VDD105.n374 VSS 0.0199f
C16870 VDD105.n375 VSS 0.0511f
C16871 VDD105.n376 VSS 0.0363f
C16872 VDD105.n377 VSS 0.0293f
C16873 VDD105.t174 VSS 0.00577f
C16874 VDD105.n378 VSS 0.0266f
C16875 VDD105.n379 VSS 0.0199f
C16876 VDD105.n380 VSS 0.0309f
C16877 VDD105.t173 VSS 0.0553f
C16878 VDD105.t167 VSS 0.0606f
C16879 VDD105.t282 VSS 0.0217f
C16880 VDD105.n381 VSS 0.0309f
C16881 VDD105.n382 VSS 0.0199f
C16882 VDD105.n383 VSS 0.0266f
C16883 VDD105.n384 VSS 0.0286f
C16884 VDD105.t334 VSS 0.00577f
C16885 VDD105.n385 VSS 0.0252f
C16886 VDD105.n386 VSS 0.0199f
C16887 VDD105.n387 VSS 0.0309f
C16888 VDD105.t333 VSS 0.0553f
C16889 VDD105.t435 VSS 0.0676f
C16890 VDD105.t473 VSS 0.0291f
C16891 VDD105.n388 VSS 0.0578f
C16892 VDD105.n389 VSS 0.0563f
C16893 VDD105.n390 VSS 0.0224f
C16894 VDD105.t37 VSS 0.00577f
C16895 VDD105.t36 VSS 0.0537f
C16896 VDD105.t286 VSS 0.0847f
C16897 VDD105.n391 VSS 0.0731f
C16898 VDD105.t440 VSS 0.068f
C16899 VDD105.t348 VSS 0.19f
C16900 VDD105.t469 VSS 0.00602f
C16901 VDD105.n392 VSS 0.00988f
C16902 VDD105.n393 VSS 0.0253f
C16903 VDD105.n394 VSS 0.0271f
C16904 VDD105.n395 VSS 0.0168f
C16905 VDD105.n396 VSS 0.0259f
C16906 VDD105.n397 VSS 0.0273f
C16907 VDD105.n398 VSS 0.019f
C16908 VDD105.n399 VSS 0.00585f
C16909 VDD105.n400 VSS 0.0313f
C16910 VDD105.n401 VSS 0.0203f
C16911 VDD105.n402 VSS 0.0283f
C16912 VDD105.n403 VSS 0.0202f
C16913 VDD105.n404 VSS 0.0269f
C16914 VDD105.n405 VSS 0.0203f
C16915 VDD105.n406 VSS 0.0283f
C16916 VDD105.n407 VSS 0.0202f
C16917 VDD105.n408 VSS 0.0269f
C16918 VDD105.n409 VSS 0.0203f
C16919 VDD105.n410 VSS 0.0283f
C16920 VDD105.n411 VSS 0.0202f
C16921 VDD105.n412 VSS 0.0726f
C16922 VDD105.n413 VSS 0.00577f
C16923 VDD105.n414 VSS 0.0189f
C16924 VDD105.n415 VSS 0.0611f
C16925 VDD105.n416 VSS 0.0236f
C16926 VDD105.n417 VSS 0.0179f
C16927 VDD105.n418 VSS 0.0358f
C16928 VDD105.t242 VSS 0.0393f
C16929 VDD105.t101 VSS 0.0849f
C16930 VDD105.t153 VSS 0.0697f
C16931 VDD105.t298 VSS 0.076f
C16932 VDD105.n419 VSS 0.0358f
C16933 VDD105.n420 VSS 0.02f
C16934 VDD105.n421 VSS 0.0286f
C16935 VDD105.n422 VSS 0.0265f
C16936 VDD105.t224 VSS 0.00577f
C16937 VDD105.n423 VSS 0.00577f
C16938 VDD105.n424 VSS 0.0265f
C16939 VDD105.n425 VSS 0.0286f
C16940 VDD105.n426 VSS 0.02f
C16941 VDD105.n427 VSS 0.0358f
C16942 VDD105.t223 VSS 0.076f
C16943 VDD105.t17 VSS 0.0697f
C16944 VDD105.t104 VSS 0.075f
C16945 VDD105.n428 VSS 0.0358f
C16946 VDD105.n429 VSS 0.02f
C16947 VDD105.n430 VSS 0.0293f
C16948 VDD105.n431 VSS 0.0407f
C16949 VDD105.n432 VSS 0.0181f
C16950 VDD105.t441 VSS 0.051f
C16951 VDD105.n433 VSS 0.0536f
C16952 VDD105.n434 VSS 0.0273f
C16953 VDD105.t459 VSS 0.00237f
C16954 VDD105.n435 VSS 0.00237f
C16955 VDD105.n436 VSS 0.00518f
C16956 VDD105.n437 VSS 0.00577f
C16957 VDD105.n438 VSS 0.0252f
C16958 VDD105.n439 VSS 0.0236f
C16959 VDD105.n440 VSS 0.0179f
C16960 VDD105.n441 VSS 0.0358f
C16961 VDD105.t458 VSS 0.0393f
C16962 VDD105.t215 VSS 0.0849f
C16963 VDD105.t159 VSS 0.0697f
C16964 VDD105.t464 VSS 0.076f
C16965 VDD105.n442 VSS 0.0358f
C16966 VDD105.n443 VSS 0.02f
C16967 VDD105.n444 VSS 0.0286f
C16968 VDD105.n445 VSS 0.0265f
C16969 VDD105.t34 VSS 0.00577f
C16970 VDD105.n446 VSS 0.00577f
C16971 VDD105.n447 VSS 0.0265f
C16972 VDD105.n448 VSS 0.0286f
C16973 VDD105.n449 VSS 0.02f
C16974 VDD105.n450 VSS 0.0358f
C16975 VDD105.t33 VSS 0.076f
C16976 VDD105.t77 VSS 0.0697f
C16977 VDD105.t213 VSS 0.075f
C16978 VDD105.n451 VSS 0.0358f
C16979 VDD105.n452 VSS 0.02f
C16980 VDD105.n453 VSS 0.0278f
C16981 VDD105.t347 VSS 0.00577f
C16982 VDD105.t466 VSS 0.0697f
C16983 VDD105.n454 VSS 0.00577f
C16984 VDD105.t406 VSS 0.00237f
C16985 VDD105.n455 VSS 0.00237f
C16986 VDD105.n456 VSS 0.00518f
C16987 VDD105.n457 VSS 0.00577f
C16988 VDD105.n458 VSS 0.0337f
C16989 VDD105.t42 VSS 0.0695f
C16990 VDD105.n459 VSS 0.00172f
C16991 VDD105.n460 VSS 0.00119f
C16992 VDD105.t488 VSS 0.00375f
C16993 VDD105.t66 VSS 0.00495f
C16994 VDD105.n461 VSS 0.00967f
C16995 VDD105.n462 VSS 0.00225f
C16996 VDD105.n463 VSS 5.93e-19
C16997 VDD105.n464 VSS 0.00529f
C16998 VDD105.n465 VSS 0.00144f
C16999 VDD105.n466 VSS 0.00154f
C17000 VDD105.t45 VSS 0.00492f
C17001 VDD105.t492 VSS 0.00376f
C17002 VDD105.n467 VSS 0.0097f
C17003 VDD105.n468 VSS 0.00182f
C17004 VDD105.n469 VSS 5.93e-19
C17005 VDD105.n470 VSS 0.0187f
C17006 VDD105.n471 VSS 0.00164f
C17007 VDD105.t477 VSS 0.00375f
C17008 VDD105.n472 VSS 0.00515f
C17009 VDD105.t73 VSS 0.00485f
C17010 VDD105.n473 VSS 0.00461f
C17011 VDD105.n474 VSS 0.00227f
C17012 VDD105.n475 VSS 0.0725f
C17013 VDD105.n476 VSS 0.106f
C17014 VDD105.n477 VSS 0.00144f
C17015 VDD105.n478 VSS 0.00149f
C17016 VDD105.t59 VSS 0.00492f
C17017 VDD105.t484 VSS 0.00376f
C17018 VDD105.n479 VSS 0.0097f
C17019 VDD105.n480 VSS 0.00189f
C17020 VDD105.n481 VSS 5.93e-19
C17021 VDD105.n482 VSS 0.0187f
C17022 VDD105.t487 VSS 0.00384f
C17023 VDD105.t52 VSS 0.00485f
C17024 VDD105.n483 VSS 0.00968f
C17025 VDD105.n484 VSS 0.00351f
C17026 VDD105.n485 VSS 0.0245f
C17027 VDD105.n486 VSS 0.117f
C17028 VDD105.t483 VSS 0.00375f
C17029 VDD105.t41 VSS 0.00495f
C17030 VDD105.n487 VSS 0.00967f
C17031 VDD105.n488 VSS 0.0486f
C17032 VDD105.n489 VSS 0.0035f
C17033 VDD105.n490 VSS 0.00539f
C17034 VDD105.n491 VSS 0.0151f
C17035 VDD105.t445 VSS 0.00237f
C17036 VDD105.n492 VSS 0.00237f
C17037 VDD105.n493 VSS 0.00518f
C17038 VDD105.n494 VSS 0.0329f
C17039 VDD105.n495 VSS 0.033f
C17040 VDD105.n496 VSS 0.0358f
C17041 VDD105.t444 VSS 0.0393f
C17042 VDD105.t343 VSS 0.0849f
C17043 VDD105.t197 VSS 0.0697f
C17044 VDD105.t28 VSS 0.0849f
C17045 VDD105.t405 VSS 0.0393f
C17046 VDD105.n497 VSS 0.0358f
C17047 VDD105.n498 VSS 0.0179f
C17048 VDD105.n499 VSS 0.0329f
C17049 VDD105.n500 VSS 0.0336f
C17050 VDD105.t32 VSS 0.00577f
C17051 VDD105.n501 VSS 0.00577f
C17052 VDD105.n502 VSS 0.0265f
C17053 VDD105.n503 VSS 0.0286f
C17054 VDD105.n504 VSS 0.02f
C17055 VDD105.n505 VSS 0.0358f
C17056 VDD105.t31 VSS 0.076f
C17057 VDD105.t409 VSS 0.0697f
C17058 VDD105.t346 VSS 0.075f
C17059 VDD105.n506 VSS 0.0358f
C17060 VDD105.n507 VSS 0.02f
C17061 VDD105.n508 VSS 0.05f
C17062 VDD105.n509 VSS 0.0663f
C17063 VDD105.n510 VSS 0.00129f
C17064 VDD105.n511 VSS 0.00577f
C17065 VDD105.n512 VSS 0.0232f
C17066 VDD108.t314 VSS 0.00797f
C17067 VDD108.t19 VSS 0.00634f
C17068 VDD108.t253 VSS 0.0837f
C17069 VDD108.n0 VSS 0.00633f
C17070 VDD108.t259 VSS 0.00634f
C17071 VDD108.n1 VSS 0.00633f
C17072 VDD108.n2 VSS 0.115f
C17073 VDD108.t428 VSS 0.0825f
C17074 VDD108.n3 VSS 0.00633f
C17075 VDD108.n4 VSS 0.00633f
C17076 VDD108.t421 VSS 0.0825f
C17077 VDD108.n5 VSS 0.0393f
C17078 VDD108.t250 VSS 0.00634f
C17079 VDD108.n6 VSS 0.00633f
C17080 VDD108.t249 VSS 0.0764f
C17081 VDD108.t431 VSS 0.0837f
C17082 VDD108.n7 VSS 0.0393f
C17083 VDD108.t252 VSS 0.00634f
C17084 VDD108.t257 VSS 0.00261f
C17085 VDD108.n8 VSS 0.00261f
C17086 VDD108.n9 VSS 0.00569f
C17087 VDD108.t251 VSS 0.0764f
C17088 VDD108.t256 VSS 0.0933f
C17089 VDD108.t341 VSS 0.0433f
C17090 VDD108.n10 VSS 0.0393f
C17091 VDD108.t330 VSS 0.00634f
C17092 VDD108.t425 VSS 0.00261f
C17093 VDD108.n11 VSS 0.00261f
C17094 VDD108.n12 VSS 0.00569f
C17095 VDD108.t329 VSS 0.0764f
C17096 VDD108.t424 VSS 0.0933f
C17097 VDD108.t310 VSS 0.0433f
C17098 VDD108.t31 VSS 0.0762f
C17099 VDD108.n13 VSS 0.0393f
C17100 VDD108.t32 VSS 0.00634f
C17101 VDD108.t17 VSS 0.00544f
C17102 VDD108.t461 VSS 0.00412f
C17103 VDD108.n14 VSS 0.0109f
C17104 VDD108.t30 VSS 0.00544f
C17105 VDD108.t456 VSS 0.00412f
C17106 VDD108.n15 VSS 0.0106f
C17107 VDD108.n16 VSS 0.00368f
C17108 VDD108.n17 VSS 0.0444f
C17109 VDD108.n18 VSS 0.0294f
C17110 VDD108.n19 VSS 0.0197f
C17111 VDD108.n20 VSS 0.0361f
C17112 VDD108.n21 VSS 0.037f
C17113 VDD108.n22 VSS 0.0197f
C17114 VDD108.n23 VSS 0.0361f
C17115 VDD108.n24 VSS 0.0369f
C17116 VDD108.n25 VSS 0.0219f
C17117 VDD108.n26 VSS 0.0314f
C17118 VDD108.n27 VSS 0.0292f
C17119 VDD108.n28 VSS 0.0219f
C17120 VDD108.n29 VSS 0.055f
C17121 VDD108.t417 VSS 0.00797f
C17122 VDD108.n30 VSS 0.0924f
C17123 VDD108.t416 VSS 0.0559f
C17124 VDD108.t418 VSS 0.0433f
C17125 VDD108.t197 VSS 0.00261f
C17126 VDD108.n31 VSS 0.00261f
C17127 VDD108.n32 VSS 0.00569f
C17128 VDD108.t199 VSS 0.00634f
C17129 VDD108.n33 VSS 0.00633f
C17130 VDD108.n34 VSS 0.115f
C17131 VDD108.t282 VSS 0.0837f
C17132 VDD108.n35 VSS 0.00633f
C17133 VDD108.t304 VSS 0.00634f
C17134 VDD108.n36 VSS 0.00633f
C17135 VDD108.n37 VSS 0.00633f
C17136 VDD108.t209 VSS 0.0825f
C17137 VDD108.n38 VSS 0.0393f
C17138 VDD108.t61 VSS 0.00634f
C17139 VDD108.n39 VSS 0.00633f
C17140 VDD108.t60 VSS 0.0764f
C17141 VDD108.t285 VSS 0.0837f
C17142 VDD108.n40 VSS 0.0393f
C17143 VDD108.t205 VSS 0.00634f
C17144 VDD108.t203 VSS 0.00261f
C17145 VDD108.n41 VSS 0.00261f
C17146 VDD108.n42 VSS 0.00569f
C17147 VDD108.t204 VSS 0.0764f
C17148 VDD108.t202 VSS 0.0933f
C17149 VDD108.t344 VSS 0.0433f
C17150 VDD108.n43 VSS 0.0393f
C17151 VDD108.t56 VSS 0.00634f
C17152 VDD108.t213 VSS 0.00261f
C17153 VDD108.n44 VSS 0.00261f
C17154 VDD108.n45 VSS 0.00569f
C17155 VDD108.t55 VSS 0.0764f
C17156 VDD108.t212 VSS 0.0933f
C17157 VDD108.t413 VSS 0.0433f
C17158 VDD108.t24 VSS 0.0762f
C17159 VDD108.n46 VSS 0.0393f
C17160 VDD108.t25 VSS 0.00634f
C17161 VDD108.t10 VSS 0.00544f
C17162 VDD108.t463 VSS 0.00412f
C17163 VDD108.n47 VSS 0.0107f
C17164 VDD108.n48 VSS 0.00875f
C17165 VDD108.t23 VSS 0.00544f
C17166 VDD108.t458 VSS 0.00412f
C17167 VDD108.n49 VSS 0.0107f
C17168 VDD108.n50 VSS 0.0488f
C17169 VDD108.n51 VSS 0.0295f
C17170 VDD108.n52 VSS 0.0197f
C17171 VDD108.n53 VSS 0.0361f
C17172 VDD108.n54 VSS 0.037f
C17173 VDD108.n55 VSS 0.0197f
C17174 VDD108.n56 VSS 0.0361f
C17175 VDD108.n57 VSS 0.0369f
C17176 VDD108.n58 VSS 0.0219f
C17177 VDD108.n59 VSS 0.0314f
C17178 VDD108.n60 VSS 0.0292f
C17179 VDD108.n61 VSS 0.0219f
C17180 VDD108.n62 VSS 0.055f
C17181 VDD108.n63 VSS 0.00631f
C17182 VDD108.t446 VSS 0.0559f
C17183 VDD108.n64 VSS 0.0588f
C17184 VDD108.n65 VSS 0.00632f
C17185 VDD108.t399 VSS 0.0435f
C17186 VDD108.n66 VSS 0.0393f
C17187 VDD108.t453 VSS 0.00261f
C17188 VDD108.n67 VSS 0.00261f
C17189 VDD108.n68 VSS 0.00567f
C17190 VDD108.n69 VSS 0.00632f
C17191 VDD108.t452 VSS 0.0432f
C17192 VDD108.t123 VSS 0.0933f
C17193 VDD108.t126 VSS 0.0766f
C17194 VDD108.n70 VSS 0.0393f
C17195 VDD108.t139 VSS 0.00632f
C17196 VDD108.n71 VSS 0.00632f
C17197 VDD108.t138 VSS 0.0835f
C17198 VDD108.t129 VSS 0.0766f
C17199 VDD108.n72 VSS 0.0393f
C17200 VDD108.t245 VSS 0.00632f
C17201 VDD108.n73 VSS 0.00632f
C17202 VDD108.t244 VSS 0.0835f
C17203 VDD108.t155 VSS 0.0766f
C17204 VDD108.t121 VSS 0.0823f
C17205 VDD108.n74 VSS 0.0393f
C17206 VDD108.t122 VSS 0.00632f
C17207 VDD108.t218 VSS 0.00633f
C17208 VDD108.t135 VSS 0.0766f
C17209 VDD108.n75 VSS 0.00634f
C17210 VDD108.t353 VSS 0.00261f
C17211 VDD108.n76 VSS 0.00261f
C17212 VDD108.n77 VSS 0.00569f
C17213 VDD108.n78 VSS 0.00634f
C17214 VDD108.n79 VSS 0.037f
C17215 VDD108.t14 VSS 0.0763f
C17216 VDD108.n80 VSS 0.00592f
C17217 VDD108.n81 VSS 6.26e-19
C17218 VDD108.t36 VSS 0.00544f
C17219 VDD108.t455 VSS 0.00412f
C17220 VDD108.n82 VSS 0.0106f
C17221 VDD108.n83 VSS 0.0706f
C17222 VDD108.n84 VSS 0.0697f
C17223 VDD108.t466 VSS 0.00411f
C17224 VDD108.t13 VSS 0.00534f
C17225 VDD108.n85 VSS 0.00516f
C17226 VDD108.n86 VSS 0.00557f
C17227 VDD108.n87 VSS 8.95e-19
C17228 VDD108.n88 VSS 0.00473f
C17229 VDD108.n89 VSS 0.0148f
C17230 VDD108.t443 VSS 0.00261f
C17231 VDD108.n90 VSS 0.00261f
C17232 VDD108.n91 VSS 0.00569f
C17233 VDD108.n92 VSS 0.0361f
C17234 VDD108.n93 VSS 0.0362f
C17235 VDD108.n94 VSS 0.0393f
C17236 VDD108.t442 VSS 0.0432f
C17237 VDD108.t214 VSS 0.0933f
C17238 VDD108.t298 VSS 0.0766f
C17239 VDD108.t132 VSS 0.0933f
C17240 VDD108.t352 VSS 0.0432f
C17241 VDD108.n95 VSS 0.0393f
C17242 VDD108.n96 VSS 0.0196f
C17243 VDD108.n97 VSS 0.0361f
C17244 VDD108.n98 VSS 0.0369f
C17245 VDD108.t243 VSS 0.00633f
C17246 VDD108.n99 VSS 0.00634f
C17247 VDD108.n100 VSS 0.0291f
C17248 VDD108.n101 VSS 0.0314f
C17249 VDD108.n102 VSS 0.0219f
C17250 VDD108.n103 VSS 0.0393f
C17251 VDD108.t242 VSS 0.0835f
C17252 VDD108.t184 VSS 0.0766f
C17253 VDD108.t217 VSS 0.0823f
C17254 VDD108.n104 VSS 0.0393f
C17255 VDD108.n105 VSS 0.0219f
C17256 VDD108.n106 VSS 0.0546f
C17257 VDD108.n107 VSS 0.00631f
C17258 VDD108.t439 VSS 0.0559f
C17259 VDD108.n108 VSS 0.0588f
C17260 VDD108.t438 VSS 0.00261f
C17261 VDD108.n109 VSS 0.00261f
C17262 VDD108.n110 VSS 0.00569f
C17263 VDD108.n111 VSS 0.0205f
C17264 VDD108.n112 VSS 0.00634f
C17265 VDD108.t449 VSS 0.0763f
C17266 VDD108.n113 VSS 0.0393f
C17267 VDD108.t223 VSS 0.00633f
C17268 VDD108.n114 VSS 0.00631f
C17269 VDD108.t222 VSS 0.0498f
C17270 VDD108.t158 VSS 0.057f
C17271 VDD108.n115 VSS 0.0987f
C17272 VDD108.n116 VSS 0.0152f
C17273 VDD108.t246 VSS 0.0539f
C17274 VDD108.n117 VSS 0.0382f
C17275 VDD108.n118 VSS 0.00631f
C17276 VDD108.t409 VSS 0.0567f
C17277 VDD108.t143 VSS 0.0562f
C17278 VDD108.n119 VSS 0.0651f
C17279 VDD108.n120 VSS 0.0339f
C17280 VDD108.n121 VSS 0.0338f
C17281 VDD108.n122 VSS 0.0343f
C17282 VDD108.n123 VSS 0.0223f
C17283 VDD108.n124 VSS 0.0311f
C17284 VDD108.n125 VSS 0.0222f
C17285 VDD108.n126 VSS 0.0436f
C17286 VDD108.t219 VSS 0.0435f
C17287 VDD108.n127 VSS 0.00634f
C17288 VDD108.n128 VSS 0.0276f
C17289 VDD108.n129 VSS 0.0219f
C17290 VDD108.n130 VSS 0.00634f
C17291 VDD108.t316 VSS 0.00633f
C17292 VDD108.n131 VSS 0.0314f
C17293 VDD108.n132 VSS 0.0291f
C17294 VDD108.n133 VSS 0.0219f
C17295 VDD108.n134 VSS 0.00634f
C17296 VDD108.t332 VSS 0.00633f
C17297 VDD108.n135 VSS 0.0314f
C17298 VDD108.n136 VSS 0.0291f
C17299 VDD108.t403 VSS 0.00633f
C17300 VDD108.t408 VSS 0.00633f
C17301 VDD108.n137 VSS 0.0688f
C17302 VDD108.t37 VSS 0.0613f
C17303 VDD108.t444 VSS 0.0348f
C17304 VDD108.t410 VSS 0.0613f
C17305 VDD108.t171 VSS 0.0613f
C17306 VDD108.t356 VSS 0.0348f
C17307 VDD108.t320 VSS 0.0218f
C17308 VDD108.n138 VSS 0.00679f
C17309 VDD108.n139 VSS 0.132f
C17310 VDD108.n140 VSS 0.00634f
C17311 VDD108.t445 VSS 0.00261f
C17312 VDD108.n141 VSS 0.00261f
C17313 VDD108.n142 VSS 0.00569f
C17314 VDD108.n143 VSS 0.0361f
C17315 VDD108.n144 VSS 0.037f
C17316 VDD108.t357 VSS 0.00261f
C17317 VDD108.n145 VSS 0.00261f
C17318 VDD108.n146 VSS 0.00569f
C17319 VDD108.n147 VSS 0.00634f
C17320 VDD108.t334 VSS 0.00633f
C17321 VDD108.n148 VSS 0.00634f
C17322 VDD108.n149 VSS 0.0291f
C17323 VDD108.n150 VSS 0.0314f
C17324 VDD108.n151 VSS 0.0219f
C17325 VDD108.n152 VSS 0.0369f
C17326 VDD108.n153 VSS 0.0361f
C17327 VDD108.n154 VSS 0.0196f
C17328 VDD108.n155 VSS 0.0712f
C17329 VDD108.n156 VSS 0.085f
C17330 VDD108.t317 VSS 0.0568f
C17331 VDD108.t333 VSS 0.0613f
C17332 VDD108.t231 VSS 0.0613f
C17333 VDD108.t407 VSS 0.0614f
C17334 VDD108.n157 VSS 0.079f
C17335 VDD108.n158 VSS 0.0219f
C17336 VDD108.n159 VSS 0.0223f
C17337 VDD108.n160 VSS 0.00592f
C17338 VDD108.n161 VSS 6.26e-19
C17339 VDD108.t40 VSS 0.00544f
C17340 VDD108.t464 VSS 0.00412f
C17341 VDD108.n162 VSS 0.0106f
C17342 VDD108.n163 VSS 0.0706f
C17343 VDD108.n164 VSS 0.0697f
C17344 VDD108.t467 VSS 0.00411f
C17345 VDD108.t26 VSS 0.00534f
C17346 VDD108.n165 VSS 0.00516f
C17347 VDD108.n166 VSS 0.00557f
C17348 VDD108.n167 VSS 8.95e-19
C17349 VDD108.n168 VSS 0.00473f
C17350 VDD108.n169 VSS 0.00964f
C17351 VDD108.t27 VSS 0.0763f
C17352 VDD108.n170 VSS 0.0393f
C17353 VDD108.t387 VSS 0.00261f
C17354 VDD108.n171 VSS 0.00261f
C17355 VDD108.n172 VSS 0.00569f
C17356 VDD108.n173 VSS 0.00634f
C17357 VDD108.t386 VSS 0.0432f
C17358 VDD108.t106 VSS 0.0933f
C17359 VDD108.t163 VSS 0.0766f
C17360 VDD108.n174 VSS 0.0393f
C17361 VDD108.t355 VSS 0.00261f
C17362 VDD108.n175 VSS 0.00261f
C17363 VDD108.n176 VSS 0.00569f
C17364 VDD108.n177 VSS 0.00634f
C17365 VDD108.t354 VSS 0.0432f
C17366 VDD108.t234 VSS 0.0933f
C17367 VDD108.t168 VSS 0.0766f
C17368 VDD108.n178 VSS 0.0393f
C17369 VDD108.t73 VSS 0.00633f
C17370 VDD108.n179 VSS 0.00634f
C17371 VDD108.t72 VSS 0.0835f
C17372 VDD108.t140 VSS 0.0766f
C17373 VDD108.t109 VSS 0.0823f
C17374 VDD108.n180 VSS 0.0393f
C17375 VDD108.t110 VSS 0.00633f
C17376 VDD108.n181 VSS 0.00631f
C17377 VDD108.n182 VSS 0.0199f
C17378 VDD108.t149 VSS 0.00633f
C17379 VDD108.t237 VSS 0.0766f
C17380 VDD108.n183 VSS 0.00634f
C17381 VDD108.n184 VSS 0.037f
C17382 VDD108.t5 VSS 0.0571f
C17383 VDD108.t167 VSS 0.00633f
C17384 VDD108.n185 VSS 0.00633f
C17385 VDD108.n186 VSS 0.0452f
C17386 VDD108.n187 VSS 0.0563f
C17387 VDD108.t67 VSS 0.0567f
C17388 VDD108.t382 VSS 0.00261f
C17389 VDD108.n188 VSS 0.00261f
C17390 VDD108.n189 VSS 0.00569f
C17391 VDD108.n190 VSS 0.0446f
C17392 VDD108.t1 VSS 0.0152f
C17393 VDD108.n191 VSS 0.00634f
C17394 VDD108.t176 VSS 0.0435f
C17395 VDD108.t306 VSS 0.00631f
C17396 VDD108.t305 VSS 0.0563f
C17397 VDD108.n192 VSS 0.0651f
C17398 VDD108.n193 VSS 0.0206f
C17399 VDD108.n194 VSS 0.00634f
C17400 VDD108.n195 VSS 0.00661f
C17401 VDD108.t378 VSS 0.0559f
C17402 VDD108.n196 VSS 0.0588f
C17403 VDD108.n197 VSS 0.0268f
C17404 VDD108.n198 VSS 0.0258f
C17405 VDD108.n199 VSS 0.0234f
C17406 VDD108.n200 VSS 0.0393f
C17407 VDD108.t381 VSS 0.0432f
C17408 VDD108.t150 VSS 0.0933f
C17409 VDD108.t116 VSS 0.0766f
C17410 VDD108.t166 VSS 0.0835f
C17411 VDD108.n201 VSS 0.0393f
C17412 VDD108.t6 VSS 0.00797f
C17413 VDD108.n202 VSS 0.015f
C17414 VDD108.n203 VSS 0.0154f
C17415 VDD108.n204 VSS 0.0549f
C17416 VDD108.n205 VSS 0.047f
C17417 VDD108.n206 VSS 0.0257f
C17418 VDD108.n207 VSS 0.0382f
C17419 VDD108.t0 VSS 0.0539f
C17420 VDD108.n208 VSS 0.0987f
C17421 VDD108.t292 VSS 0.0499f
C17422 VDD108.t96 VSS 0.0762f
C17423 VDD108.n209 VSS 0.0393f
C17424 VDD108.n210 VSS 0.0275f
C17425 VDD108.t97 VSS 0.00634f
C17426 VDD108.t75 VSS 0.00633f
C17427 VDD108.t228 VSS 0.00261f
C17428 VDD108.n211 VSS 0.00261f
C17429 VDD108.n212 VSS 0.00569f
C17430 VDD108.n213 VSS 0.0244f
C17431 VDD108.t274 VSS 0.0837f
C17432 VDD108.n214 VSS 0.00633f
C17433 VDD108.t190 VSS 0.00634f
C17434 VDD108.n215 VSS 0.00633f
C17435 VDD108.n216 VSS 0.0314f
C17436 VDD108.t224 VSS 0.0825f
C17437 VDD108.n217 VSS 0.00633f
C17438 VDD108.n218 VSS 0.00633f
C17439 VDD108.t64 VSS 0.0825f
C17440 VDD108.n219 VSS 0.0393f
C17441 VDD108.t147 VSS 0.00634f
C17442 VDD108.n220 VSS 0.00633f
C17443 VDD108.t146 VSS 0.0764f
C17444 VDD108.t396 VSS 0.0837f
C17445 VDD108.n221 VSS 0.0393f
C17446 VDD108.t273 VSS 0.00634f
C17447 VDD108.t188 VSS 0.00261f
C17448 VDD108.n222 VSS 0.00261f
C17449 VDD108.n223 VSS 0.00569f
C17450 VDD108.t272 VSS 0.0764f
C17451 VDD108.t187 VSS 0.0933f
C17452 VDD108.t338 VSS 0.0433f
C17453 VDD108.n224 VSS 0.0393f
C17454 VDD108.t302 VSS 0.00634f
C17455 VDD108.t63 VSS 0.00261f
C17456 VDD108.n225 VSS 0.00261f
C17457 VDD108.n226 VSS 0.00569f
C17458 VDD108.t301 VSS 0.0764f
C17459 VDD108.t62 VSS 0.0933f
C17460 VDD108.t93 VSS 0.0433f
C17461 VDD108.t21 VSS 0.0762f
C17462 VDD108.n227 VSS 0.0393f
C17463 VDD108.t22 VSS 0.00679f
C17464 VDD108.n228 VSS 0.0488f
C17465 VDD108.n229 VSS 0.0361f
C17466 VDD108.n230 VSS 0.037f
C17467 VDD108.n231 VSS 0.0197f
C17468 VDD108.n232 VSS 0.0361f
C17469 VDD108.n233 VSS 0.0369f
C17470 VDD108.n234 VSS 0.0219f
C17471 VDD108.n235 VSS 0.0314f
C17472 VDD108.n236 VSS 0.0292f
C17473 VDD108.n237 VSS 0.0219f
C17474 VDD108.n238 VSS 0.0597f
C17475 VDD108.n239 VSS 0.0679f
C17476 VDD108.t192 VSS 0.00634f
C17477 VDD108.n240 VSS 0.0292f
C17478 VDD108.n241 VSS 0.0219f
C17479 VDD108.n242 VSS 0.0393f
C17480 VDD108.t191 VSS 0.0764f
C17481 VDD108.t393 VSS 0.0837f
C17482 VDD108.t189 VSS 0.0764f
C17483 VDD108.n243 VSS 0.0393f
C17484 VDD108.n244 VSS 0.0219f
C17485 VDD108.n245 VSS 0.0292f
C17486 VDD108.n246 VSS 0.0314f
C17487 VDD108.t359 VSS 0.00634f
C17488 VDD108.n247 VSS 0.0276f
C17489 VDD108.n248 VSS 0.0219f
C17490 VDD108.n249 VSS 0.0393f
C17491 VDD108.t358 VSS 0.0764f
C17492 VDD108.t227 VSS 0.0933f
C17493 VDD108.t90 VSS 0.0433f
C17494 VDD108.n250 VSS 0.0393f
C17495 VDD108.t291 VSS 0.00634f
C17496 VDD108.t89 VSS 0.00631f
C17497 VDD108.n251 VSS 0.00633f
C17498 VDD108.t295 VSS 0.0666f
C17499 VDD108.n252 VSS 0.0339f
C17500 VDD108.t154 VSS 0.00634f
C17501 VDD108.n253 VSS 0.00633f
C17502 VDD108.t153 VSS 0.0608f
C17503 VDD108.t47 VSS 0.0666f
C17504 VDD108.n254 VSS 0.0339f
C17505 VDD108.t84 VSS 0.00634f
C17506 VDD108.t82 VSS 0.00261f
C17507 VDD108.n255 VSS 0.00261f
C17508 VDD108.n256 VSS 0.00569f
C17509 VDD108.n257 VSS 0.0339f
C17510 VDD108.t162 VSS 0.00634f
C17511 VDD108.t289 VSS 0.00261f
C17512 VDD108.n258 VSS 0.00261f
C17513 VDD108.n259 VSS 0.00569f
C17514 VDD108.t161 VSS 0.0608f
C17515 VDD108.t288 VSS 0.0742f
C17516 VDD108.t103 VSS 0.0345f
C17517 VDD108.t83 VSS 0.0554f
C17518 VDD108.t349 VSS 0.0345f
C17519 VDD108.t81 VSS 0.0264f
C17520 VDD108.n260 VSS 0.219f
C17521 VDD108.t34 VSS 0.0697f
C17522 VDD108.n261 VSS 0.0339f
C17523 VDD108.n262 VSS 0.00164f
C17524 VDD108.t457 VSS 0.00412f
C17525 VDD108.t33 VSS 0.00528f
C17526 VDD108.n263 VSS 0.00512f
C17527 VDD108.t462 VSS 0.00412f
C17528 VDD108.t20 VSS 0.00544f
C17529 VDD108.n264 VSS 0.0106f
C17530 VDD108.n265 VSS 0.0596f
C17531 VDD108.n266 VSS 0.0778f
C17532 VDD108.n267 VSS 5.26e-20
C17533 VDD108.n268 VSS 0.00139f
C17534 VDD108.n269 VSS 0.00566f
C17535 VDD108.n270 VSS 7.54e-19
C17536 VDD108.n271 VSS 6.27e-19
C17537 VDD108.n272 VSS 0.00471f
C17538 VDD108.t35 VSS 0.00592f
C17539 VDD108.n273 VSS 0.0148f
C17540 VDD108.n274 VSS 0.0362f
C17541 VDD108.n275 VSS 0.0361f
C17542 VDD108.n276 VSS 0.037f
C17543 VDD108.n277 VSS 0.0197f
C17544 VDD108.n278 VSS 0.0361f
C17545 VDD108.n279 VSS 0.0369f
C17546 VDD108.n280 VSS 0.0219f
C17547 VDD108.n281 VSS 0.0314f
C17548 VDD108.n282 VSS 0.0292f
C17549 VDD108.n283 VSS 0.0219f
C17550 VDD108.n284 VSS 0.0547f
C17551 VDD108.n285 VSS 0.00633f
C17552 VDD108.t360 VSS 0.0825f
C17553 VDD108.n286 VSS 0.0393f
C17554 VDD108.n287 VSS 0.00633f
C17555 VDD108.n288 VSS 0.00634f
C17556 VDD108.t53 VSS 0.0764f
C17557 VDD108.t50 VSS 0.0837f
C17558 VDD108.n289 VSS 0.0393f
C17559 VDD108.t383 VSS 0.0763f
C17560 VDD108.n290 VSS 0.0393f
C17561 VDD108.t80 VSS 0.00634f
C17562 VDD108.t112 VSS 0.00633f
C17563 VDD108.n291 VSS 0.00633f
C17564 VDD108.t111 VSS 0.0498f
C17565 VDD108.t373 VSS 0.057f
C17566 VDD108.n292 VSS 0.0987f
C17567 VDD108.n293 VSS 0.00795f
C17568 VDD108.t79 VSS 0.0764f
C17569 VDD108.t85 VSS 0.0837f
C17570 VDD108.n294 VSS 0.0393f
C17571 VDD108.t366 VSS 0.00634f
C17572 VDD108.n295 VSS 0.0152f
C17573 VDD108.t57 VSS 0.0539f
C17574 VDD108.n296 VSS 0.0382f
C17575 VDD108.t364 VSS 0.00261f
C17576 VDD108.n297 VSS 0.00261f
C17577 VDD108.n298 VSS 0.00569f
C17578 VDD108.t365 VSS 0.0764f
C17579 VDD108.t363 VSS 0.0933f
C17580 VDD108.t98 VSS 0.0433f
C17581 VDD108.n299 VSS 0.0393f
C17582 VDD108.n300 VSS 0.00631f
C17583 VDD108.t372 VSS 0.0567f
C17584 VDD108.t2 VSS 0.0562f
C17585 VDD108.n301 VSS 0.0651f
C17586 VDD108.n302 VSS 0.0206f
C17587 VDD108.t230 VSS 0.00666f
C17588 VDD108.t229 VSS 0.0433f
C17589 VDD108.t101 VSS 0.056f
C17590 VDD108.n303 VSS 0.0588f
C17591 VDD108.t102 VSS 0.0065f
C17592 VDD108.n304 VSS 0.0695f
C17593 VDD108.n305 VSS 0.0214f
C17594 VDD108.n306 VSS 0.0234f
C17595 VDD108.n307 VSS 0.0446f
C17596 VDD108.n308 VSS 0.0259f
C17597 VDD108.n309 VSS 0.0468f
C17598 VDD108.n310 VSS 0.055f
C17599 VDD108.n311 VSS 0.0154f
C17600 VDD108.n312 VSS 0.0152f
C17601 VDD108.n313 VSS 0.0562f
C17602 VDD108.n314 VSS 0.0452f
C17603 VDD108.n315 VSS 0.037f
C17604 VDD108.n316 VSS 0.0277f
C17605 VDD108.n317 VSS 0.0267f
C17606 VDD108.n318 VSS 0.037f
C17607 VDD108.n319 VSS 0.0285f
C17608 VDD108.t392 VSS 0.00261f
C17609 VDD108.n320 VSS 0.00261f
C17610 VDD108.n321 VSS 0.00569f
C17611 VDD108.n322 VSS 0.0205f
C17612 VDD108.n323 VSS 0.00634f
C17613 VDD108.n324 VSS 0.0279f
C17614 VDD108.t388 VSS 0.0559f
C17615 VDD108.n325 VSS 0.0588f
C17616 VDD108.t113 VSS 0.0435f
C17617 VDD108.t280 VSS 0.0835f
C17618 VDD108.n326 VSS 0.00634f
C17619 VDD108.n327 VSS 0.0276f
C17620 VDD108.t281 VSS 0.00633f
C17621 VDD108.n328 VSS 0.00634f
C17622 VDD108.t263 VSS 0.0766f
C17623 VDD108.n329 VSS 0.0393f
C17624 VDD108.t71 VSS 0.00633f
C17625 VDD108.n330 VSS 0.00634f
C17626 VDD108.t70 VSS 0.0835f
C17627 VDD108.t326 VSS 0.0766f
C17628 VDD108.t182 VSS 0.0823f
C17629 VDD108.n331 VSS 0.0393f
C17630 VDD108.t183 VSS 0.00633f
C17631 VDD108.t368 VSS 0.00633f
C17632 VDD108.n332 VSS 0.0688f
C17633 VDD108.t41 VSS 0.0613f
C17634 VDD108.t376 VSS 0.0348f
C17635 VDD108.t369 VSS 0.0613f
C17636 VDD108.t44 VSS 0.0613f
C17637 VDD108.t347 VSS 0.0348f
C17638 VDD108.t266 VSS 0.0218f
C17639 VDD108.n333 VSS 0.00679f
C17640 VDD108.n334 VSS 0.132f
C17641 VDD108.n335 VSS 0.00634f
C17642 VDD108.t377 VSS 0.00261f
C17643 VDD108.n336 VSS 0.00261f
C17644 VDD108.n337 VSS 0.00569f
C17645 VDD108.n338 VSS 0.0361f
C17646 VDD108.n339 VSS 0.037f
C17647 VDD108.t348 VSS 0.00261f
C17648 VDD108.n340 VSS 0.00261f
C17649 VDD108.n341 VSS 0.00569f
C17650 VDD108.n342 VSS 0.00634f
C17651 VDD108.t69 VSS 0.00633f
C17652 VDD108.n343 VSS 0.00634f
C17653 VDD108.n344 VSS 0.0291f
C17654 VDD108.n345 VSS 0.0314f
C17655 VDD108.n346 VSS 0.0219f
C17656 VDD108.n347 VSS 0.0369f
C17657 VDD108.n348 VSS 0.0361f
C17658 VDD108.n349 VSS 0.0196f
C17659 VDD108.n350 VSS 0.0712f
C17660 VDD108.n351 VSS 0.085f
C17661 VDD108.t277 VSS 0.0568f
C17662 VDD108.t68 VSS 0.0613f
C17663 VDD108.t7 VSS 0.0613f
C17664 VDD108.t367 VSS 0.0614f
C17665 VDD108.n352 VSS 0.079f
C17666 VDD108.n353 VSS 0.0219f
C17667 VDD108.n354 VSS 0.0596f
C17668 VDD108.n355 VSS 0.0678f
C17669 VDD108.n356 VSS 0.0219f
C17670 VDD108.n357 VSS 0.0291f
C17671 VDD108.n358 VSS 0.0314f
C17672 VDD108.n359 VSS 0.0219f
C17673 VDD108.n360 VSS 0.0291f
C17674 VDD108.n361 VSS 0.0314f
C17675 VDD108.n362 VSS 0.0219f
C17676 VDD108.n363 VSS 0.0393f
C17677 VDD108.t260 VSS 0.0766f
C17678 VDD108.t179 VSS 0.0933f
C17679 VDD108.t391 VSS 0.0432f
C17680 VDD108.n364 VSS 0.0393f
C17681 VDD108.n365 VSS 0.0146f
C17682 VDD108.n366 VSS 0.0494f
C17683 VDD108.n367 VSS 0.0402f
C17684 VDD108.t54 VSS 0.00652f
C17685 VDD108.n368 VSS 0.0499f
C17686 VDD108.n369 VSS 0.0328f
C17687 VDD108.n370 VSS 0.0548f
C17688 VDD108.n371 VSS 0.074f
C17689 VDD108.n372 VSS 0.0436f
C17690 VDD108.t88 VSS 0.056f
C17691 VDD108.t290 VSS 0.0433f
C17692 VDD108.n373 VSS 0.0588f
C17693 VDD108.n374 VSS 0.0607f
C17694 VDD108.n375 VSS 0.0279f
C17695 VDD108.n376 VSS 0.0465f
C17696 VDD108.n377 VSS 0.00608f
C17697 VDD108.n378 VSS 0.0144f
C17698 VDD108.n379 VSS 0.0627f
C17699 VDD108.n380 VSS 0.0284f
C17700 VDD108.n381 VSS 0.037f
C17701 VDD108.n382 VSS 0.0268f
C17702 VDD108.n383 VSS 0.0393f
C17703 VDD108.t74 VSS 0.0835f
C17704 VDD108.t76 VSS 0.0766f
C17705 VDD108.t148 VSS 0.0823f
C17706 VDD108.n384 VSS 0.0393f
C17707 VDD108.n385 VSS 0.0219f
C17708 VDD108.n386 VSS 0.0321f
C17709 VDD108.n387 VSS 0.0448f
C17710 VDD108.n388 VSS 0.0561f
C17711 VDD108.n389 VSS 0.0219f
C17712 VDD108.n390 VSS 0.0291f
C17713 VDD108.n391 VSS 0.0314f
C17714 VDD108.n392 VSS 0.0219f
C17715 VDD108.n393 VSS 0.0369f
C17716 VDD108.n394 VSS 0.0361f
C17717 VDD108.n395 VSS 0.0196f
C17718 VDD108.n396 VSS 0.037f
C17719 VDD108.n397 VSS 0.0361f
C17720 VDD108.n398 VSS 0.0196f
C17721 VDD108.n399 VSS 0.0706f
C17722 VDD108.n400 VSS 0.0883f
C17723 VDD108.n401 VSS 0.0668f
C17724 VDD108.n402 VSS 0.0219f
C17725 VDD108.t402 VSS 0.0823f
C17726 VDD108.n403 VSS 0.0393f
C17727 VDD108.t335 VSS 0.0766f
C17728 VDD108.t331 VSS 0.0835f
C17729 VDD108.n404 VSS 0.0393f
C17730 VDD108.t323 VSS 0.0766f
C17731 VDD108.t315 VSS 0.0835f
C17732 VDD108.n405 VSS 0.0393f
C17733 VDD108.t269 VSS 0.0766f
C17734 VDD108.t404 VSS 0.0933f
C17735 VDD108.t437 VSS 0.0432f
C17736 VDD108.n406 VSS 0.0393f
C17737 VDD108.n407 VSS 0.0146f
C17738 VDD108.n408 VSS 0.0484f
C17739 VDD108.n409 VSS 0.00655f
C17740 VDD108.n410 VSS 0.0364f
C17741 VDD108.n411 VSS 0.028f
C17742 VDD108.n412 VSS 0.0507f
C17743 VDD108.n413 VSS 0.0329f
C17744 VDD108.n414 VSS 0.0231f
C17745 VDD108.n415 VSS 0.0312f
C17746 VDD108.n416 VSS 0.0338f
C17747 VDD108.n417 VSS 0.0231f
C17748 VDD108.n418 VSS 0.0312f
C17749 VDD108.n419 VSS 0.0338f
C17750 VDD108.n420 VSS 0.0231f
C17751 VDD108.n421 VSS 0.0296f
C17752 VDD108.n422 VSS 0.028f
C17753 VDD108.n423 VSS 0.0204f
C17754 VDD108.n424 VSS 0.0361f
C17755 VDD108.n425 VSS 0.231f
C17756 VDD108.n426 VSS 0.566f
C17757 VDD108.n427 VSS 0.112f
C17758 VDD108.t193 VSS 0.0825f
C17759 VDD108.t303 VSS 0.0764f
C17760 VDD108.n428 VSS 0.0393f
C17761 VDD108.n429 VSS 0.0584f
C17762 VDD108.n430 VSS 0.103f
C17763 VDD108.n431 VSS 0.115f
C17764 VDD108.t201 VSS 0.00634f
C17765 VDD108.n432 VSS 0.103f
C17766 VDD108.n433 VSS 0.0584f
C17767 VDD108.n434 VSS 0.0393f
C17768 VDD108.t200 VSS 0.0764f
C17769 VDD108.t206 VSS 0.0837f
C17770 VDD108.t196 VSS 0.0933f
C17771 VDD108.t198 VSS 0.0764f
C17772 VDD108.n435 VSS 0.0393f
C17773 VDD108.n436 VSS 0.0584f
C17774 VDD108.n437 VSS 0.0956f
C17775 VDD108.n438 VSS 0.0993f
C17776 VDD108.t12 VSS 0.00634f
C17777 VDD108.n439 VSS 0.124f
C17778 VDD108.n440 VSS 0.0472f
C17779 VDD108.n441 VSS 0.0393f
C17780 VDD108.t11 VSS 0.0433f
C17781 VDD108.n442 VSS 0.0588f
C17782 VDD108.n443 VSS 0.0927f
C17783 VDD108.n444 VSS 0.112f
C17784 VDD108.t241 VSS 0.00634f
C17785 VDD108.n445 VSS 0.104f
C17786 VDD108.n446 VSS 0.0586f
C17787 VDD108.n447 VSS 0.0393f
C17788 VDD108.t240 VSS 0.0764f
C17789 VDD108.t434 VSS 0.0837f
C17790 VDD108.t258 VSS 0.0764f
C17791 VDD108.n448 VSS 0.0393f
C17792 VDD108.n449 VSS 0.0586f
C17793 VDD108.n450 VSS 0.104f
C17794 VDD108.n451 VSS 0.115f
C17795 VDD108.t175 VSS 0.00634f
C17796 VDD108.t427 VSS 0.00261f
C17797 VDD108.n452 VSS 0.00261f
C17798 VDD108.n453 VSS 0.00569f
C17799 VDD108.n454 VSS 0.0997f
C17800 VDD108.n455 VSS 0.0959f
C17801 VDD108.n456 VSS 0.0586f
C17802 VDD108.n457 VSS 0.0393f
C17803 VDD108.t174 VSS 0.0764f
C17804 VDD108.t426 VSS 0.0933f
C17805 VDD108.t307 VSS 0.0433f
C17806 VDD108.t18 VSS 0.0433f
C17807 VDD108.n458 VSS 0.0393f
C17808 VDD108.n459 VSS 0.0473f
C17809 VDD108.n460 VSS 0.124f
C17810 VDD108.n461 VSS 0.0927f
C17811 VDD108.t313 VSS 0.0559f
C17812 VDD108.n462 VSS 0.0588f
C17813 VDD108.n463 VSS 0.00637f
C17814 VDD108.n464 VSS 0.00131f
C17815 VDD108.n465 VSS 0.0169f
C17816 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n0 VSS 0.0877f
C17817 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t8 VSS 0.0189f
C17818 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t3 VSS 0.0237f
C17819 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n1 VSS 0.0561f
C17820 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t5 VSS 0.0333f
C17821 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t4 VSS 0.0212f
C17822 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n2 VSS 0.0588f
C17823 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t6 VSS 0.0306f
C17824 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t7 VSS 0.0235f
C17825 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n3 VSS 0.0604f
C17826 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n4 VSS 1.13f
C17827 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n5 VSS 0.378f
C17828 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.t0 VSS 0.0148f
C17829 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n6 VSS 0.0148f
C17830 CLK_div_90_mag_0.CLK_div_10_mag_0.JK_FF_mag_2.K.n7 VSS 0.0349f
C17831 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n0 VSS 0.192f
C17832 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n1 VSS 0.0484f
C17833 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n2 VSS 0.156f
C17834 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n3 VSS 0.00958f
C17835 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n4 VSS 0.186f
C17836 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n5 VSS 0.00958f
C17837 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n6 VSS 0.186f
C17838 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n7 VSS 0.00958f
C17839 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n8 VSS 0.186f
C17840 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n9 VSS 0.00958f
C17841 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n10 VSS 0.0653f
C17842 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n11 VSS 0.0653f
C17843 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n12 VSS 0.0653f
C17844 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n13 VSS 0.0653f
C17845 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n14 VSS 0.0478f
C17846 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n15 VSS 0.0478f
C17847 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n16 VSS 0.0478f
C17848 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n17 VSS 0.0092f
C17849 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t0 VSS 0.00793f
C17850 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t1 VSS 0.0264f
C17851 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n18 VSS 0.0913f
C17852 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t2 VSS 0.0155f
C17853 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t16 VSS 0.0235f
C17854 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n19 VSS 0.0416f
C17855 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t10 VSS 0.0155f
C17856 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t24 VSS 0.0235f
C17857 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n20 VSS 0.0416f
C17858 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t9 VSS 0.0194f
C17859 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t26 VSS 0.00496f
C17860 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n21 VSS 0.0321f
C17861 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t6 VSS 0.0155f
C17862 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t20 VSS 0.0235f
C17863 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n22 VSS 0.0416f
C17864 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t3 VSS 0.0155f
C17865 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t17 VSS 0.0235f
C17866 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n23 VSS 0.0416f
C17867 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t18 VSS 0.0194f
C17868 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t11 VSS 0.00496f
C17869 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n24 VSS 0.0322f
C17870 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t4 VSS 0.0155f
C17871 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t19 VSS 0.0235f
C17872 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n25 VSS 0.0416f
C17873 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t12 VSS 0.0155f
C17874 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t27 VSS 0.0235f
C17875 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n26 VSS 0.0416f
C17876 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t22 VSS 0.0194f
C17877 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t13 VSS 0.00496f
C17878 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n27 VSS 0.0322f
C17879 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t8 VSS 0.0155f
C17880 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t25 VSS 0.0235f
C17881 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n28 VSS 0.0418f
C17882 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t15 VSS 0.0155f
C17883 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t7 VSS 0.0235f
C17884 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n29 VSS 0.0416f
C17885 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t23 VSS 0.0155f
C17886 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t14 VSS 0.0235f
C17887 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n30 VSS 0.0416f
C17888 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t21 VSS 0.00496f
C17889 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.t5 VSS 0.0194f
C17890 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n31 VSS 0.0322f
C17891 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n32 VSS 0.368f
C17892 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n33 VSS 1.93f
C17893 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n34 VSS 1.85f
C17894 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n35 VSS 0.321f
C17895 CLK_div_99_mag_0.CLK_div_3_mag_0.Vdiv3.n36 VSS 0.0147f
C17896 VDD110.t442 VSS 0.00724f
C17897 VDD110.n0 VSS 0.0332f
C17898 VDD110.t441 VSS 0.0684f
C17899 VDD110.n1 VSS 0.0776f
C17900 VDD110.t168 VSS 0.0812f
C17901 VDD110.t324 VSS 0.0816f
C17902 VDD110.n2 VSS 0.0512f
C17903 VDD110.t325 VSS 0.0191f
C17904 VDD110.n3 VSS 0.11f
C17905 VDD110.t343 VSS 0.00724f
C17906 VDD110.n4 VSS 0.0334f
C17907 VDD110.t342 VSS 0.0684f
C17908 VDD110.n5 VSS 0.0776f
C17909 VDD110.t454 VSS 0.0812f
C17910 VDD110.t176 VSS 0.0816f
C17911 VDD110.n6 VSS 0.0512f
C17912 VDD110.t177 VSS 0.019f
C17913 VDD110.n7 VSS 0.111f
C17914 VDD110.t428 VSS 0.00694f
C17915 VDD110.t32 VSS 0.0151f
C17916 VDD110.n8 VSS 0.171f
C17917 VDD110.t292 VSS 0.00727f
C17918 VDD110.t476 VSS 0.00299f
C17919 VDD110.n9 VSS 0.00299f
C17920 VDD110.n10 VSS 0.00653f
C17921 VDD110.t44 VSS 0.00727f
C17922 VDD110.n11 VSS 0.00727f
C17923 VDD110.n12 VSS 0.131f
C17924 VDD110.t116 VSS 0.0856f
C17925 VDD110.t43 VSS 0.0703f
C17926 VDD110.t293 VSS 0.0352f
C17927 VDD110.t117 VSS 0.00914f
C17928 VDD110.t170 VSS 0.0158f
C17929 VDD110.t250 VSS 0.014f
C17930 VDD110.n13 VSS 0.0977f
C17931 VDD110.t249 VSS 0.0479f
C17932 VDD110.t171 VSS 0.093f
C17933 VDD110.t172 VSS 0.0151f
C17934 VDD110.n14 VSS 0.0538f
C17935 VDD110.t248 VSS 0.00728f
C17936 VDD110.t247 VSS 0.0857f
C17937 VDD110.n15 VSS 0.0564f
C17938 VDD110.t89 VSS 0.177f
C17939 VDD110.t118 VSS 0.0589f
C17940 VDD110.t63 VSS 0.0428f
C17941 VDD110.n16 VSS 0.04f
C17942 VDD110.n17 VSS 0.0683f
C17943 VDD110.t62 VSS 0.188f
C17944 VDD110.n18 VSS 0.106f
C17945 VDD110.n19 VSS 0.124f
C17946 VDD110.n20 VSS 0.0732f
C17947 VDD110.n21 VSS 0.102f
C17948 VDD110.t169 VSS 0.0509f
C17949 VDD110.n22 VSS 0.0677f
C17950 VDD110.n23 VSS 0.159f
C17951 VDD110.n24 VSS 0.0705f
C17952 VDD110.n25 VSS 0.0856f
C17953 VDD110.n26 VSS 0.162f
C17954 VDD110.n27 VSS 0.169f
C17955 VDD110.t475 VSS 0.0703f
C17956 VDD110.t291 VSS 0.0703f
C17957 VDD110.t329 VSS 0.053f
C17958 VDD110.n28 VSS 0.0436f
C17959 VDD110.n29 VSS 0.185f
C17960 VDD110.t31 VSS 0.0721f
C17961 VDD110.t427 VSS 0.0866f
C17962 VDD110.n30 VSS 0.0753f
C17963 VDD110.n31 VSS 0.099f
C17964 VDD110.n32 VSS 0.11f
C17965 VDD110.t440 VSS 0.00299f
C17966 VDD110.n33 VSS 0.00299f
C17967 VDD110.n34 VSS 0.00653f
C17968 VDD110.n35 VSS 0.028f
C17969 VDD110.t269 VSS 0.096f
C17970 VDD110.n36 VSS 0.00727f
C17971 VDD110.t277 VSS 0.00727f
C17972 VDD110.n37 VSS 0.00727f
C17973 VDD110.n38 VSS 0.0397f
C17974 VDD110.t436 VSS 0.0947f
C17975 VDD110.n39 VSS 0.00727f
C17976 VDD110.n40 VSS 0.00727f
C17977 VDD110.t431 VSS 0.0947f
C17978 VDD110.n41 VSS 0.0451f
C17979 VDD110.t30 VSS 0.00727f
C17980 VDD110.n42 VSS 0.00727f
C17981 VDD110.t29 VSS 0.0877f
C17982 VDD110.t296 VSS 0.096f
C17983 VDD110.n43 VSS 0.0451f
C17984 VDD110.t273 VSS 0.00727f
C17985 VDD110.t275 VSS 0.00299f
C17986 VDD110.n44 VSS 0.00299f
C17987 VDD110.n45 VSS 0.00653f
C17988 VDD110.t272 VSS 0.0877f
C17989 VDD110.t274 VSS 0.107f
C17990 VDD110.t407 VSS 0.0497f
C17991 VDD110.n46 VSS 0.0451f
C17992 VDD110.t120 VSS 0.00727f
C17993 VDD110.t430 VSS 0.00299f
C17994 VDD110.n47 VSS 0.00299f
C17995 VDD110.n48 VSS 0.00653f
C17996 VDD110.t119 VSS 0.0877f
C17997 VDD110.t429 VSS 0.107f
C17998 VDD110.t469 VSS 0.0497f
C17999 VDD110.t445 VSS 0.0874f
C18000 VDD110.n49 VSS 0.0451f
C18001 VDD110.t446 VSS 0.00779f
C18002 VDD110.n50 VSS 0.056f
C18003 VDD110.n51 VSS 0.0414f
C18004 VDD110.n52 VSS 0.0425f
C18005 VDD110.n53 VSS 0.0226f
C18006 VDD110.n54 VSS 0.0414f
C18007 VDD110.n55 VSS 0.0424f
C18008 VDD110.n56 VSS 0.0251f
C18009 VDD110.n57 VSS 0.036f
C18010 VDD110.n58 VSS 0.0335f
C18011 VDD110.n59 VSS 0.0251f
C18012 VDD110.n60 VSS 0.0631f
C18013 VDD110.t488 VSS 0.00724f
C18014 VDD110.t244 VSS 0.00727f
C18015 VDD110.n61 VSS 0.0421f
C18016 VDD110.t487 VSS 0.0642f
C18017 VDD110.t463 VSS 0.0497f
C18018 VDD110.t456 VSS 0.00299f
C18019 VDD110.n62 VSS 0.00299f
C18020 VDD110.n63 VSS 0.00653f
C18021 VDD110.t414 VSS 0.00727f
C18022 VDD110.n64 VSS 0.00727f
C18023 VDD110.n65 VSS 0.0394f
C18024 VDD110.t306 VSS 0.096f
C18025 VDD110.n66 VSS 0.00727f
C18026 VDD110.t61 VSS 0.00727f
C18027 VDD110.n67 VSS 0.00727f
C18028 VDD110.n68 VSS 0.00727f
C18029 VDD110.t50 VSS 0.0947f
C18030 VDD110.n69 VSS 0.0451f
C18031 VDD110.t313 VSS 0.00727f
C18032 VDD110.n70 VSS 0.00727f
C18033 VDD110.t312 VSS 0.0877f
C18034 VDD110.t309 VSS 0.096f
C18035 VDD110.n71 VSS 0.0451f
C18036 VDD110.t290 VSS 0.00727f
C18037 VDD110.t124 VSS 0.00299f
C18038 VDD110.n72 VSS 0.00299f
C18039 VDD110.n73 VSS 0.00653f
C18040 VDD110.t289 VSS 0.0877f
C18041 VDD110.t123 VSS 0.107f
C18042 VDD110.t389 VSS 0.0497f
C18043 VDD110.n74 VSS 0.0451f
C18044 VDD110.t232 VSS 0.00727f
C18045 VDD110.t49 VSS 0.00299f
C18046 VDD110.n75 VSS 0.00299f
C18047 VDD110.n76 VSS 0.00653f
C18048 VDD110.t231 VSS 0.0877f
C18049 VDD110.t48 VSS 0.107f
C18050 VDD110.t491 VSS 0.0497f
C18051 VDD110.t245 VSS 0.0874f
C18052 VDD110.n77 VSS 0.0451f
C18053 VDD110.t246 VSS 0.00779f
C18054 VDD110.n78 VSS 0.056f
C18055 VDD110.n79 VSS 0.0414f
C18056 VDD110.n80 VSS 0.0425f
C18057 VDD110.n81 VSS 0.0226f
C18058 VDD110.n82 VSS 0.0414f
C18059 VDD110.n83 VSS 0.0424f
C18060 VDD110.n84 VSS 0.0251f
C18061 VDD110.n85 VSS 0.036f
C18062 VDD110.n86 VSS 0.0335f
C18063 VDD110.n87 VSS 0.0251f
C18064 VDD110.n88 VSS 0.0855f
C18065 VDD110.t478 VSS 0.00724f
C18066 VDD110.t279 VSS 0.00727f
C18067 VDD110.n89 VSS 0.0428f
C18068 VDD110.t477 VSS 0.0642f
C18069 VDD110.t479 VSS 0.0497f
C18070 VDD110.t336 VSS 0.00299f
C18071 VDD110.n90 VSS 0.00299f
C18072 VDD110.n91 VSS 0.00653f
C18073 VDD110.t379 VSS 0.00727f
C18074 VDD110.n92 VSS 0.00727f
C18075 VDD110.n93 VSS 0.04f
C18076 VDD110.t236 VSS 0.096f
C18077 VDD110.n94 VSS 0.00727f
C18078 VDD110.t167 VSS 0.00727f
C18079 VDD110.n95 VSS 0.00727f
C18080 VDD110.n96 VSS 0.00727f
C18081 VDD110.t326 VSS 0.0947f
C18082 VDD110.n97 VSS 0.0451f
C18083 VDD110.t122 VSS 0.00727f
C18084 VDD110.n98 VSS 0.00727f
C18085 VDD110.t121 VSS 0.0877f
C18086 VDD110.t233 VSS 0.096f
C18087 VDD110.n99 VSS 0.0451f
C18088 VDD110.t453 VSS 0.00727f
C18089 VDD110.t315 VSS 0.00299f
C18090 VDD110.n100 VSS 0.00299f
C18091 VDD110.n101 VSS 0.00653f
C18092 VDD110.t452 VSS 0.0877f
C18093 VDD110.t314 VSS 0.107f
C18094 VDD110.t392 VSS 0.0497f
C18095 VDD110.n102 VSS 0.0451f
C18096 VDD110.t283 VSS 0.00727f
C18097 VDD110.t319 VSS 0.00299f
C18098 VDD110.n103 VSS 0.00299f
C18099 VDD110.n104 VSS 0.00653f
C18100 VDD110.t282 VSS 0.0877f
C18101 VDD110.t318 VSS 0.107f
C18102 VDD110.t466 VSS 0.0497f
C18103 VDD110.t280 VSS 0.0874f
C18104 VDD110.n105 VSS 0.0451f
C18105 VDD110.t281 VSS 0.00779f
C18106 VDD110.n106 VSS 0.056f
C18107 VDD110.n107 VSS 0.0414f
C18108 VDD110.n108 VSS 0.0425f
C18109 VDD110.n109 VSS 0.0226f
C18110 VDD110.n110 VSS 0.0414f
C18111 VDD110.n111 VSS 0.0424f
C18112 VDD110.n112 VSS 0.0251f
C18113 VDD110.n113 VSS 0.036f
C18114 VDD110.n114 VSS 0.0335f
C18115 VDD110.n115 VSS 0.0251f
C18116 VDD110.n116 VSS 0.0857f
C18117 VDD110.n117 VSS 0.0988f
C18118 VDD110.t332 VSS 0.0947f
C18119 VDD110.t166 VSS 0.0877f
C18120 VDD110.n118 VSS 0.0451f
C18121 VDD110.n119 VSS 0.0269f
C18122 VDD110.n120 VSS 0.037f
C18123 VDD110.n121 VSS 0.04f
C18124 VDD110.t317 VSS 0.00727f
C18125 VDD110.n122 VSS 0.037f
C18126 VDD110.n123 VSS 0.0269f
C18127 VDD110.n124 VSS 0.0451f
C18128 VDD110.t316 VSS 0.0877f
C18129 VDD110.t449 VSS 0.096f
C18130 VDD110.t335 VSS 0.107f
C18131 VDD110.t378 VSS 0.0877f
C18132 VDD110.n125 VSS 0.0451f
C18133 VDD110.n126 VSS 0.0269f
C18134 VDD110.n127 VSS 0.0349f
C18135 VDD110.n128 VSS 0.0332f
C18136 VDD110.n129 VSS 0.0239f
C18137 VDD110.n130 VSS 0.0451f
C18138 VDD110.t278 VSS 0.0497f
C18139 VDD110.n131 VSS 0.0675f
C18140 VDD110.n132 VSS 0.0406f
C18141 VDD110.n133 VSS 0.0453f
C18142 VDD110.n134 VSS 0.0405f
C18143 VDD110.t457 VSS 0.0947f
C18144 VDD110.t60 VSS 0.0877f
C18145 VDD110.n135 VSS 0.0451f
C18146 VDD110.n136 VSS 0.0266f
C18147 VDD110.n137 VSS 0.0365f
C18148 VDD110.n138 VSS 0.0394f
C18149 VDD110.t126 VSS 0.00727f
C18150 VDD110.n139 VSS 0.0365f
C18151 VDD110.n140 VSS 0.0266f
C18152 VDD110.n141 VSS 0.0451f
C18153 VDD110.t125 VSS 0.0877f
C18154 VDD110.t286 VSS 0.096f
C18155 VDD110.t455 VSS 0.107f
C18156 VDD110.t413 VSS 0.0877f
C18157 VDD110.n142 VSS 0.0451f
C18158 VDD110.n143 VSS 0.0266f
C18159 VDD110.n144 VSS 0.0344f
C18160 VDD110.n145 VSS 0.0327f
C18161 VDD110.n146 VSS 0.0237f
C18162 VDD110.n147 VSS 0.0451f
C18163 VDD110.t243 VSS 0.0497f
C18164 VDD110.n148 VSS 0.0675f
C18165 VDD110.n149 VSS 0.0389f
C18166 VDD110.n150 VSS 0.0639f
C18167 VDD110.n151 VSS 0.0388f
C18168 VDD110.t416 VSS 0.00727f
C18169 VDD110.n152 VSS 0.0367f
C18170 VDD110.n153 VSS 0.0267f
C18171 VDD110.n154 VSS 0.0451f
C18172 VDD110.t415 VSS 0.0877f
C18173 VDD110.t299 VSS 0.096f
C18174 VDD110.t276 VSS 0.0877f
C18175 VDD110.n155 VSS 0.0451f
C18176 VDD110.n156 VSS 0.0267f
C18177 VDD110.n157 VSS 0.0367f
C18178 VDD110.n158 VSS 0.0397f
C18179 VDD110.t285 VSS 0.00727f
C18180 VDD110.n159 VSS 0.0347f
C18181 VDD110.n160 VSS 0.0267f
C18182 VDD110.n161 VSS 0.0451f
C18183 VDD110.t284 VSS 0.0877f
C18184 VDD110.t439 VSS 0.107f
C18185 VDD110.t484 VSS 0.0497f
C18186 VDD110.n162 VSS 0.0451f
C18187 VDD110.t448 VSS 0.00727f
C18188 VDD110.t447 VSS 0.0497f
C18189 VDD110.t482 VSS 0.0642f
C18190 VDD110.n163 VSS 0.0675f
C18191 VDD110.t483 VSS 0.00724f
C18192 VDD110.n164 VSS 0.00727f
C18193 VDD110.t90 VSS 0.0947f
C18194 VDD110.n165 VSS 0.0451f
C18195 VDD110.t444 VSS 0.00727f
C18196 VDD110.n166 VSS 0.00727f
C18197 VDD110.t443 VSS 0.0877f
C18198 VDD110.t253 VSS 0.096f
C18199 VDD110.n167 VSS 0.0451f
C18200 VDD110.t139 VSS 0.00727f
C18201 VDD110.t65 VSS 0.00299f
C18202 VDD110.n168 VSS 0.00299f
C18203 VDD110.n169 VSS 0.00653f
C18204 VDD110.t138 VSS 0.0877f
C18205 VDD110.t64 VSS 0.107f
C18206 VDD110.t401 VSS 0.0497f
C18207 VDD110.n170 VSS 0.0451f
C18208 VDD110.t99 VSS 0.00727f
C18209 VDD110.t88 VSS 0.00299f
C18210 VDD110.n171 VSS 0.00299f
C18211 VDD110.n172 VSS 0.00653f
C18212 VDD110.t98 VSS 0.0877f
C18213 VDD110.t87 VSS 0.107f
C18214 VDD110.t460 VSS 0.0497f
C18215 VDD110.t241 VSS 0.0874f
C18216 VDD110.n173 VSS 0.0451f
C18217 VDD110.t242 VSS 0.00779f
C18218 VDD110.n174 VSS 0.056f
C18219 VDD110.n175 VSS 0.0414f
C18220 VDD110.n176 VSS 0.0425f
C18221 VDD110.n177 VSS 0.0226f
C18222 VDD110.n178 VSS 0.0414f
C18223 VDD110.n179 VSS 0.0424f
C18224 VDD110.n180 VSS 0.0251f
C18225 VDD110.n181 VSS 0.036f
C18226 VDD110.n182 VSS 0.0335f
C18227 VDD110.n183 VSS 0.0251f
C18228 VDD110.n184 VSS 0.0631f
C18229 VDD110.n185 VSS 0.00727f
C18230 VDD110.t173 VSS 0.0947f
C18231 VDD110.n186 VSS 0.0451f
C18232 VDD110.t69 VSS 0.00727f
C18233 VDD110.n187 VSS 0.00727f
C18234 VDD110.t68 VSS 0.0877f
C18235 VDD110.t256 VSS 0.096f
C18236 VDD110.n188 VSS 0.0451f
C18237 VDD110.t67 VSS 0.00727f
C18238 VDD110.n189 VSS 0.00727f
C18239 VDD110.t66 VSS 0.0877f
C18240 VDD110.t135 VSS 0.096f
C18241 VDD110.n190 VSS 0.0451f
C18242 VDD110.t181 VSS 0.00727f
C18243 VDD110.t179 VSS 0.00299f
C18244 VDD110.n191 VSS 0.00299f
C18245 VDD110.n192 VSS 0.00653f
C18246 VDD110.t180 VSS 0.0877f
C18247 VDD110.t178 VSS 0.107f
C18248 VDD110.t472 VSS 0.0497f
C18249 VDD110.n193 VSS 0.0451f
C18250 VDD110.t240 VSS 0.00727f
C18251 VDD110.t239 VSS 0.0497f
C18252 VDD110.t489 VSS 0.0642f
C18253 VDD110.n194 VSS 0.0636f
C18254 VDD110.n195 VSS 0.0601f
C18255 VDD110.t490 VSS 0.00724f
C18256 VDD110.n196 VSS 0.0368f
C18257 VDD110.t57 VSS 0.00724f
C18258 VDD110.n197 VSS 0.00727f
C18259 VDD110.t56 VSS 0.0695f
C18260 VDD110.n198 VSS 0.066f
C18261 VDD110.t53 VSS 0.0569f
C18262 VDD110.t320 VSS 0.0874f
C18263 VDD110.n199 VSS 0.0451f
C18264 VDD110.n200 VSS 0.00629f
C18265 VDD110.n201 VSS 0.0777f
C18266 VDD110.t28 VSS 0.0173f
C18267 VDD110.t365 VSS 0.00724f
C18268 VDD110.t435 VSS 0.00299f
C18269 VDD110.n202 VSS 0.00299f
C18270 VDD110.n203 VSS 0.00653f
C18271 VDD110.n204 VSS 0.00727f
C18272 VDD110.n205 VSS 0.0545f
C18273 VDD110.t196 VSS 0.00724f
C18274 VDD110.t45 VSS 0.175f
C18275 VDD110.t47 VSS 0.00727f
C18276 VDD110.t46 VSS 0.00727f
C18277 VDD110.n206 VSS 0.067f
C18278 VDD110.n207 VSS 0.0306f
C18279 VDD110.n208 VSS 0.0902f
C18280 VDD110.t84 VSS 0.0994f
C18281 VDD110.t434 VSS 0.137f
C18282 VDD110.t27 VSS 0.0234f
C18283 VDD110.t195 VSS 0.0967f
C18284 VDD110.t165 VSS 0.00724f
C18285 VDD110.n210 VSS 0.018f
C18286 VDD110.n211 VSS 0.00105f
C18287 VDD110.t77 VSS 0.00724f
C18288 VDD110.n212 VSS 0.15f
C18289 VDD110.n213 VSS 0.201f
C18290 VDD110.t20 VSS 0.00727f
C18291 VDD110.n214 VSS 0.0673f
C18292 VDD110.t76 VSS 0.0643f
C18293 VDD110.t70 VSS 0.0497f
C18294 VDD110.t201 VSS 0.00299f
C18295 VDD110.n215 VSS 0.00299f
C18296 VDD110.n216 VSS 0.00653f
C18297 VDD110.t8 VSS 0.00727f
C18298 VDD110.n217 VSS 0.0308f
C18299 VDD110.n218 VSS 0.223f
C18300 VDD110.t426 VSS 0.00727f
C18301 VDD110.n219 VSS 0.0313f
C18302 VDD110.n220 VSS 0.00727f
C18303 VDD110.t78 VSS 0.096f
C18304 VDD110.n221 VSS 0.00727f
C18305 VDD110.t228 VSS 0.00727f
C18306 VDD110.n222 VSS 0.00727f
C18307 VDD110.n223 VSS 0.00727f
C18308 VDD110.t209 VSS 0.0764f
C18309 VDD110.n224 VSS 0.0389f
C18310 VDD110.t6 VSS 0.00727f
C18311 VDD110.n225 VSS 0.00727f
C18312 VDD110.t5 VSS 0.0697f
C18313 VDD110.t81 VSS 0.0764f
C18314 VDD110.n226 VSS 0.0389f
C18315 VDD110.t338 VSS 0.00727f
C18316 VDD110.t424 VSS 0.00299f
C18317 VDD110.n227 VSS 0.00299f
C18318 VDD110.n228 VSS 0.00653f
C18319 VDD110.n229 VSS 0.0389f
C18320 VDD110.t34 VSS 0.00727f
C18321 VDD110.t206 VSS 0.00299f
C18322 VDD110.n230 VSS 0.00299f
C18323 VDD110.n231 VSS 0.00653f
C18324 VDD110.t33 VSS 0.0697f
C18325 VDD110.t205 VSS 0.0851f
C18326 VDD110.t73 VSS 0.0396f
C18327 VDD110.t337 VSS 0.0636f
C18328 VDD110.t398 VSS 0.0396f
C18329 VDD110.t423 VSS 0.0303f
C18330 VDD110.n232 VSS 0.251f
C18331 VDD110.t22 VSS 0.08f
C18332 VDD110.n233 VSS 0.0389f
C18333 VDD110.t23 VSS 0.00779f
C18334 VDD110.n234 VSS 0.056f
C18335 VDD110.n235 VSS 0.0414f
C18336 VDD110.n236 VSS 0.0425f
C18337 VDD110.n237 VSS 0.0226f
C18338 VDD110.n238 VSS 0.0414f
C18339 VDD110.n239 VSS 0.0424f
C18340 VDD110.n240 VSS 0.0251f
C18341 VDD110.n241 VSS 0.036f
C18342 VDD110.n242 VSS 0.0335f
C18343 VDD110.n243 VSS 0.0251f
C18344 VDD110.n244 VSS 0.0628f
C18345 VDD110.n245 VSS 0.254f
C18346 VDD110.n246 VSS 0.0255f
C18347 VDD110.t190 VSS 0.00727f
C18348 VDD110.t223 VSS 0.0643f
C18349 VDD110.t382 VSS 0.096f
C18350 VDD110.n247 VSS 0.00727f
C18351 VDD110.t386 VSS 0.00727f
C18352 VDD110.n248 VSS 0.0986f
C18353 VDD110.t158 VSS 0.0947f
C18354 VDD110.n249 VSS 0.00727f
C18355 VDD110.n250 VSS 0.0402f
C18356 VDD110.t154 VSS 0.00727f
C18357 VDD110.n251 VSS 0.00727f
C18358 VDD110.n252 VSS 0.0642f
C18359 VDD110.t267 VSS 0.0646f
C18360 VDD110.t268 VSS 0.00724f
C18361 VDD110.n253 VSS 0.054f
C18362 VDD110.t147 VSS 0.0573f
C18363 VDD110.n254 VSS 0.00727f
C18364 VDD110.t101 VSS 0.00724f
C18365 VDD110.t219 VSS 0.00727f
C18366 VDD110.n255 VSS 0.0688f
C18367 VDD110.t100 VSS 0.0646f
C18368 VDD110.t357 VSS 0.0573f
C18369 VDD110.n256 VSS 0.00727f
C18370 VDD110.t252 VSS 0.00724f
C18371 VDD110.t230 VSS 0.00724f
C18372 VDD110.n257 VSS 0.086f
C18373 VDD110.t302 VSS 0.093f
C18374 VDD110.t303 VSS 0.0151f
C18375 VDD110.t305 VSS 0.0282f
C18376 VDD110.n258 VSS 0.0446f
C18377 VDD110.t419 VSS 0.185f
C18378 VDD110.t264 VSS 0.0589f
C18379 VDD110.n259 VSS 0.0683f
C18380 VDD110.t304 VSS 0.188f
C18381 VDD110.n260 VSS 0.0881f
C18382 VDD110.n261 VSS 0.0933f
C18383 VDD110.n262 VSS 0.0569f
C18384 VDD110.n263 VSS 0.102f
C18385 VDD110.t229 VSS 0.0602f
C18386 VDD110.t251 VSS 0.103f
C18387 VDD110.n264 VSS 0.0671f
C18388 VDD110.n265 VSS 0.054f
C18389 VDD110.n266 VSS 0.0642f
C18390 VDD110.n267 VSS 0.0384f
C18391 VDD110.n268 VSS 0.0451f
C18392 VDD110.t218 VSS 0.0497f
C18393 VDD110.n269 VSS 0.106f
C18394 VDD110.n270 VSS 0.054f
C18395 VDD110.n271 VSS 0.0642f
C18396 VDD110.t363 VSS 0.00727f
C18397 VDD110.n272 VSS 0.0688f
C18398 VDD110.n273 VSS 0.0384f
C18399 VDD110.n274 VSS 0.0451f
C18400 VDD110.t362 VSS 0.0497f
C18401 VDD110.n275 VSS 0.106f
C18402 VDD110.t354 VSS 0.0573f
C18403 VDD110.t153 VSS 0.0874f
C18404 VDD110.n276 VSS 0.0451f
C18405 VDD110.n277 VSS 0.0384f
C18406 VDD110.n278 VSS 0.067f
C18407 VDD110.n279 VSS 0.206f
C18408 VDD110.t26 VSS 0.00727f
C18409 VDD110.n280 VSS 0.0505f
C18410 VDD110.t140 VSS 0.0643f
C18411 VDD110.t144 VSS 0.0497f
C18412 VDD110.t347 VSS 0.00299f
C18413 VDD110.n281 VSS 0.00299f
C18414 VDD110.n282 VSS 0.00653f
C18415 VDD110.t59 VSS 0.0073f
C18416 VDD110.n283 VSS 0.00727f
C18417 VDD110.n284 VSS 0.036f
C18418 VDD110.t130 VSS 0.096f
C18419 VDD110.n285 VSS 0.00727f
C18420 VDD110.t134 VSS 0.00727f
C18421 VDD110.n286 VSS 0.00727f
C18422 VDD110.t208 VSS 0.00724f
C18423 VDD110.t113 VSS 0.00727f
C18424 VDD110.n287 VSS 0.0343f
C18425 VDD110.t207 VSS 0.0643f
C18426 VDD110.t215 VSS 0.0497f
C18427 VDD110.t192 VSS 0.00299f
C18428 VDD110.n288 VSS 0.00299f
C18429 VDD110.n289 VSS 0.00653f
C18430 VDD110.t115 VSS 0.00727f
C18431 VDD110.n290 VSS 0.00727f
C18432 VDD110.n291 VSS 0.036f
C18433 VDD110.t373 VSS 0.096f
C18434 VDD110.n292 VSS 0.00727f
C18435 VDD110.t377 VSS 0.00727f
C18436 VDD110.n293 VSS 0.00727f
C18437 VDD110.n294 VSS 0.00727f
C18438 VDD110.t420 VSS 0.0947f
C18439 VDD110.n295 VSS 0.0451f
C18440 VDD110.t194 VSS 0.00727f
C18441 VDD110.n296 VSS 0.00727f
C18442 VDD110.t193 VSS 0.0877f
C18443 VDD110.t370 VSS 0.096f
C18444 VDD110.n297 VSS 0.0451f
C18445 VDD110.t4 VSS 0.00727f
C18446 VDD110.t369 VSS 0.00299f
C18447 VDD110.n298 VSS 0.00299f
C18448 VDD110.n299 VSS 0.00653f
C18449 VDD110.t3 VSS 0.0877f
C18450 VDD110.t368 VSS 0.107f
C18451 VDD110.t404 VSS 0.0497f
C18452 VDD110.n300 VSS 0.0451f
C18453 VDD110.t103 VSS 0.00727f
C18454 VDD110.t418 VSS 0.00299f
C18455 VDD110.n301 VSS 0.00299f
C18456 VDD110.n302 VSS 0.00653f
C18457 VDD110.t102 VSS 0.0877f
C18458 VDD110.t417 VSS 0.107f
C18459 VDD110.t220 VSS 0.0497f
C18460 VDD110.t13 VSS 0.0874f
C18461 VDD110.n303 VSS 0.0451f
C18462 VDD110.n304 VSS 0.00216f
C18463 VDD110.t499 VSS 0.00473f
C18464 VDD110.t9 VSS 0.00624f
C18465 VDD110.n305 VSS 0.0122f
C18466 VDD110.n306 VSS 0.00287f
C18467 VDD110.n307 VSS 0.00148f
C18468 VDD110.n308 VSS 7.48e-19
C18469 VDD110.n309 VSS 0.00666f
C18470 VDD110.n310 VSS 0.00182f
C18471 VDD110.t18 VSS 0.0062f
C18472 VDD110.t496 VSS 0.00473f
C18473 VDD110.n311 VSS 0.0122f
C18474 VDD110.n312 VSS 0.0023f
C18475 VDD110.n313 VSS 0.00194f
C18476 VDD110.n314 VSS 7.48e-19
C18477 VDD110.n315 VSS 0.0236f
C18478 VDD110.n316 VSS 7.19e-19
C18479 VDD110.t495 VSS 0.00473f
C18480 VDD110.t21 VSS 0.00589f
C18481 VDD110.n317 VSS 0.00603f
C18482 VDD110.n318 VSS 0.00202f
C18483 VDD110.n319 VSS 0.00649f
C18484 VDD110.n320 VSS 0.0022f
C18485 VDD110.n321 VSS 0.0914f
C18486 VDD110.n322 VSS 0.133f
C18487 VDD110.n323 VSS 0.00182f
C18488 VDD110.t24 VSS 0.0062f
C18489 VDD110.t494 VSS 0.00473f
C18490 VDD110.n324 VSS 0.0122f
C18491 VDD110.n325 VSS 0.00238f
C18492 VDD110.n326 VSS 0.00187f
C18493 VDD110.n327 VSS 7.48e-19
C18494 VDD110.n328 VSS 0.0236f
C18495 VDD110.t497 VSS 0.00483f
C18496 VDD110.t15 VSS 0.00612f
C18497 VDD110.n329 VSS 0.0122f
C18498 VDD110.n330 VSS 0.00445f
C18499 VDD110.n331 VSS 0.0308f
C18500 VDD110.n332 VSS 0.148f
C18501 VDD110.t498 VSS 0.00473f
C18502 VDD110.t12 VSS 0.00624f
C18503 VDD110.n333 VSS 0.0122f
C18504 VDD110.n334 VSS 0.0623f
C18505 VDD110.n335 VSS 7.06e-19
C18506 VDD110.n336 VSS 0.00584f
C18507 VDD110.t14 VSS 0.00679f
C18508 VDD110.n337 VSS 0.0169f
C18509 VDD110.n338 VSS 0.0415f
C18510 VDD110.n339 VSS 0.0414f
C18511 VDD110.n340 VSS 0.0425f
C18512 VDD110.n341 VSS 0.0226f
C18513 VDD110.n342 VSS 0.0414f
C18514 VDD110.n343 VSS 0.0424f
C18515 VDD110.n344 VSS 0.0251f
C18516 VDD110.n345 VSS 0.036f
C18517 VDD110.n346 VSS 0.0335f
C18518 VDD110.n347 VSS 0.0251f
C18519 VDD110.n348 VSS 0.0686f
C18520 VDD110.n349 VSS 0.0779f
C18521 VDD110.t186 VSS 0.0947f
C18522 VDD110.t376 VSS 0.0877f
C18523 VDD110.n350 VSS 0.0451f
C18524 VDD110.n351 VSS 0.0251f
C18525 VDD110.n352 VSS 0.0335f
C18526 VDD110.n353 VSS 0.036f
C18527 VDD110.t367 VSS 0.00727f
C18528 VDD110.n354 VSS 0.0335f
C18529 VDD110.n355 VSS 0.0251f
C18530 VDD110.n356 VSS 0.0451f
C18531 VDD110.t366 VSS 0.0877f
C18532 VDD110.t0 VSS 0.096f
C18533 VDD110.t191 VSS 0.107f
C18534 VDD110.t114 VSS 0.0877f
C18535 VDD110.n357 VSS 0.0451f
C18536 VDD110.n358 VSS 0.0251f
C18537 VDD110.n359 VSS 0.0317f
C18538 VDD110.n360 VSS 0.0297f
C18539 VDD110.n361 VSS 0.0226f
C18540 VDD110.n362 VSS 0.0451f
C18541 VDD110.t112 VSS 0.0497f
C18542 VDD110.n363 VSS 0.0675f
C18543 VDD110.n364 VSS 0.0228f
C18544 VDD110.n365 VSS 0.00727f
C18545 VDD110.t351 VSS 0.0764f
C18546 VDD110.n366 VSS 0.0389f
C18547 VDD110.t345 VSS 0.00727f
C18548 VDD110.n367 VSS 0.00727f
C18549 VDD110.t344 VSS 0.0697f
C18550 VDD110.t127 VSS 0.0764f
C18551 VDD110.n368 VSS 0.0389f
C18552 VDD110.t260 VSS 0.00727f
C18553 VDD110.t111 VSS 0.00299f
C18554 VDD110.n369 VSS 0.00299f
C18555 VDD110.n370 VSS 0.00653f
C18556 VDD110.n371 VSS 0.0389f
C18557 VDD110.t226 VSS 0.00727f
C18558 VDD110.t361 VSS 0.00299f
C18559 VDD110.n372 VSS 0.00299f
C18560 VDD110.n373 VSS 0.00653f
C18561 VDD110.t225 VSS 0.0697f
C18562 VDD110.t360 VSS 0.0851f
C18563 VDD110.t155 VSS 0.0396f
C18564 VDD110.t259 VSS 0.0636f
C18565 VDD110.t410 VSS 0.0396f
C18566 VDD110.t110 VSS 0.0303f
C18567 VDD110.n374 VSS 0.251f
C18568 VDD110.t16 VSS 0.08f
C18569 VDD110.n375 VSS 0.0389f
C18570 VDD110.t17 VSS 0.00779f
C18571 VDD110.n376 VSS 0.056f
C18572 VDD110.n377 VSS 0.0414f
C18573 VDD110.n378 VSS 0.0425f
C18574 VDD110.n379 VSS 0.0226f
C18575 VDD110.n380 VSS 0.0414f
C18576 VDD110.n381 VSS 0.0424f
C18577 VDD110.n382 VSS 0.0251f
C18578 VDD110.n383 VSS 0.036f
C18579 VDD110.n384 VSS 0.0335f
C18580 VDD110.n385 VSS 0.0251f
C18581 VDD110.n386 VSS 0.0644f
C18582 VDD110.n387 VSS 0.0514f
C18583 VDD110.n388 VSS 0.0369f
C18584 VDD110.t348 VSS 0.0947f
C18585 VDD110.t133 VSS 0.0877f
C18586 VDD110.n389 VSS 0.0451f
C18587 VDD110.n390 VSS 0.0251f
C18588 VDD110.n391 VSS 0.0335f
C18589 VDD110.n392 VSS 0.036f
C18590 VDD110.t109 VSS 0.00727f
C18591 VDD110.n393 VSS 0.0335f
C18592 VDD110.n394 VSS 0.0251f
C18593 VDD110.n395 VSS 0.0451f
C18594 VDD110.t108 VSS 0.0877f
C18595 VDD110.t261 VSS 0.096f
C18596 VDD110.t346 VSS 0.107f
C18597 VDD110.t58 VSS 0.0877f
C18598 VDD110.n396 VSS 0.0451f
C18599 VDD110.n397 VSS 0.0251f
C18600 VDD110.n398 VSS 0.0358f
C18601 VDD110.n399 VSS 0.101f
C18602 VDD110.n400 VSS 0.0545f
C18603 VDD110.n401 VSS 0.0318f
C18604 VDD110.n402 VSS 0.0451f
C18605 VDD110.t25 VSS 0.0497f
C18606 VDD110.n403 VSS 0.0675f
C18607 VDD110.t141 VSS 0.00724f
C18608 VDD110.n404 VSS 0.00727f
C18609 VDD110.t150 VSS 0.0764f
C18610 VDD110.n405 VSS 0.0389f
C18611 VDD110.t266 VSS 0.00727f
C18612 VDD110.n406 VSS 0.00727f
C18613 VDD110.t265 VSS 0.0697f
C18614 VDD110.t38 VSS 0.0764f
C18615 VDD110.n407 VSS 0.0389f
C18616 VDD110.t381 VSS 0.00727f
C18617 VDD110.t388 VSS 0.00299f
C18618 VDD110.n408 VSS 0.00299f
C18619 VDD110.n409 VSS 0.00653f
C18620 VDD110.n410 VSS 0.0389f
C18621 VDD110.t183 VSS 0.00727f
C18622 VDD110.t143 VSS 0.00299f
C18623 VDD110.n411 VSS 0.00299f
C18624 VDD110.n412 VSS 0.00653f
C18625 VDD110.t182 VSS 0.0697f
C18626 VDD110.t142 VSS 0.0851f
C18627 VDD110.t212 VSS 0.0396f
C18628 VDD110.t380 VSS 0.0636f
C18629 VDD110.t395 VSS 0.0396f
C18630 VDD110.t387 VSS 0.0303f
C18631 VDD110.n413 VSS 0.251f
C18632 VDD110.t10 VSS 0.08f
C18633 VDD110.n414 VSS 0.0389f
C18634 VDD110.t11 VSS 0.00779f
C18635 VDD110.n415 VSS 0.056f
C18636 VDD110.n416 VSS 0.0414f
C18637 VDD110.n417 VSS 0.0425f
C18638 VDD110.n418 VSS 0.0226f
C18639 VDD110.n419 VSS 0.0414f
C18640 VDD110.n420 VSS 0.0424f
C18641 VDD110.n421 VSS 0.0251f
C18642 VDD110.n422 VSS 0.036f
C18643 VDD110.n423 VSS 0.0335f
C18644 VDD110.n424 VSS 0.0251f
C18645 VDD110.n425 VSS 0.0628f
C18646 VDD110.n426 VSS 0.0844f
C18647 VDD110.n427 VSS 0.0497f
C18648 VDD110.n428 VSS 0.117f
C18649 VDD110.n429 VSS 0.252f
C18650 VDD110.n430 VSS 0.243f
C18651 VDD110.n431 VSS 0.242f
C18652 VDD110.n432 VSS 0.0984f
C18653 VDD110.t105 VSS 0.00727f
C18654 VDD110.n433 VSS 0.00727f
C18655 VDD110.n434 VSS 0.0549f
C18656 VDD110.n435 VSS 0.0585f
C18657 VDD110.n436 VSS 0.0372f
C18658 VDD110.n437 VSS 0.0451f
C18659 VDD110.t104 VSS 0.0877f
C18660 VDD110.t35 VSS 0.096f
C18661 VDD110.t385 VSS 0.0877f
C18662 VDD110.n438 VSS 0.0451f
C18663 VDD110.n439 VSS 0.0243f
C18664 VDD110.n440 VSS 0.0585f
C18665 VDD110.n441 VSS 0.0642f
C18666 VDD110.t107 VSS 0.00727f
C18667 VDD110.t162 VSS 0.00299f
C18668 VDD110.n442 VSS 0.00299f
C18669 VDD110.n443 VSS 0.00653f
C18670 VDD110.n444 VSS 0.0545f
C18671 VDD110.n445 VSS 0.05f
C18672 VDD110.n446 VSS 0.0928f
C18673 VDD110.n447 VSS 0.0374f
C18674 VDD110.n448 VSS 0.0451f
C18675 VDD110.t106 VSS 0.0877f
C18676 VDD110.t161 VSS 0.107f
C18677 VDD110.t202 VSS 0.0497f
C18678 VDD110.n449 VSS 0.0451f
C18679 VDD110.t189 VSS 0.0497f
C18680 VDD110.n450 VSS 0.0675f
C18681 VDD110.t224 VSS 0.00724f
C18682 VDD110.n451 VSS 0.0427f
C18683 VDD110.n452 VSS 0.0359f
C18684 VDD110.n453 VSS 0.093f
C18685 VDD110.n454 VSS 0.244f
C18686 VDD110.n455 VSS 0.228f
C18687 VDD110.n456 VSS 0.0831f
C18688 VDD110.n457 VSS 0.0645f
C18689 VDD110.n458 VSS 0.0624f
C18690 VDD110.t197 VSS 0.0947f
C18691 VDD110.t227 VSS 0.0877f
C18692 VDD110.n459 VSS 0.0451f
C18693 VDD110.n460 VSS 0.0374f
C18694 VDD110.n461 VSS 0.0318f
C18695 VDD110.n462 VSS 0.106f
C18696 VDD110.n463 VSS 0.0614f
C18697 VDD110.n464 VSS 0.0374f
C18698 VDD110.n465 VSS 0.0451f
C18699 VDD110.t425 VSS 0.0877f
C18700 VDD110.t339 VSS 0.096f
C18701 VDD110.t200 VSS 0.107f
C18702 VDD110.t7 VSS 0.0877f
C18703 VDD110.n466 VSS 0.0451f
C18704 VDD110.n467 VSS 0.0374f
C18705 VDD110.n468 VSS 0.0619f
C18706 VDD110.n469 VSS 0.106f
C18707 VDD110.n470 VSS 0.213f
C18708 VDD110.n471 VSS 0.212f
C18709 VDD110.n472 VSS 0.102f
C18710 VDD110.n473 VSS 0.0521f
C18711 VDD110.n474 VSS 0.0983f
C18712 VDD110.n475 VSS 0.0318f
C18713 VDD110.n476 VSS 0.0451f
C18714 VDD110.t19 VSS 0.0497f
C18715 VDD110.n477 VSS 0.0675f
C18716 VDD110.n478 VSS 0.117f
C18717 VDD110.n479 VSS 0.914f
C18718 VDD110.n480 VSS 0.5f
C18719 VDD110.n481 VSS 0.305f
C18720 VDD110.n482 VSS 0.00738f
C18721 VDD110.n484 VSS 0.00369f
C18722 VDD110.n485 VSS 0.0554f
C18723 VDD110.t164 VSS 0.0645f
C18724 VDD110.n486 VSS 0.0756f
C18725 VDD110.t163 VSS 0.0607f
C18726 VDD110.n487 VSS 0.026f
C18727 VDD110.n488 VSS 0.0914f
C18728 VDD110.n489 VSS 0.0541f
C18729 VDD110.n490 VSS 0.0257f
C18730 VDD110.n491 VSS 0.0139f
C18731 VDD110.n492 VSS 0.0756f
C18732 VDD110.t364 VSS 0.0892f
C18733 VDD110.n493 VSS 0.0619f
C18734 VDD110.n494 VSS 0.0327f
C18735 VDD110.n495 VSS 0.0362f
C18736 VDD110.n496 VSS 0.0248f
C18737 VDD110.t321 VSS 0.00739f
C18738 VDD110.n497 VSS 0.0404f
C18739 VDD110.n498 VSS 0.0255f
C18740 VDD110.n499 VSS 0.0357f
C18741 VDD110.n500 VSS 0.0334f
C18742 VDD110.n501 VSS 0.0299f
C18743 VDD110.n502 VSS 0.0373f
C18744 VDD110.n503 VSS 0.0237f
C18745 VDD110.n504 VSS 0.0327f
C18746 VDD110.n505 VSS 0.0344f
C18747 VDD110.n506 VSS 0.0266f
C18748 VDD110.n507 VSS 0.0394f
C18749 VDD110.n508 VSS 0.0365f
C18750 VDD110.n509 VSS 0.0266f
C18751 VDD110.n510 VSS 0.0394f
C18752 VDD110.n511 VSS 0.0365f
C18753 VDD110.n512 VSS 0.0266f
C18754 VDD110.n513 VSS 0.0385f
C18755 VDD110.n514 VSS 0.0647f
C18756 VDD110.n515 VSS 0.0404f
C18757 VDD110.n516 VSS 0.0425f
C18758 VDD110.n517 VSS 0.0238f
C18759 VDD110.n518 VSS 0.111f
C18760 VDD110.n519 VSS 1.12f
C18761 VDD110.n520 VSS 0.553f
C18762 VDD110.n521 VSS 0.522f
C18763 VDD110.t42 VSS 0.00727f
C18764 VDD110.n522 VSS 0.00727f
C18765 VDD110.n523 VSS 0.0357f
C18766 VDD110.t96 VSS 0.0856f
C18767 VDD110.t41 VSS 0.0703f
C18768 VDD110.t93 VSS 0.0352f
C18769 VDD110.t97 VSS 0.00724f
C18770 VDD110.n524 VSS 0.0256f
C18771 VDD110.n525 VSS 0.0705f
C18772 VDD110.n526 VSS 0.0511f
C18773 VDD110.n527 VSS 0.0975f
C18774 VDD110.n528 VSS 0.00396f
C18775 VDD110.n529 VSS 6.48e-19
C18776 VDD110.n530 VSS 0.00727f
C18777 VDD110.n531 VSS 7.79e-19
C18778 VDD110.n532 VSS 0.00112f
C18779 VDD110.n533 VSS 0.00246f
C18780 VDD110.n534 VSS 0.00263f
C18781 VDD110.n535 VSS 7.58e-19
C18782 VDD110.n536 VSS 0.00781f
C18783 VDD110.n537 VSS 0.897f
C18784 VDD110.n538 VSS 0.714f
C18785 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n0 VSS 0.826f
C18786 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n1 VSS 0.0344f
C18787 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n2 VSS 0.254f
C18788 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n3 VSS 0.0151f
C18789 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n4 VSS 0.241f
C18790 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n5 VSS 0.0151f
C18791 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n6 VSS 0.15f
C18792 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n7 VSS 0.103f
C18793 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n8 VSS 0.103f
C18794 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n9 VSS 0.035f
C18795 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t0 VSS 0.0201f
C18796 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t2 VSS 0.0165f
C18797 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n10 VSS 0.0165f
C18798 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n11 VSS 0.0397f
C18799 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n12 VSS 0.124f
C18800 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t5 VSS 0.0368f
C18801 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t4 VSS 0.0243f
C18802 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n13 VSS 0.0654f
C18803 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n14 VSS 0.257f
C18804 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t20 VSS 0.0264f
C18805 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t19 VSS 0.0211f
C18806 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n15 VSS 0.0614f
C18807 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n16 VSS 0.0381f
C18808 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n17 VSS 0.488f
C18809 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t10 VSS 0.0368f
C18810 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t7 VSS 0.0243f
C18811 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n18 VSS 0.0651f
C18812 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t11 VSS 0.0368f
C18813 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t6 VSS 0.0243f
C18814 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n19 VSS 0.0651f
C18815 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t17 VSS 0.0304f
C18816 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t3 VSS 0.00786f
C18817 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n20 VSS 0.0504f
C18818 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t18 VSS 0.0368f
C18819 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t16 VSS 0.0243f
C18820 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n21 VSS 0.0651f
C18821 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t15 VSS 0.0368f
C18822 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t13 VSS 0.0243f
C18823 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n22 VSS 0.0651f
C18824 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n23 VSS 0.11f
C18825 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t8 VSS 0.0342f
C18826 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t12 VSS 0.0189f
C18827 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n24 VSS 0.0652f
C18828 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n25 VSS 0.869f
C18829 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t9 VSS 0.0304f
C18830 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.t14 VSS 0.00786f
C18831 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n26 VSS 0.0504f
C18832 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n27 VSS 0.124f
C18833 CLK_div_100_mag_0.CLK_div_10_mag_1.Q0.n28 VSS 0.0156f
C18834 F0.n0 VSS 0.103f
C18835 F0.t20 VSS 0.013f
C18836 F0.t13 VSS 0.0163f
C18837 F0.n1 VSS 0.0385f
C18838 F0.n2 VSS 0.0202f
C18839 F0.n3 VSS 0.00376f
C18840 F0.t18 VSS 0.00474f
C18841 F0.t3 VSS 0.0188f
C18842 F0.n4 VSS 0.0307f
C18843 F0.n5 VSS 0.0105f
C18844 F0.n6 VSS 0.0748f
C18845 F0.n7 VSS 0.186f
C18846 F0.n8 VSS 0.109f
C18847 F0.n9 VSS 0.00552f
C18848 F0.t8 VSS 0.013f
C18849 F0.t2 VSS 0.0163f
C18850 F0.n10 VSS 0.0385f
C18851 F0.n11 VSS 2.22e-19
C18852 F0.n12 VSS 0.0098f
C18853 F0.n13 VSS 0.00537f
C18854 F0.n14 VSS 0.00395f
C18855 F0.t4 VSS 0.0188f
C18856 F0.t6 VSS 0.00474f
C18857 F0.n15 VSS 0.0307f
C18858 F0.n16 VSS 0.0105f
C18859 F0.t11 VSS 0.013f
C18860 F0.t24 VSS 0.0163f
C18861 F0.n17 VSS 0.0385f
C18862 F0.n18 VSS 0.0202f
C18863 F0.n19 VSS 0.00376f
C18864 F0.t19 VSS 0.0188f
C18865 F0.t22 VSS 0.00474f
C18866 F0.n20 VSS 0.0307f
C18867 F0.n21 VSS 0.0105f
C18868 F0.n22 VSS 0.0749f
C18869 F0.n23 VSS 0.186f
C18870 F0.n24 VSS 0.00553f
C18871 F0.t17 VSS 0.013f
C18872 F0.t9 VSS 0.0163f
C18873 F0.n25 VSS 0.0385f
C18874 F0.n26 VSS 0.0157f
C18875 F0.n27 VSS 2.22e-19
C18876 F0.n28 VSS 0.109f
C18877 F0.n29 VSS 0.0768f
C18878 F0.n30 VSS 0.0762f
C18879 F0.n31 VSS 0.00395f
C18880 F0.n32 VSS 0.108f
C18881 F0.n33 VSS 0.108f
C18882 F0.t14 VSS 0.00474f
C18883 F0.t23 VSS 0.0188f
C18884 F0.n34 VSS 0.0307f
C18885 F0.n35 VSS 0.0105f
C18886 F0.n36 VSS 0.0739f
C18887 F0.n37 VSS 2.51f
C18888 F0.n38 VSS 0.00182f
C18889 F0.t12 VSS 0.0226f
C18890 F0.t10 VSS 0.0149f
C18891 F0.n39 VSS 0.0401f
C18892 F0.n40 VSS 7.39e-19
C18893 F0.n41 VSS 0.00109f
C18894 F0.n42 VSS 0.0024f
C18895 F0.n43 VSS 0.00265f
C18896 F0.n44 VSS 0.0112f
C18897 F0.n45 VSS 0.00859f
C18898 F0.t16 VSS 0.0226f
C18899 F0.t15 VSS 0.0149f
C18900 F0.n46 VSS 0.0399f
C18901 F0.n47 VSS 0.00272f
C18902 F0.n48 VSS 0.00608f
C18903 F0.t0 VSS 0.0143f
C18904 F0.n49 VSS 0.0134f
C18905 F0.n50 VSS 0.0012f
C18906 F0.t1 VSS 0.0225f
C18907 F0.n51 VSS 0.0275f
C18908 F0.n52 VSS 0.00232f
C18909 F0.n53 VSS 0.00538f
C18910 F0.n54 VSS 0.00289f
C18911 F0.t7 VSS 0.0226f
C18912 F0.t5 VSS 0.0149f
C18913 F0.n55 VSS 0.0401f
C18914 F0.n56 VSS 0.00227f
C18915 F0.n57 VSS 0.106f
C18916 F0.n58 VSS 0.204f
C18917 F0.n59 VSS 0.196f
C18918 F0.n60 VSS 0.157f
C18919 F0.t25 VSS 0.00414f
C18920 F0.n61 VSS 0.0105f
C18921 F0.t21 VSS 0.0186f
C18922 F0.n62 VSS 0.021f
C18923 F0.n63 VSS 0.00202f
C18924 F0.n64 VSS 0.00129f
C18925 F0.n65 VSS 0.00486f
C18926 F0.n66 VSS 0.00666f
C18927 F0.n67 VSS 0.0694f
C18928 F0.n68 VSS 0.078f
C18929 F0.n69 VSS 4.79f
C18930 VDD100.t483 VSS 0.00407f
C18931 VDD100.t89 VSS 0.00537f
C18932 VDD100.n0 VSS 0.0105f
C18933 VDD100.n1 VSS 0.00186f
C18934 VDD100.n2 VSS 0.00128f
C18935 VDD100.t492 VSS 0.00407f
C18936 VDD100.t71 VSS 0.00537f
C18937 VDD100.n3 VSS 0.0105f
C18938 VDD100.n4 VSS 0.00244f
C18939 VDD100.n5 VSS 6.43e-19
C18940 VDD100.n6 VSS 0.00573f
C18941 VDD100.n7 VSS 0.00156f
C18942 VDD100.n8 VSS 0.00167f
C18943 VDD100.t85 VSS 0.00534f
C18944 VDD100.t487 VSS 0.00407f
C18945 VDD100.n9 VSS 0.0105f
C18946 VDD100.n10 VSS 0.00197f
C18947 VDD100.n11 VSS 6.43e-19
C18948 VDD100.n12 VSS 0.0203f
C18949 VDD100.n13 VSS 0.00177f
C18950 VDD100.t489 VSS 0.00407f
C18951 VDD100.n14 VSS 0.00559f
C18952 VDD100.t75 VSS 0.00526f
C18953 VDD100.n15 VSS 0.005f
C18954 VDD100.n16 VSS 0.00246f
C18955 VDD100.n17 VSS 0.0786f
C18956 VDD100.n18 VSS 0.115f
C18957 VDD100.n19 VSS 0.00156f
C18958 VDD100.n20 VSS 0.00161f
C18959 VDD100.t64 VSS 0.00534f
C18960 VDD100.t481 VSS 0.00407f
C18961 VDD100.n21 VSS 0.0105f
C18962 VDD100.n22 VSS 0.00205f
C18963 VDD100.n23 VSS 6.43e-19
C18964 VDD100.n24 VSS 0.0203f
C18965 VDD100.t477 VSS 0.00416f
C18966 VDD100.t102 VSS 0.00526f
C18967 VDD100.n25 VSS 0.0105f
C18968 VDD100.n26 VSS 0.00381f
C18969 VDD100.n27 VSS 0.0265f
C18970 VDD100.n28 VSS 0.127f
C18971 VDD100.n29 VSS 0.0527f
C18972 VDD100.n30 VSS 0.00379f
C18973 VDD100.n31 VSS 0.00584f
C18974 VDD100.n32 VSS 0.0163f
C18975 VDD100.t90 VSS 0.0754f
C18976 VDD100.t341 VSS 0.0921f
C18977 VDD100.t403 VSS 0.0426f
C18978 VDD100.n33 VSS 0.0388f
C18979 VDD100.n34 VSS 0.0357f
C18980 VDD100.t404 VSS 0.00257f
C18981 VDD100.n35 VSS 0.00257f
C18982 VDD100.n36 VSS 0.00562f
C18983 VDD100.n37 VSS 0.00626f
C18984 VDD100.t8 VSS 0.0756f
C18985 VDD100.n38 VSS 0.0388f
C18986 VDD100.t376 VSS 0.00257f
C18987 VDD100.n39 VSS 0.00257f
C18988 VDD100.n40 VSS 0.00562f
C18989 VDD100.n41 VSS 0.00626f
C18990 VDD100.t375 VSS 0.0426f
C18991 VDD100.t322 VSS 0.0921f
C18992 VDD100.t3 VSS 0.0756f
C18993 VDD100.n42 VSS 0.0388f
C18994 VDD100.t114 VSS 0.00625f
C18995 VDD100.n43 VSS 0.00626f
C18996 VDD100.t113 VSS 0.0825f
C18997 VDD100.t0 VSS 0.0756f
C18998 VDD100.t344 VSS 0.0813f
C18999 VDD100.n44 VSS 0.0388f
C19000 VDD100.t345 VSS 0.00625f
C19001 VDD100.t128 VSS 0.00625f
C19002 VDD100.t325 VSS 0.0756f
C19003 VDD100.n45 VSS 0.00626f
C19004 VDD100.t7 VSS 0.00625f
C19005 VDD100.t14 VSS 0.0429f
C19006 VDD100.n46 VSS 0.00626f
C19007 VDD100.n47 VSS 0.00623f
C19008 VDD100.t228 VSS 0.00625f
C19009 VDD100.t31 VSS 0.0756f
C19010 VDD100.n48 VSS 0.00626f
C19011 VDD100.t378 VSS 0.00257f
C19012 VDD100.n49 VSS 0.00257f
C19013 VDD100.n50 VSS 0.00562f
C19014 VDD100.n51 VSS 0.00626f
C19015 VDD100.n52 VSS 0.0366f
C19016 VDD100.t103 VSS 0.0754f
C19017 VDD100.n53 VSS 0.00671f
C19018 VDD100.t423 VSS 0.00257f
C19019 VDD100.n54 VSS 0.00257f
C19020 VDD100.n55 VSS 0.00562f
C19021 VDD100.n56 VSS 0.0357f
C19022 VDD100.n57 VSS 0.0482f
C19023 VDD100.n58 VSS 0.0388f
C19024 VDD100.t422 VSS 0.0426f
C19025 VDD100.t229 VSS 0.0921f
C19026 VDD100.t148 VSS 0.0756f
C19027 VDD100.t286 VSS 0.0921f
C19028 VDD100.t377 VSS 0.0426f
C19029 VDD100.n59 VSS 0.0388f
C19030 VDD100.n60 VSS 0.0194f
C19031 VDD100.n61 VSS 0.0357f
C19032 VDD100.n62 VSS 0.0364f
C19033 VDD100.t193 VSS 0.00625f
C19034 VDD100.n63 VSS 0.00626f
C19035 VDD100.n64 VSS 0.0288f
C19036 VDD100.n65 VSS 0.031f
C19037 VDD100.n66 VSS 0.0217f
C19038 VDD100.n67 VSS 0.0388f
C19039 VDD100.t192 VSS 0.0825f
C19040 VDD100.t432 VSS 0.0756f
C19041 VDD100.t227 VSS 0.0813f
C19042 VDD100.n68 VSS 0.0388f
C19043 VDD100.n69 VSS 0.0217f
C19044 VDD100.n70 VSS 0.0553f
C19045 VDD100.t436 VSS 0.00625f
C19046 VDD100.t289 VSS 0.0756f
C19047 VDD100.n71 VSS 0.00626f
C19048 VDD100.t35 VSS 0.00625f
C19049 VDD100.t65 VSS 0.0429f
C19050 VDD100.n72 VSS 0.00626f
C19051 VDD100.n73 VSS 0.0296f
C19052 VDD100.t421 VSS 0.00257f
C19053 VDD100.n74 VSS 0.00257f
C19054 VDD100.n75 VSS 0.00562f
C19055 VDD100.n76 VSS 0.00626f
C19056 VDD100.t427 VSS 0.0754f
C19057 VDD100.n77 VSS 0.0388f
C19058 VDD100.t223 VSS 0.00625f
C19059 VDD100.n78 VSS 0.00623f
C19060 VDD100.t222 VSS 0.0491f
C19061 VDD100.t41 VSS 0.0556f
C19062 VDD100.n79 VSS 0.0909f
C19063 VDD100.n80 VSS 0.00626f
C19064 VDD100.t224 VSS 0.0429f
C19065 VDD100.n81 VSS 0.0388f
C19066 VDD100.t431 VSS 0.00625f
C19067 VDD100.n82 VSS 0.00623f
C19068 VDD100.t430 VSS 0.0491f
C19069 VDD100.t283 VSS 0.0556f
C19070 VDD100.n83 VSS 0.0909f
C19071 VDD100.n84 VSS 0.00626f
C19072 VDD100.t239 VSS 0.0429f
C19073 VDD100.n85 VSS 0.0388f
C19074 VDD100.t233 VSS 0.00625f
C19075 VDD100.n86 VSS 0.00623f
C19076 VDD100.t232 VSS 0.0491f
C19077 VDD100.n87 VSS 0.0577f
C19078 VDD100.t304 VSS 0.0888f
C19079 VDD100.t280 VSS 0.0518f
C19080 VDD100.n88 VSS 0.0882f
C19081 VDD100.n89 VSS 0.00623f
C19082 VDD100.t390 VSS 0.08f
C19083 VDD100.n90 VSS 0.0482f
C19084 VDD100.t411 VSS 0.00257f
C19085 VDD100.n91 VSS 0.00257f
C19086 VDD100.n92 VSS 0.00564f
C19087 VDD100.n93 VSS 0.0198f
C19088 VDD100.n94 VSS 0.191f
C19089 VDD100.t274 VSS 0.0497f
C19090 VDD100.n95 VSS 0.00625f
C19091 VDD100.t308 VSS 0.00626f
C19092 VDD100.n96 VSS 0.00625f
C19093 VDD100.n97 VSS 0.031f
C19094 VDD100.t412 VSS 0.0657f
C19095 VDD100.n98 VSS 0.00625f
C19096 VDD100.t462 VSS 0.00623f
C19097 VDD100.t248 VSS 0.00626f
C19098 VDD100.n99 VSS 0.0295f
C19099 VDD100.t247 VSS 0.034f
C19100 VDD100.t153 VSS 0.0444f
C19101 VDD100.n100 VSS 0.00625f
C19102 VDD100.t154 VSS 0.00626f
C19103 VDD100.n101 VSS 0.00625f
C19104 VDD100.n102 VSS 0.031f
C19105 VDD100.t165 VSS 0.0657f
C19106 VDD100.n103 VSS 0.00625f
C19107 VDD100.t172 VSS 0.00623f
C19108 VDD100.t70 VSS 0.00626f
C19109 VDD100.n104 VSS 0.0295f
C19110 VDD100.t69 VSS 0.034f
C19111 VDD100.t117 VSS 0.0444f
C19112 VDD100.n105 VSS 0.00625f
C19113 VDD100.t118 VSS 0.00626f
C19114 VDD100.n106 VSS 0.00625f
C19115 VDD100.n107 VSS 0.031f
C19116 VDD100.t48 VSS 0.0657f
C19117 VDD100.n108 VSS 0.00625f
C19118 VDD100.t452 VSS 0.00623f
C19119 VDD100.t156 VSS 0.00626f
C19120 VDD100.n109 VSS 0.0295f
C19121 VDD100.t451 VSS 0.0552f
C19122 VDD100.t448 VSS 0.0428f
C19123 VDD100.t250 VSS 0.00257f
C19124 VDD100.n110 VSS 0.00257f
C19125 VDD100.n111 VSS 0.00562f
C19126 VDD100.t158 VSS 0.00626f
C19127 VDD100.n112 VSS 0.00625f
C19128 VDD100.n113 VSS 0.031f
C19129 VDD100.t28 VSS 0.0826f
C19130 VDD100.n114 VSS 0.00625f
C19131 VDD100.t402 VSS 0.00626f
C19132 VDD100.n115 VSS 0.00625f
C19133 VDD100.n116 VSS 0.00625f
C19134 VDD100.t314 VSS 0.0814f
C19135 VDD100.n117 VSS 0.0388f
C19136 VDD100.t145 VSS 0.00626f
C19137 VDD100.n118 VSS 0.00625f
C19138 VDD100.t144 VSS 0.0754f
C19139 VDD100.t25 VSS 0.0826f
C19140 VDD100.n119 VSS 0.0388f
C19141 VDD100.t56 VSS 0.00626f
C19142 VDD100.t54 VSS 0.00257f
C19143 VDD100.n120 VSS 0.00257f
C19144 VDD100.n121 VSS 0.00562f
C19145 VDD100.t55 VSS 0.0754f
C19146 VDD100.t53 VSS 0.0921f
C19147 VDD100.t369 VSS 0.0428f
C19148 VDD100.n122 VSS 0.0388f
C19149 VDD100.t197 VSS 0.00626f
C19150 VDD100.t312 VSS 0.00257f
C19151 VDD100.n123 VSS 0.00257f
C19152 VDD100.n124 VSS 0.00562f
C19153 VDD100.t196 VSS 0.0754f
C19154 VDD100.t311 VSS 0.0921f
C19155 VDD100.t440 VSS 0.0428f
C19156 VDD100.t94 VSS 0.0752f
C19157 VDD100.n125 VSS 0.0388f
C19158 VDD100.t95 VSS 0.00584f
C19159 VDD100.t93 VSS 0.00537f
C19160 VDD100.t480 VSS 0.00407f
C19161 VDD100.n126 VSS 0.0105f
C19162 VDD100.n127 VSS 0.00186f
C19163 VDD100.t96 VSS 0.00537f
C19164 VDD100.t479 VSS 0.00407f
C19165 VDD100.n128 VSS 0.0105f
C19166 VDD100.n129 VSS 0.00247f
C19167 VDD100.n130 VSS 0.00127f
C19168 VDD100.n131 VSS 6.43e-19
C19169 VDD100.n132 VSS 0.00573f
C19170 VDD100.n133 VSS 6.18e-19
C19171 VDD100.t79 VSS 0.00521f
C19172 VDD100.n134 VSS 0.00515f
C19173 VDD100.t486 VSS 0.00406f
C19174 VDD100.n135 VSS 0.00174f
C19175 VDD100.n136 VSS 0.0055f
C19176 VDD100.n137 VSS 0.0019f
C19177 VDD100.n138 VSS 0.00156f
C19178 VDD100.t99 VSS 0.00534f
C19179 VDD100.t478 VSS 0.00407f
C19180 VDD100.n139 VSS 0.0105f
C19181 VDD100.n140 VSS 0.00197f
C19182 VDD100.n141 VSS 0.00167f
C19183 VDD100.n142 VSS 6.43e-19
C19184 VDD100.n143 VSS 0.0203f
C19185 VDD100.n144 VSS 0.0786f
C19186 VDD100.n145 VSS 0.115f
C19187 VDD100.t485 VSS 0.00415f
C19188 VDD100.t82 VSS 0.00527f
C19189 VDD100.n146 VSS 0.0105f
C19190 VDD100.n147 VSS 0.00383f
C19191 VDD100.n148 VSS 0.00156f
C19192 VDD100.t490 VSS 0.00407f
C19193 VDD100.t68 VSS 0.00534f
C19194 VDD100.n149 VSS 0.0105f
C19195 VDD100.n150 VSS 0.00205f
C19196 VDD100.n151 VSS 0.00161f
C19197 VDD100.n152 VSS 6.43e-19
C19198 VDD100.n153 VSS 0.0203f
C19199 VDD100.n154 VSS 0.0265f
C19200 VDD100.n155 VSS 0.127f
C19201 VDD100.n156 VSS 0.0536f
C19202 VDD100.n157 VSS 6.07e-19
C19203 VDD100.n158 VSS 0.00503f
C19204 VDD100.n159 VSS 0.0145f
C19205 VDD100.n160 VSS 0.0357f
C19206 VDD100.n161 VSS 0.0356f
C19207 VDD100.n162 VSS 0.0366f
C19208 VDD100.n163 VSS 0.0194f
C19209 VDD100.n164 VSS 0.0356f
C19210 VDD100.n165 VSS 0.0365f
C19211 VDD100.n166 VSS 0.0216f
C19212 VDD100.n167 VSS 0.031f
C19213 VDD100.n168 VSS 0.0288f
C19214 VDD100.n169 VSS 0.0216f
C19215 VDD100.n170 VSS 0.059f
C19216 VDD100.n171 VSS 0.0671f
C19217 VDD100.t251 VSS 0.0814f
C19218 VDD100.t401 VSS 0.0754f
C19219 VDD100.n172 VSS 0.0388f
C19220 VDD100.n173 VSS 0.0216f
C19221 VDD100.n174 VSS 0.0288f
C19222 VDD100.n175 VSS 0.031f
C19223 VDD100.t52 VSS 0.00626f
C19224 VDD100.n176 VSS 0.0288f
C19225 VDD100.n177 VSS 0.0216f
C19226 VDD100.n178 VSS 0.0388f
C19227 VDD100.t51 VSS 0.0754f
C19228 VDD100.t57 VSS 0.0826f
C19229 VDD100.t249 VSS 0.0921f
C19230 VDD100.t157 VSS 0.0754f
C19231 VDD100.n179 VSS 0.0388f
C19232 VDD100.n180 VSS 0.0216f
C19233 VDD100.n181 VSS 0.0273f
C19234 VDD100.n182 VSS 0.0256f
C19235 VDD100.n183 VSS 0.0194f
C19236 VDD100.n184 VSS 0.0388f
C19237 VDD100.t155 VSS 0.0428f
C19238 VDD100.n185 VSS 0.0581f
C19239 VDD100.n186 VSS 0.0196f
C19240 VDD100.n187 VSS 0.00625f
C19241 VDD100.t205 VSS 0.0814f
C19242 VDD100.n188 VSS 0.0388f
C19243 VDD100.t45 VSS 0.00626f
C19244 VDD100.n189 VSS 0.00625f
C19245 VDD100.t44 VSS 0.0754f
C19246 VDD100.t267 VSS 0.0826f
C19247 VDD100.n190 VSS 0.0388f
C19248 VDD100.t21 VSS 0.00626f
C19249 VDD100.t120 VSS 0.00257f
C19250 VDD100.n191 VSS 0.00257f
C19251 VDD100.n192 VSS 0.00562f
C19252 VDD100.t20 VSS 0.0754f
C19253 VDD100.t119 VSS 0.0921f
C19254 VDD100.t379 VSS 0.0428f
C19255 VDD100.n193 VSS 0.0388f
C19256 VDD100.t294 VSS 0.00626f
C19257 VDD100.t217 VSS 0.00257f
C19258 VDD100.n194 VSS 0.00257f
C19259 VDD100.n195 VSS 0.00562f
C19260 VDD100.t293 VSS 0.0754f
C19261 VDD100.t216 VSS 0.0921f
C19262 VDD100.t181 VSS 0.0428f
C19263 VDD100.t83 VSS 0.0752f
C19264 VDD100.n196 VSS 0.0388f
C19265 VDD100.t84 VSS 0.00671f
C19266 VDD100.n197 VSS 0.0482f
C19267 VDD100.n198 VSS 0.0356f
C19268 VDD100.n199 VSS 0.0366f
C19269 VDD100.n200 VSS 0.0194f
C19270 VDD100.n201 VSS 0.0356f
C19271 VDD100.n202 VSS 0.0365f
C19272 VDD100.n203 VSS 0.0216f
C19273 VDD100.n204 VSS 0.031f
C19274 VDD100.n205 VSS 0.0288f
C19275 VDD100.n206 VSS 0.0216f
C19276 VDD100.n207 VSS 0.0554f
C19277 VDD100.n208 VSS 0.0443f
C19278 VDD100.n209 VSS 0.0317f
C19279 VDD100.t329 VSS 0.00626f
C19280 VDD100.n210 VSS 0.0288f
C19281 VDD100.n211 VSS 0.0216f
C19282 VDD100.n212 VSS 0.0335f
C19283 VDD100.t328 VSS 0.06f
C19284 VDD100.t264 VSS 0.0657f
C19285 VDD100.n213 VSS 0.0335f
C19286 VDD100.n214 VSS 0.0216f
C19287 VDD100.n215 VSS 0.0288f
C19288 VDD100.n216 VSS 0.031f
C19289 VDD100.n217 VSS 0.0216f
C19290 VDD100.t47 VSS 0.00257f
C19291 VDD100.n218 VSS 0.00257f
C19292 VDD100.n219 VSS 0.00562f
C19293 VDD100.t185 VSS 0.00626f
C19294 VDD100.n220 VSS 0.00625f
C19295 VDD100.n221 VSS 0.0307f
C19296 VDD100.t219 VSS 0.00623f
C19297 VDD100.n222 VSS 0.022f
C19298 VDD100.t218 VSS 0.0555f
C19299 VDD100.t173 VSS 0.0493f
C19300 VDD100.n223 VSS 0.00625f
C19301 VDD100.t61 VSS 0.00623f
C19302 VDD100.t457 VSS 0.00626f
C19303 VDD100.n224 VSS 0.0291f
C19304 VDD100.t60 VSS 0.0555f
C19305 VDD100.t208 VSS 0.0493f
C19306 VDD100.n225 VSS 0.00625f
C19307 VDD100.t160 VSS 0.00623f
C19308 VDD100.t162 VSS 0.00635f
C19309 VDD100.n226 VSS 0.034f
C19310 VDD100.t121 VSS 0.08f
C19311 VDD100.t122 VSS 0.00623f
C19312 VDD100.n227 VSS 0.0281f
C19313 VDD100.t86 VSS 0.0586f
C19314 VDD100.t124 VSS 0.0243f
C19315 VDD100.n228 VSS 0.00626f
C19316 VDD100.n229 VSS 0.00653f
C19317 VDD100.t313 VSS 0.206f
C19318 VDD100.t292 VSS 0.0738f
C19319 VDD100.t123 VSS 0.0918f
C19320 VDD100.n230 VSS 0.0793f
C19321 VDD100.n231 VSS 0.0108f
C19322 VDD100.n232 VSS 0.0275f
C19323 VDD100.n233 VSS 0.0294f
C19324 VDD100.n234 VSS 0.0181f
C19325 VDD100.n235 VSS 0.061f
C19326 VDD100.t262 VSS 0.0825f
C19327 VDD100.n236 VSS 0.00626f
C19328 VDD100.t360 VSS 0.00257f
C19329 VDD100.n237 VSS 0.00257f
C19330 VDD100.n238 VSS 0.00564f
C19331 VDD100.n239 VSS 0.0197f
C19332 VDD100.n240 VSS 0.0273f
C19333 VDD100.t263 VSS 0.00625f
C19334 VDD100.n241 VSS 0.00626f
C19335 VDD100.t141 VSS 0.0756f
C19336 VDD100.n242 VSS 0.0388f
C19337 VDD100.t364 VSS 0.00625f
C19338 VDD100.n243 VSS 0.00626f
C19339 VDD100.t363 VSS 0.0825f
C19340 VDD100.t332 VSS 0.0756f
C19341 VDD100.t203 VSS 0.0813f
C19342 VDD100.n244 VSS 0.0388f
C19343 VDD100.t204 VSS 0.00625f
C19344 VDD100.n245 VSS 0.00623f
C19345 VDD100.t242 VSS 0.0553f
C19346 VDD100.n246 VSS 0.0581f
C19347 VDD100.n247 VSS 0.00626f
C19348 VDD100.t132 VSS 0.0429f
C19349 VDD100.n248 VSS 0.0388f
C19350 VDD100.t258 VSS 0.00257f
C19351 VDD100.n249 VSS 0.00257f
C19352 VDD100.n250 VSS 0.00562f
C19353 VDD100.n251 VSS 0.00626f
C19354 VDD100.t257 VSS 0.0426f
C19355 VDD100.t319 VSS 0.0921f
C19356 VDD100.t347 VSS 0.0756f
C19357 VDD100.n252 VSS 0.0388f
C19358 VDD100.t400 VSS 0.00625f
C19359 VDD100.n253 VSS 0.00626f
C19360 VDD100.t399 VSS 0.0825f
C19361 VDD100.t186 VSS 0.0756f
C19362 VDD100.n254 VSS 0.0388f
C19363 VDD100.t351 VSS 0.00625f
C19364 VDD100.n255 VSS 0.00626f
C19365 VDD100.t350 VSS 0.0825f
C19366 VDD100.t354 VSS 0.0756f
C19367 VDD100.t317 VSS 0.0813f
C19368 VDD100.n256 VSS 0.0388f
C19369 VDD100.t318 VSS 0.00625f
C19370 VDD100.n257 VSS 0.00623f
C19371 VDD100.t424 VSS 0.0553f
C19372 VDD100.n258 VSS 0.0581f
C19373 VDD100.n259 VSS 0.0196f
C19374 VDD100.t419 VSS 0.00625f
C19375 VDD100.t396 VSS 0.0756f
C19376 VDD100.n260 VSS 0.00626f
C19377 VDD100.t386 VSS 0.00257f
C19378 VDD100.n261 VSS 0.00257f
C19379 VDD100.n262 VSS 0.00562f
C19380 VDD100.n263 VSS 0.00626f
C19381 VDD100.n264 VSS 0.0366f
C19382 VDD100.t72 VSS 0.0754f
C19383 VDD100.n265 VSS 0.00671f
C19384 VDD100.t238 VSS 0.00257f
C19385 VDD100.n266 VSS 0.00257f
C19386 VDD100.n267 VSS 0.00562f
C19387 VDD100.n268 VSS 0.0357f
C19388 VDD100.n269 VSS 0.0482f
C19389 VDD100.n270 VSS 0.0388f
C19390 VDD100.t237 VSS 0.0426f
C19391 VDD100.t415 VSS 0.0921f
C19392 VDD100.t295 VSS 0.0756f
C19393 VDD100.t189 VSS 0.0921f
C19394 VDD100.t385 VSS 0.0426f
C19395 VDD100.n271 VSS 0.0388f
C19396 VDD100.n272 VSS 0.0194f
C19397 VDD100.n273 VSS 0.0357f
C19398 VDD100.n274 VSS 0.0364f
C19399 VDD100.t353 VSS 0.00625f
C19400 VDD100.n275 VSS 0.00626f
C19401 VDD100.n276 VSS 0.0288f
C19402 VDD100.n277 VSS 0.031f
C19403 VDD100.n278 VSS 0.0217f
C19404 VDD100.n279 VSS 0.0388f
C19405 VDD100.t352 VSS 0.0825f
C19406 VDD100.t277 VSS 0.0756f
C19407 VDD100.t418 VSS 0.0813f
C19408 VDD100.n280 VSS 0.0388f
C19409 VDD100.n281 VSS 0.0217f
C19410 VDD100.n282 VSS 0.0553f
C19411 VDD100.n283 VSS 0.0441f
C19412 VDD100.n284 VSS 0.0317f
C19413 VDD100.n285 VSS 0.0217f
C19414 VDD100.n286 VSS 0.0288f
C19415 VDD100.n287 VSS 0.031f
C19416 VDD100.n288 VSS 0.0217f
C19417 VDD100.n289 VSS 0.0288f
C19418 VDD100.n290 VSS 0.031f
C19419 VDD100.n291 VSS 0.0217f
C19420 VDD100.n292 VSS 0.0273f
C19421 VDD100.n293 VSS 0.0256f
C19422 VDD100.n294 VSS 0.0194f
C19423 VDD100.n295 VSS 0.0296f
C19424 VDD100.n296 VSS 0.0192f
C19425 VDD100.t409 VSS 0.00625f
C19426 VDD100.t259 VSS 0.0756f
C19427 VDD100.n297 VSS 0.00626f
C19428 VDD100.t368 VSS 0.00257f
C19429 VDD100.n298 VSS 0.00257f
C19430 VDD100.n299 VSS 0.00562f
C19431 VDD100.n300 VSS 0.00626f
C19432 VDD100.n301 VSS 0.0366f
C19433 VDD100.t76 VSS 0.0754f
C19434 VDD100.n302 VSS 0.00671f
C19435 VDD100.t358 VSS 0.00257f
C19436 VDD100.n303 VSS 0.00257f
C19437 VDD100.n304 VSS 0.00562f
C19438 VDD100.n305 VSS 0.0357f
C19439 VDD100.n306 VSS 0.0482f
C19440 VDD100.n307 VSS 0.0388f
C19441 VDD100.t357 VSS 0.0426f
C19442 VDD100.t254 VSS 0.0921f
C19443 VDD100.t234 VSS 0.0756f
C19444 VDD100.t138 VSS 0.0921f
C19445 VDD100.t367 VSS 0.0426f
C19446 VDD100.n308 VSS 0.0388f
C19447 VDD100.n309 VSS 0.0194f
C19448 VDD100.n310 VSS 0.0357f
C19449 VDD100.n311 VSS 0.0364f
C19450 VDD100.t366 VSS 0.00625f
C19451 VDD100.n312 VSS 0.00626f
C19452 VDD100.n313 VSS 0.0288f
C19453 VDD100.n314 VSS 0.031f
C19454 VDD100.n315 VSS 0.0217f
C19455 VDD100.n316 VSS 0.0388f
C19456 VDD100.t365 VSS 0.0825f
C19457 VDD100.t393 VSS 0.0756f
C19458 VDD100.t408 VSS 0.0813f
C19459 VDD100.n317 VSS 0.0388f
C19460 VDD100.n318 VSS 0.0217f
C19461 VDD100.n319 VSS 0.0553f
C19462 VDD100.n320 VSS 0.0392f
C19463 VDD100.n321 VSS 0.0317f
C19464 VDD100.n322 VSS 0.0217f
C19465 VDD100.n323 VSS 0.0288f
C19466 VDD100.n324 VSS 0.031f
C19467 VDD100.n325 VSS 0.0217f
C19468 VDD100.n326 VSS 0.0288f
C19469 VDD100.n327 VSS 0.031f
C19470 VDD100.n328 VSS 0.0217f
C19471 VDD100.n329 VSS 0.0388f
C19472 VDD100.t11 VSS 0.0756f
C19473 VDD100.t200 VSS 0.0921f
C19474 VDD100.t359 VSS 0.0397f
C19475 VDD100.n330 VSS 0.0606f
C19476 VDD100.n331 VSS 0.0482f
C19477 VDD100.n332 VSS 0.0296f
C19478 VDD100.n333 VSS 0.0205f
C19479 VDD100.n334 VSS 0.0882f
C19480 VDD100.t161 VSS 0.0521f
C19481 VDD100.t159 VSS 0.0884f
C19482 VDD100.n335 VSS 0.0577f
C19483 VDD100.n336 VSS 0.022f
C19484 VDD100.n337 VSS 0.0307f
C19485 VDD100.n338 VSS 0.0219f
C19486 VDD100.n339 VSS 0.0388f
C19487 VDD100.t456 VSS 0.0428f
C19488 VDD100.n340 VSS 0.0909f
C19489 VDD100.n341 VSS 0.022f
C19490 VDD100.n342 VSS 0.0307f
C19491 VDD100.t215 VSS 0.00626f
C19492 VDD100.n343 VSS 0.0291f
C19493 VDD100.n344 VSS 0.0219f
C19494 VDD100.n345 VSS 0.0388f
C19495 VDD100.t214 VSS 0.0428f
C19496 VDD100.n346 VSS 0.0909f
C19497 VDD100.t211 VSS 0.0493f
C19498 VDD100.t184 VSS 0.0752f
C19499 VDD100.n347 VSS 0.0388f
C19500 VDD100.n348 VSS 0.0219f
C19501 VDD100.n349 VSS 0.0563f
C19502 VDD100.t199 VSS 0.00626f
C19503 VDD100.n350 VSS 0.0205f
C19504 VDD100.n351 VSS 0.0314f
C19505 VDD100.n352 VSS 0.0256f
C19506 VDD100.n353 VSS 0.0194f
C19507 VDD100.n354 VSS 0.0335f
C19508 VDD100.t168 VSS 0.034f
C19509 VDD100.t46 VSS 0.0733f
C19510 VDD100.t198 VSS 0.06f
C19511 VDD100.n355 VSS 0.0335f
C19512 VDD100.t22 VSS 0.0288f
C19513 VDD100.n356 VSS 0.174f
C19514 VDD100.n357 VSS 0.0958f
C19515 VDD100.t171 VSS 0.0689f
C19516 VDD100.n358 VSS 0.0196f
C19517 VDD100.n359 VSS 0.00625f
C19518 VDD100.t176 VSS 0.0814f
C19519 VDD100.n360 VSS 0.0388f
C19520 VDD100.t147 VSS 0.00626f
C19521 VDD100.n361 VSS 0.00625f
C19522 VDD100.t146 VSS 0.0754f
C19523 VDD100.t463 VSS 0.0826f
C19524 VDD100.n362 VSS 0.0388f
C19525 VDD100.t40 VSS 0.00626f
C19526 VDD100.t152 VSS 0.00257f
C19527 VDD100.n363 VSS 0.00257f
C19528 VDD100.n364 VSS 0.00562f
C19529 VDD100.t39 VSS 0.0754f
C19530 VDD100.t151 VSS 0.0921f
C19531 VDD100.t382 VSS 0.0428f
C19532 VDD100.n365 VSS 0.0388f
C19533 VDD100.t107 VSS 0.00626f
C19534 VDD100.t180 VSS 0.00257f
C19535 VDD100.n366 VSS 0.00257f
C19536 VDD100.n367 VSS 0.00562f
C19537 VDD100.t106 VSS 0.0754f
C19538 VDD100.t179 VSS 0.0921f
C19539 VDD100.t445 VSS 0.0428f
C19540 VDD100.t97 VSS 0.0752f
C19541 VDD100.n368 VSS 0.0388f
C19542 VDD100.t98 VSS 0.00671f
C19543 VDD100.n369 VSS 0.0482f
C19544 VDD100.n370 VSS 0.0356f
C19545 VDD100.n371 VSS 0.0366f
C19546 VDD100.n372 VSS 0.0194f
C19547 VDD100.n373 VSS 0.0356f
C19548 VDD100.n374 VSS 0.0365f
C19549 VDD100.n375 VSS 0.0216f
C19550 VDD100.n376 VSS 0.031f
C19551 VDD100.n377 VSS 0.0288f
C19552 VDD100.n378 VSS 0.0216f
C19553 VDD100.n379 VSS 0.0554f
C19554 VDD100.n380 VSS 0.0443f
C19555 VDD100.n381 VSS 0.0317f
C19556 VDD100.t271 VSS 0.00626f
C19557 VDD100.n382 VSS 0.0288f
C19558 VDD100.n383 VSS 0.0216f
C19559 VDD100.n384 VSS 0.0335f
C19560 VDD100.t270 VSS 0.06f
C19561 VDD100.t466 VSS 0.0657f
C19562 VDD100.n385 VSS 0.0335f
C19563 VDD100.n386 VSS 0.0216f
C19564 VDD100.n387 VSS 0.0288f
C19565 VDD100.n388 VSS 0.031f
C19566 VDD100.n389 VSS 0.0216f
C19567 VDD100.t164 VSS 0.00257f
C19568 VDD100.n390 VSS 0.00257f
C19569 VDD100.n391 VSS 0.00562f
C19570 VDD100.t126 VSS 0.00626f
C19571 VDD100.n392 VSS 0.0273f
C19572 VDD100.n393 VSS 0.0256f
C19573 VDD100.n394 VSS 0.0194f
C19574 VDD100.n395 VSS 0.0335f
C19575 VDD100.t453 VSS 0.034f
C19576 VDD100.t163 VSS 0.0733f
C19577 VDD100.t125 VSS 0.06f
C19578 VDD100.n396 VSS 0.0335f
C19579 VDD100.t36 VSS 0.0288f
C19580 VDD100.n397 VSS 0.174f
C19581 VDD100.n398 VSS 0.0958f
C19582 VDD100.t461 VSS 0.0689f
C19583 VDD100.n399 VSS 0.0192f
C19584 VDD100.n400 VSS 0.00625f
C19585 VDD100.t458 VSS 0.0814f
C19586 VDD100.n401 VSS 0.0388f
C19587 VDD100.t63 VSS 0.00626f
C19588 VDD100.n402 VSS 0.00625f
C19589 VDD100.t62 VSS 0.0754f
C19590 VDD100.t298 VSS 0.0826f
C19591 VDD100.n403 VSS 0.0388f
C19592 VDD100.t273 VSS 0.00626f
C19593 VDD100.t310 VSS 0.00257f
C19594 VDD100.n404 VSS 0.00257f
C19595 VDD100.n405 VSS 0.00562f
C19596 VDD100.t272 VSS 0.0754f
C19597 VDD100.t309 VSS 0.0921f
C19598 VDD100.t372 VSS 0.0428f
C19599 VDD100.n406 VSS 0.0388f
C19600 VDD100.t336 VSS 0.00626f
C19601 VDD100.t444 VSS 0.00257f
C19602 VDD100.n407 VSS 0.00257f
C19603 VDD100.n408 VSS 0.00562f
C19604 VDD100.t335 VSS 0.0754f
C19605 VDD100.t443 VSS 0.0921f
C19606 VDD100.t473 VSS 0.0428f
C19607 VDD100.t80 VSS 0.0752f
C19608 VDD100.n409 VSS 0.0388f
C19609 VDD100.t81 VSS 0.00671f
C19610 VDD100.n410 VSS 0.0482f
C19611 VDD100.n411 VSS 0.0356f
C19612 VDD100.n412 VSS 0.0366f
C19613 VDD100.n413 VSS 0.0194f
C19614 VDD100.n414 VSS 0.0356f
C19615 VDD100.n415 VSS 0.0365f
C19616 VDD100.n416 VSS 0.0216f
C19617 VDD100.n417 VSS 0.031f
C19618 VDD100.n418 VSS 0.0288f
C19619 VDD100.n419 VSS 0.0216f
C19620 VDD100.n420 VSS 0.0554f
C19621 VDD100.n421 VSS 0.0393f
C19622 VDD100.n422 VSS 0.0317f
C19623 VDD100.t112 VSS 0.00626f
C19624 VDD100.n423 VSS 0.0288f
C19625 VDD100.n424 VSS 0.0216f
C19626 VDD100.n425 VSS 0.0335f
C19627 VDD100.t111 VSS 0.06f
C19628 VDD100.t301 VSS 0.0657f
C19629 VDD100.t307 VSS 0.0235f
C19630 VDD100.n426 VSS 0.0335f
C19631 VDD100.n427 VSS 0.0216f
C19632 VDD100.n428 VSS 0.0288f
C19633 VDD100.n429 VSS 0.031f
C19634 VDD100.t331 VSS 0.00626f
C19635 VDD100.n430 VSS 0.0273f
C19636 VDD100.n431 VSS 0.0216f
C19637 VDD100.n432 VSS 0.0335f
C19638 VDD100.t330 VSS 0.06f
C19639 VDD100.t410 VSS 0.0733f
C19640 VDD100.t470 VSS 0.0316f
C19641 VDD100.n433 VSS 0.0626f
C19642 VDD100.n434 VSS 0.061f
C19643 VDD100.n435 VSS 0.0243f
C19644 VDD100.t101 VSS 0.00626f
C19645 VDD100.t100 VSS 0.0582f
C19646 VDD100.t108 VSS 0.0918f
C19647 VDD100.n436 VSS 0.0793f
C19648 VDD100.t337 VSS 0.0738f
C19649 VDD100.t346 VSS 0.206f
C19650 VDD100.t469 VSS 0.00653f
C19651 VDD100.n437 VSS 0.0107f
C19652 VDD100.n438 VSS 0.0274f
C19653 VDD100.n439 VSS 0.0294f
C19654 VDD100.n440 VSS 0.0182f
C19655 VDD100.n441 VSS 0.0281f
C19656 VDD100.n442 VSS 0.0296f
C19657 VDD100.n443 VSS 0.0206f
C19658 VDD100.n444 VSS 0.00635f
C19659 VDD100.n445 VSS 0.034f
C19660 VDD100.n446 VSS 0.022f
C19661 VDD100.n447 VSS 0.0307f
C19662 VDD100.n448 VSS 0.0219f
C19663 VDD100.n449 VSS 0.0292f
C19664 VDD100.n450 VSS 0.022f
C19665 VDD100.n451 VSS 0.0307f
C19666 VDD100.n452 VSS 0.0219f
C19667 VDD100.n453 VSS 0.0292f
C19668 VDD100.n454 VSS 0.022f
C19669 VDD100.n455 VSS 0.0307f
C19670 VDD100.n456 VSS 0.0219f
C19671 VDD100.n457 VSS 0.0788f
C19672 VDD100.n458 VSS 0.00626f
C19673 VDD100.n459 VSS 0.0205f
C19674 VDD100.n460 VSS 0.0663f
C19675 VDD100.n461 VSS 0.0256f
C19676 VDD100.n462 VSS 0.0194f
C19677 VDD100.n463 VSS 0.0388f
C19678 VDD100.t420 VSS 0.0426f
C19679 VDD100.t437 VSS 0.0921f
C19680 VDD100.t135 VSS 0.0756f
C19681 VDD100.t34 VSS 0.0825f
C19682 VDD100.n464 VSS 0.0388f
C19683 VDD100.n465 VSS 0.0217f
C19684 VDD100.n466 VSS 0.031f
C19685 VDD100.n467 VSS 0.0288f
C19686 VDD100.t195 VSS 0.00625f
C19687 VDD100.n468 VSS 0.00626f
C19688 VDD100.n469 VSS 0.0288f
C19689 VDD100.n470 VSS 0.031f
C19690 VDD100.n471 VSS 0.0217f
C19691 VDD100.n472 VSS 0.0388f
C19692 VDD100.t194 VSS 0.0825f
C19693 VDD100.t387 VSS 0.0756f
C19694 VDD100.t435 VSS 0.0813f
C19695 VDD100.n473 VSS 0.0388f
C19696 VDD100.n474 VSS 0.0217f
C19697 VDD100.n475 VSS 0.0317f
C19698 VDD100.n476 VSS 0.0441f
C19699 VDD100.n477 VSS 0.0196f
C19700 VDD100.t405 VSS 0.0553f
C19701 VDD100.n478 VSS 0.0581f
C19702 VDD100.n479 VSS 0.0296f
C19703 VDD100.t246 VSS 0.00257f
C19704 VDD100.n480 VSS 0.00257f
C19705 VDD100.n481 VSS 0.00562f
C19706 VDD100.n482 VSS 0.00626f
C19707 VDD100.n483 VSS 0.0273f
C19708 VDD100.n484 VSS 0.0256f
C19709 VDD100.n485 VSS 0.0194f
C19710 VDD100.n486 VSS 0.0388f
C19711 VDD100.t245 VSS 0.0426f
C19712 VDD100.t129 VSS 0.0921f
C19713 VDD100.t17 VSS 0.0756f
C19714 VDD100.t6 VSS 0.0825f
C19715 VDD100.n487 VSS 0.0388f
C19716 VDD100.n488 VSS 0.0217f
C19717 VDD100.n489 VSS 0.031f
C19718 VDD100.n490 VSS 0.0288f
C19719 VDD100.t116 VSS 0.00625f
C19720 VDD100.n491 VSS 0.00626f
C19721 VDD100.n492 VSS 0.0288f
C19722 VDD100.n493 VSS 0.031f
C19723 VDD100.n494 VSS 0.0217f
C19724 VDD100.n495 VSS 0.0388f
C19725 VDD100.t115 VSS 0.0825f
C19726 VDD100.t338 VSS 0.0756f
C19727 VDD100.t127 VSS 0.0813f
C19728 VDD100.n496 VSS 0.0388f
C19729 VDD100.n497 VSS 0.0217f
C19730 VDD100.n498 VSS 0.0657f
C19731 VDD100.n499 VSS 0.00629f
C19732 VDD100.n500 VSS 0.00172f
C19733 VDD100.n501 VSS 0.0128f
C19734 VDD100.n502 VSS 0.0697f
C19735 VDD100.n503 VSS 0.0227f
C19736 VDD100.n504 VSS 0.0217f
C19737 VDD100.n505 VSS 0.0288f
C19738 VDD100.n506 VSS 0.031f
C19739 VDD100.n507 VSS 0.0217f
C19740 VDD100.n508 VSS 0.0364f
C19741 VDD100.n509 VSS 0.0357f
C19742 VDD100.n510 VSS 0.0194f
C19743 VDD100.n511 VSS 0.0366f
C19744 VDD100.n512 VSS 0.0357f
C19745 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n0 VSS 0.353f
C19746 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n1 VSS 0.227f
C19747 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t1 VSS 0.0191f
C19748 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t2 VSS 0.0157f
C19749 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n2 VSS 0.0157f
C19750 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n3 VSS 0.0378f
C19751 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t9 VSS 0.035f
C19752 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t11 VSS 0.0231f
C19753 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n4 VSS 0.0622f
C19754 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t3 VSS 0.0201f
C19755 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t15 VSS 0.0252f
C19756 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n5 VSS 0.0596f
C19757 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t16 VSS 0.0201f
C19758 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t13 VSS 0.0252f
C19759 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n6 VSS 0.0596f
C19760 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n7 VSS 1.06f
C19761 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n8 VSS 0.789f
C19762 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t4 VSS 0.0251f
C19763 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t8 VSS 0.0201f
C19764 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n9 VSS 0.0584f
C19765 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n10 VSS 0.362f
C19766 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t5 VSS 0.029f
C19767 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t12 VSS 0.0074f
C19768 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n11 VSS 0.048f
C19769 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t14 VSS 0.0231f
C19770 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t10 VSS 0.035f
C19771 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n12 VSS 0.0619f
C19772 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t7 VSS 0.0231f
C19773 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.t6 VSS 0.035f
C19774 CLK_div_93_mag_0.CLK_div_31_mag_0.Q1.n13 VSS 0.0619f
C19775 VDD99.t461 VSS 0.00692f
C19776 VDD99.n0 VSS 0.00693f
C19777 VDD99.n1 VSS 0.232f
C19778 VDD99.t234 VSS 0.00692f
C19779 VDD99.t95 VSS 0.0837f
C19780 VDD99.n2 VSS 0.00693f
C19781 VDD99.n3 VSS 0.226f
C19782 VDD99.t91 VSS 0.00692f
C19783 VDD99.t485 VSS 0.0475f
C19784 VDD99.n4 VSS 0.00693f
C19785 VDD99.n5 VSS 0.0273f
C19786 VDD99.n6 VSS 0.00698f
C19787 VDD99.t127 VSS 0.0613f
C19788 VDD99.n7 VSS 0.0643f
C19789 VDD99.n8 VSS 0.0925f
C19790 VDD99.n9 VSS 0.0069f
C19791 VDD99.n10 VSS 0.0225f
C19792 VDD99.t77 VSS 0.0544f
C19793 VDD99.t287 VSS 0.0625f
C19794 VDD99.t78 VSS 0.00692f
C19795 VDD99.n11 VSS 0.00693f
C19796 VDD99.n12 VSS 0.215f
C19797 VDD99.t434 VSS 0.00692f
C19798 VDD99.t190 VSS 0.0837f
C19799 VDD99.n13 VSS 0.199f
C19800 VDD99.n14 VSS 0.00693f
C19801 VDD99.t331 VSS 0.00692f
C19802 VDD99.n15 VSS 0.179f
C19803 VDD99.t471 VSS 0.0475f
C19804 VDD99.n16 VSS 0.00706f
C19805 VDD99.n17 VSS 0.00723f
C19806 VDD99.t502 VSS 0.0613f
C19807 VDD99.n18 VSS 0.0643f
C19808 VDD99.n19 VSS 0.215f
C19809 VDD99.t495 VSS 0.00285f
C19810 VDD99.n20 VSS 0.00285f
C19811 VDD99.n21 VSS 0.00622f
C19812 VDD99.n22 VSS 0.00693f
C19813 VDD99.n23 VSS 0.0242f
C19814 VDD99.n24 VSS 0.921f
C19815 VDD99.n25 VSS 0.0728f
C19816 VDD99.n26 VSS 0.0256f
C19817 VDD99.n27 VSS 0.0147f
C19818 VDD99.n28 VSS 0.043f
C19819 VDD99.t494 VSS 0.0472f
C19820 VDD99.t435 VSS 0.102f
C19821 VDD99.t411 VSS 0.0837f
C19822 VDD99.t330 VSS 0.0913f
C19823 VDD99.n29 VSS 0.043f
C19824 VDD99.n30 VSS 0.0186f
C19825 VDD99.n31 VSS 0.065f
C19826 VDD99.n32 VSS 0.0299f
C19827 VDD99.n33 VSS 0.0278f
C19828 VDD99.n34 VSS 0.0624f
C19829 VDD99.t283 VSS 0.00692f
C19830 VDD99.n35 VSS 0.00706f
C19831 VDD99.n36 VSS 0.0913f
C19832 VDD99.n37 VSS 0.0314f
C19833 VDD99.n38 VSS 0.024f
C19834 VDD99.n39 VSS 0.043f
C19835 VDD99.t282 VSS 0.0913f
C19836 VDD99.t284 VSS 0.0837f
C19837 VDD99.t433 VSS 0.09f
C19838 VDD99.n40 VSS 0.043f
C19839 VDD99.n41 VSS 0.024f
C19840 VDD99.n42 VSS 0.0313f
C19841 VDD99.t80 VSS 0.00692f
C19842 VDD99.t332 VSS 0.0837f
C19843 VDD99.n43 VSS 0.00693f
C19844 VDD99.t375 VSS 0.00285f
C19845 VDD99.n44 VSS 0.00285f
C19846 VDD99.n45 VSS 0.00622f
C19847 VDD99.n46 VSS 0.00693f
C19848 VDD99.n47 VSS 0.0405f
C19849 VDD99.t45 VSS 0.0835f
C19850 VDD99.n48 VSS 6.85e-19
C19851 VDD99.t510 VSS 0.00451f
C19852 VDD99.t48 VSS 0.00594f
C19853 VDD99.n49 VSS 0.0116f
C19854 VDD99.n50 VSS 0.0772f
C19855 VDD99.n51 VSS 0.0762f
C19856 VDD99.t511 VSS 0.00451f
C19857 VDD99.t44 VSS 0.00583f
C19858 VDD99.n52 VSS 0.00554f
C19859 VDD99.n53 VSS 0.00618f
C19860 VDD99.n54 VSS 9.79e-19
C19861 VDD99.n55 VSS 0.00517f
C19862 VDD99.n56 VSS 0.00647f
C19863 VDD99.n57 VSS 0.0162f
C19864 VDD99.t493 VSS 0.00285f
C19865 VDD99.n58 VSS 0.00285f
C19866 VDD99.n59 VSS 0.00622f
C19867 VDD99.n60 VSS 0.0395f
C19868 VDD99.n61 VSS 0.0396f
C19869 VDD99.n62 VSS 0.043f
C19870 VDD99.t492 VSS 0.0472f
C19871 VDD99.t81 VSS 0.102f
C19872 VDD99.t308 VSS 0.0837f
C19873 VDD99.t193 VSS 0.102f
C19874 VDD99.t374 VSS 0.0472f
C19875 VDD99.n63 VSS 0.043f
C19876 VDD99.n64 VSS 0.0214f
C19877 VDD99.n65 VSS 0.0395f
C19878 VDD99.n66 VSS 0.0403f
C19879 VDD99.t281 VSS 0.00692f
C19880 VDD99.n67 VSS 0.00693f
C19881 VDD99.n68 VSS 0.0318f
C19882 VDD99.n69 VSS 0.0343f
C19883 VDD99.n70 VSS 0.024f
C19884 VDD99.n71 VSS 0.043f
C19885 VDD99.t280 VSS 0.0913f
C19886 VDD99.t335 VSS 0.0837f
C19887 VDD99.t79 VSS 0.09f
C19888 VDD99.n72 VSS 0.043f
C19889 VDD99.n73 VSS 0.024f
C19890 VDD99.n74 VSS 0.0598f
C19891 VDD99.n75 VSS 0.0069f
C19892 VDD99.n76 VSS 0.00693f
C19893 VDD99.n77 VSS 0.0305f
C19894 VDD99.t499 VSS 0.0613f
C19895 VDD99.n78 VSS 0.016f
C19896 VDD99.t145 VSS 0.0913f
C19897 VDD99.n79 VSS 0.00693f
C19898 VDD99.t491 VSS 0.00285f
C19899 VDD99.n80 VSS 0.00285f
C19900 VDD99.n81 VSS 0.00622f
C19901 VDD99.n82 VSS 0.054f
C19902 VDD99.n83 VSS 0.0224f
C19903 VDD99.n84 VSS 0.0302f
C19904 VDD99.t146 VSS 0.00692f
C19905 VDD99.n85 VSS 0.00693f
C19906 VDD99.t296 VSS 0.0837f
C19907 VDD99.n86 VSS 0.043f
C19908 VDD99.t36 VSS 0.00692f
C19909 VDD99.n87 VSS 0.00693f
C19910 VDD99.t35 VSS 0.0913f
C19911 VDD99.t253 VSS 0.0837f
C19912 VDD99.t469 VSS 0.09f
C19913 VDD99.n88 VSS 0.043f
C19914 VDD99.t470 VSS 0.00692f
C19915 VDD99.t116 VSS 0.00692f
C19916 VDD99.t147 VSS 0.0837f
C19917 VDD99.n89 VSS 0.00693f
C19918 VDD99.t377 VSS 0.00285f
C19919 VDD99.n90 VSS 0.00285f
C19920 VDD99.n91 VSS 0.00622f
C19921 VDD99.n92 VSS 0.00693f
C19922 VDD99.n93 VSS 0.0405f
C19923 VDD99.t49 VSS 0.0835f
C19924 VDD99.n94 VSS 0.00743f
C19925 VDD99.t489 VSS 0.00285f
C19926 VDD99.n95 VSS 0.00285f
C19927 VDD99.n96 VSS 0.00622f
C19928 VDD99.n97 VSS 0.0395f
C19929 VDD99.n98 VSS 0.0534f
C19930 VDD99.n99 VSS 0.043f
C19931 VDD99.t488 VSS 0.0472f
C19932 VDD99.t117 VSS 0.102f
C19933 VDD99.t240 VSS 0.0837f
C19934 VDD99.t293 VSS 0.102f
C19935 VDD99.t376 VSS 0.0472f
C19936 VDD99.n100 VSS 0.043f
C19937 VDD99.n101 VSS 0.0214f
C19938 VDD99.n102 VSS 0.0395f
C19939 VDD99.n103 VSS 0.0403f
C19940 VDD99.t34 VSS 0.00692f
C19941 VDD99.n104 VSS 0.00693f
C19942 VDD99.n105 VSS 0.0318f
C19943 VDD99.n106 VSS 0.0343f
C19944 VDD99.n107 VSS 0.024f
C19945 VDD99.n108 VSS 0.043f
C19946 VDD99.t33 VSS 0.0913f
C19947 VDD99.t13 VSS 0.0837f
C19948 VDD99.t115 VSS 0.09f
C19949 VDD99.n109 VSS 0.043f
C19950 VDD99.n110 VSS 0.024f
C19951 VDD99.n111 VSS 0.0652f
C19952 VDD99.n112 VSS 0.0741f
C19953 VDD99.n113 VSS 0.024f
C19954 VDD99.n114 VSS 0.0318f
C19955 VDD99.n115 VSS 0.0343f
C19956 VDD99.n116 VSS 0.024f
C19957 VDD99.n117 VSS 0.0318f
C19958 VDD99.n118 VSS 0.0343f
C19959 VDD99.n119 VSS 0.024f
C19960 VDD99.n120 VSS 0.043f
C19961 VDD99.t403 VSS 0.0837f
C19962 VDD99.t466 VSS 0.102f
C19963 VDD99.t490 VSS 0.0472f
C19964 VDD99.n121 VSS 0.043f
C19965 VDD99.t84 VSS 0.0475f
C19966 VDD99.n122 VSS 0.0643f
C19967 VDD99.n123 VSS 0.0217f
C19968 VDD99.n124 VSS 0.0414f
C19969 VDD99.n125 VSS 0.068f
C19970 VDD99.n126 VSS 0.253f
C19971 VDD99.n127 VSS 0.199f
C19972 VDD99.n128 VSS 0.0544f
C19973 VDD99.t496 VSS 0.0835f
C19974 VDD99.n129 VSS 0.043f
C19975 VDD99.n130 VSS 0.0464f
C19976 VDD99.n131 VSS 0.0959f
C19977 VDD99.n132 VSS 0.00869f
C19978 VDD99.n133 VSS 0.0166f
C19979 VDD99.n134 VSS 0.0975f
C19980 VDD99.n135 VSS 0.069f
C19981 VDD99.n136 VSS 0.108f
C19982 VDD99.t8 VSS 0.0589f
C19983 VDD99.t219 VSS 0.0616f
C19984 VDD99.n137 VSS 0.0712f
C19985 VDD99.t120 VSS 0.062f
C19986 VDD99.n138 VSS 0.0418f
C19987 VDD99.n139 VSS 0.0721f
C19988 VDD99.n140 VSS 0.169f
C19989 VDD99.n141 VSS 0.2f
C19990 VDD99.n142 VSS 0.194f
C19991 VDD99.t135 VSS 0.00285f
C19992 VDD99.n143 VSS 0.00285f
C19993 VDD99.n144 VSS 0.00622f
C19994 VDD99.n145 VSS 0.211f
C19995 VDD99.n146 VSS 0.00693f
C19996 VDD99.n147 VSS 0.0213f
C19997 VDD99.n148 VSS 0.0708f
C19998 VDD99.n149 VSS 0.0245f
C19999 VDD99.n150 VSS 0.0699f
C20000 VDD99.n151 VSS 0.0161f
C20001 VDD99.n152 VSS 0.043f
C20002 VDD99.t134 VSS 0.0472f
C20003 VDD99.t235 VSS 0.102f
C20004 VDD99.t92 VSS 0.0837f
C20005 VDD99.t90 VSS 0.0913f
C20006 VDD99.n153 VSS 0.043f
C20007 VDD99.n154 VSS 0.024f
C20008 VDD99.n155 VSS 0.0252f
C20009 VDD99.n156 VSS 0.0681f
C20010 VDD99.n157 VSS 0.0281f
C20011 VDD99.t30 VSS 0.00692f
C20012 VDD99.n158 VSS 0.00693f
C20013 VDD99.n159 VSS 0.0265f
C20014 VDD99.n160 VSS 0.0681f
C20015 VDD99.n161 VSS 0.0268f
C20016 VDD99.n162 VSS 0.024f
C20017 VDD99.n163 VSS 0.043f
C20018 VDD99.t29 VSS 0.0913f
C20019 VDD99.t65 VSS 0.0837f
C20020 VDD99.t233 VSS 0.09f
C20021 VDD99.n164 VSS 0.043f
C20022 VDD99.n165 VSS 0.024f
C20023 VDD99.n166 VSS 0.0265f
C20024 VDD99.t456 VSS 0.00692f
C20025 VDD99.t87 VSS 0.0837f
C20026 VDD99.n167 VSS 0.00693f
C20027 VDD99.t359 VSS 0.00285f
C20028 VDD99.n168 VSS 0.00285f
C20029 VDD99.n169 VSS 0.00622f
C20030 VDD99.n170 VSS 0.00693f
C20031 VDD99.n171 VSS 0.0405f
C20032 VDD99.t41 VSS 0.0835f
C20033 VDD99.n172 VSS 9.33e-19
C20034 VDD99.t515 VSS 0.00451f
C20035 VDD99.t52 VSS 0.00594f
C20036 VDD99.n173 VSS 0.0116f
C20037 VDD99.n174 VSS 0.0772f
C20038 VDD99.t513 VSS 0.00451f
C20039 VDD99.n175 VSS 0.00618f
C20040 VDD99.t40 VSS 0.00583f
C20041 VDD99.n176 VSS 0.00554f
C20042 VDD99.n177 VSS 0.0758f
C20043 VDD99.n178 VSS 0.00335f
C20044 VDD99.n179 VSS 0.00647f
C20045 VDD99.n180 VSS 0.0182f
C20046 VDD99.t133 VSS 0.00285f
C20047 VDD99.n181 VSS 0.00285f
C20048 VDD99.n182 VSS 0.00622f
C20049 VDD99.n183 VSS 0.0395f
C20050 VDD99.n184 VSS 0.0396f
C20051 VDD99.n185 VSS 0.043f
C20052 VDD99.t132 VSS 0.0472f
C20053 VDD99.t452 VSS 0.102f
C20054 VDD99.t311 VSS 0.0837f
C20055 VDD99.t98 VSS 0.102f
C20056 VDD99.t358 VSS 0.0472f
C20057 VDD99.n186 VSS 0.043f
C20058 VDD99.n187 VSS 0.0214f
C20059 VDD99.n188 VSS 0.0395f
C20060 VDD99.n189 VSS 0.0403f
C20061 VDD99.t32 VSS 0.00692f
C20062 VDD99.n190 VSS 0.00693f
C20063 VDD99.n191 VSS 0.0318f
C20064 VDD99.n192 VSS 0.0343f
C20065 VDD99.n193 VSS 0.024f
C20066 VDD99.n194 VSS 0.043f
C20067 VDD99.t31 VSS 0.0913f
C20068 VDD99.t230 VSS 0.0837f
C20069 VDD99.t455 VSS 0.09f
C20070 VDD99.n195 VSS 0.043f
C20071 VDD99.n196 VSS 0.024f
C20072 VDD99.n197 VSS 0.0613f
C20073 VDD99.n198 VSS 0.0069f
C20074 VDD99.n199 VSS 0.00693f
C20075 VDD99.n200 VSS 0.0305f
C20076 VDD99.t121 VSS 0.0613f
C20077 VDD99.n201 VSS 0.016f
C20078 VDD99.t110 VSS 0.0913f
C20079 VDD99.n202 VSS 0.00693f
C20080 VDD99.t131 VSS 0.00285f
C20081 VDD99.n203 VSS 0.00285f
C20082 VDD99.n204 VSS 0.00622f
C20083 VDD99.n205 VSS 0.054f
C20084 VDD99.n206 VSS 0.0224f
C20085 VDD99.n207 VSS 0.0302f
C20086 VDD99.t111 VSS 0.00692f
C20087 VDD99.n208 VSS 0.00693f
C20088 VDD99.t302 VSS 0.0837f
C20089 VDD99.n209 VSS 0.043f
C20090 VDD99.t277 VSS 0.00692f
C20091 VDD99.n210 VSS 0.00693f
C20092 VDD99.t276 VSS 0.0913f
C20093 VDD99.t305 VSS 0.0837f
C20094 VDD99.t480 VSS 0.09f
C20095 VDD99.n211 VSS 0.043f
C20096 VDD99.t481 VSS 0.00692f
C20097 VDD99.t479 VSS 0.00692f
C20098 VDD99.t112 VSS 0.0837f
C20099 VDD99.n212 VSS 0.00693f
C20100 VDD99.t361 VSS 0.00285f
C20101 VDD99.n213 VSS 0.00285f
C20102 VDD99.n214 VSS 0.00622f
C20103 VDD99.n215 VSS 0.00693f
C20104 VDD99.n216 VSS 0.0405f
C20105 VDD99.t53 VSS 0.0835f
C20106 VDD99.n217 VSS 0.00743f
C20107 VDD99.t137 VSS 0.00285f
C20108 VDD99.n218 VSS 0.00285f
C20109 VDD99.n219 VSS 0.00622f
C20110 VDD99.n220 VSS 0.0395f
C20111 VDD99.n221 VSS 0.0534f
C20112 VDD99.n222 VSS 0.043f
C20113 VDD99.t136 VSS 0.0472f
C20114 VDD99.t474 VSS 0.102f
C20115 VDD99.t60 VSS 0.0837f
C20116 VDD99.t299 VSS 0.102f
C20117 VDD99.t360 VSS 0.0472f
C20118 VDD99.n223 VSS 0.043f
C20119 VDD99.n224 VSS 0.0214f
C20120 VDD99.n225 VSS 0.0395f
C20121 VDD99.n226 VSS 0.0403f
C20122 VDD99.t279 VSS 0.00692f
C20123 VDD99.n227 VSS 0.00693f
C20124 VDD99.n228 VSS 0.0318f
C20125 VDD99.n229 VSS 0.0343f
C20126 VDD99.n230 VSS 0.024f
C20127 VDD99.n231 VSS 0.043f
C20128 VDD99.t278 VSS 0.0913f
C20129 VDD99.t26 VSS 0.0837f
C20130 VDD99.t478 VSS 0.09f
C20131 VDD99.n232 VSS 0.043f
C20132 VDD99.n233 VSS 0.024f
C20133 VDD99.n234 VSS 0.0652f
C20134 VDD99.n235 VSS 0.0741f
C20135 VDD99.n236 VSS 0.024f
C20136 VDD99.n237 VSS 0.0318f
C20137 VDD99.n238 VSS 0.0343f
C20138 VDD99.n239 VSS 0.024f
C20139 VDD99.n240 VSS 0.0318f
C20140 VDD99.n241 VSS 0.0343f
C20141 VDD99.n242 VSS 0.024f
C20142 VDD99.n243 VSS 0.043f
C20143 VDD99.t273 VSS 0.0837f
C20144 VDD99.t482 VSS 0.102f
C20145 VDD99.t130 VSS 0.0472f
C20146 VDD99.n244 VSS 0.043f
C20147 VDD99.t457 VSS 0.0475f
C20148 VDD99.n245 VSS 0.0643f
C20149 VDD99.n246 VSS 0.0217f
C20150 VDD99.n247 VSS 0.0435f
C20151 VDD99.n248 VSS 0.0693f
C20152 VDD99.n249 VSS 0.278f
C20153 VDD99.n250 VSS 0.213f
C20154 VDD99.n251 VSS 0.0544f
C20155 VDD99.t124 VSS 0.0835f
C20156 VDD99.t460 VSS 0.0544f
C20157 VDD99.n252 VSS 0.043f
C20158 VDD99.n253 VSS 0.0464f
C20159 VDD99.n254 VSS 0.0959f
C20160 VDD99.t68 VSS 0.0625f
C20161 VDD99.n255 VSS 0.108f
C20162 VDD99.n256 VSS 0.00869f
C20163 VDD99.n257 VSS 0.0166f
C20164 VDD99.t406 VSS 0.0589f
C20165 VDD99.n258 VSS 0.0418f
C20166 VDD99.n259 VSS 0.0069f
C20167 VDD99.t477 VSS 0.062f
C20168 VDD99.t338 VSS 0.0616f
C20169 VDD99.n260 VSS 0.0712f
C20170 VDD99.n261 VSS 0.0225f
C20171 VDD99.t432 VSS 0.00693f
C20172 VDD99.n262 VSS 0.00692f
C20173 VDD99.n263 VSS 0.034f
C20174 VDD99.t409 VSS 0.0815f
C20175 VDD99.t431 VSS 0.067f
C20176 VDD99.t351 VSS 0.0335f
C20177 VDD99.t410 VSS 0.0069f
C20178 VDD99.n264 VSS 0.0244f
C20179 VDD99.n265 VSS 0.0672f
C20180 VDD99.n266 VSS 0.0487f
C20181 VDD99.n267 VSS 0.0309f
C20182 VDD99.t244 VSS 0.0069f
C20183 VDD99.n268 VSS 0.0316f
C20184 VDD99.t243 VSS 0.0652f
C20185 VDD99.n269 VSS 0.0739f
C20186 VDD99.t292 VSS 0.0774f
C20187 VDD99.t256 VSS 0.0777f
C20188 VDD99.n270 VSS 0.0488f
C20189 VDD99.t257 VSS 0.0182f
C20190 VDD99.n271 VSS 0.105f
C20191 VDD99.t109 VSS 0.0069f
C20192 VDD99.n272 VSS 0.0318f
C20193 VDD99.t108 VSS 0.0652f
C20194 VDD99.n273 VSS 0.0739f
C20195 VDD99.t176 VSS 0.0774f
C20196 VDD99.t106 VSS 0.0777f
C20197 VDD99.n274 VSS 0.0488f
C20198 VDD99.t107 VSS 0.0181f
C20199 VDD99.n275 VSS 0.106f
C20200 VDD99.t451 VSS 0.00661f
C20201 VDD99.t57 VSS 0.0144f
C20202 VDD99.n276 VSS 0.205f
C20203 VDD99.t139 VSS 0.00693f
C20204 VDD99.t159 VSS 0.00285f
C20205 VDD99.n277 VSS 0.00285f
C20206 VDD99.n278 VSS 0.00622f
C20207 VDD99.t424 VSS 0.00693f
C20208 VDD99.n279 VSS 0.00692f
C20209 VDD99.n280 VSS 0.163f
C20210 VDD99.t143 VSS 0.0815f
C20211 VDD99.t423 VSS 0.067f
C20212 VDD99.t140 VSS 0.0335f
C20213 VDD99.t144 VSS 0.00871f
C20214 VDD99.t72 VSS 0.0151f
C20215 VDD99.t415 VSS 0.0134f
C20216 VDD99.n281 VSS 0.123f
C20217 VDD99.t414 VSS 0.0456f
C20218 VDD99.t75 VSS 0.0886f
C20219 VDD99.t76 VSS 0.0144f
C20220 VDD99.n282 VSS -0.211f
C20221 VDD99.t344 VSS 0.00693f
C20222 VDD99.t343 VSS 0.0816f
C20223 VDD99.n283 VSS 0.0538f
C20224 VDD99.t345 VSS 0.169f
C20225 VDD99.t37 VSS 0.0561f
C20226 VDD99.t342 VSS 0.0408f
C20227 VDD99.n284 VSS 0.0381f
C20228 VDD99.n285 VSS 0.0651f
C20229 VDD99.t341 VSS 0.179f
C20230 VDD99.n286 VSS 0.101f
C20231 VDD99.n287 VSS 0.159f
C20232 VDD99.n288 VSS 0.0922f
C20233 VDD99.n289 VSS 0.0976f
C20234 VDD99.t71 VSS 0.0485f
C20235 VDD99.n290 VSS 0.0645f
C20236 VDD99.n291 VSS 0.2f
C20237 VDD99.n292 VSS 0.0672f
C20238 VDD99.n293 VSS 0.0961f
C20239 VDD99.n294 VSS 0.205f
C20240 VDD99.n295 VSS 0.216f
C20241 VDD99.t158 VSS 0.067f
C20242 VDD99.t138 VSS 0.067f
C20243 VDD99.t261 VSS 0.0505f
C20244 VDD99.n296 VSS 0.0521f
C20245 VDD99.n297 VSS 0.232f
C20246 VDD99.t56 VSS 0.0687f
C20247 VDD99.t450 VSS 0.0825f
C20248 VDD99.n298 VSS 0.0717f
C20249 VDD99.n299 VSS 0.117f
C20250 VDD99.n300 VSS 0.128f
C20251 VDD99.t439 VSS 0.00285f
C20252 VDD99.n301 VSS 0.00285f
C20253 VDD99.n302 VSS 0.00622f
C20254 VDD99.n303 VSS 0.0267f
C20255 VDD99.t198 VSS 0.0915f
C20256 VDD99.n304 VSS 0.00692f
C20257 VDD99.t396 VSS 0.00693f
C20258 VDD99.n305 VSS 0.00692f
C20259 VDD99.n306 VSS 0.0378f
C20260 VDD99.t440 VSS 0.0902f
C20261 VDD99.n307 VSS 0.00692f
C20262 VDD99.n308 VSS 0.00692f
C20263 VDD99.t443 VSS 0.0902f
C20264 VDD99.n309 VSS 0.043f
C20265 VDD99.t329 VSS 0.00693f
C20266 VDD99.n310 VSS 0.00692f
C20267 VDD99.t328 VSS 0.0835f
C20268 VDD99.t0 VSS 0.0915f
C20269 VDD99.n311 VSS 0.043f
C20270 VDD99.t197 VSS 0.00693f
C20271 VDD99.t394 VSS 0.00285f
C20272 VDD99.n312 VSS 0.00285f
C20273 VDD99.n313 VSS 0.00622f
C20274 VDD99.t196 VSS 0.0835f
C20275 VDD99.t393 VSS 0.102f
C20276 VDD99.t368 VSS 0.0474f
C20277 VDD99.n314 VSS 0.043f
C20278 VDD99.t392 VSS 0.00693f
C20279 VDD99.t449 VSS 0.00285f
C20280 VDD99.n315 VSS 0.00285f
C20281 VDD99.n316 VSS 0.00622f
C20282 VDD99.t391 VSS 0.0835f
C20283 VDD99.t448 VSS 0.102f
C20284 VDD99.t155 VSS 0.0474f
C20285 VDD99.t464 VSS 0.0833f
C20286 VDD99.n317 VSS 0.043f
C20287 VDD99.t465 VSS 0.00743f
C20288 VDD99.n318 VSS 0.0533f
C20289 VDD99.n319 VSS 0.0395f
C20290 VDD99.n320 VSS 0.0405f
C20291 VDD99.n321 VSS 0.0215f
C20292 VDD99.n322 VSS 0.0395f
C20293 VDD99.n323 VSS 0.0404f
C20294 VDD99.n324 VSS 0.0239f
C20295 VDD99.n325 VSS 0.0343f
C20296 VDD99.n326 VSS 0.0319f
C20297 VDD99.n327 VSS 0.0239f
C20298 VDD99.n328 VSS 0.0601f
C20299 VDD99.t154 VSS 0.0069f
C20300 VDD99.t388 VSS 0.00693f
C20301 VDD99.n329 VSS 0.0401f
C20302 VDD99.t153 VSS 0.0611f
C20303 VDD99.t181 VSS 0.0474f
C20304 VDD99.t172 VSS 0.00285f
C20305 VDD99.n330 VSS 0.00285f
C20306 VDD99.n331 VSS 0.00622f
C20307 VDD99.t239 VSS 0.00693f
C20308 VDD99.n332 VSS 0.00692f
C20309 VDD99.n333 VSS 0.0375f
C20310 VDD99.t222 VSS 0.0915f
C20311 VDD99.n334 VSS 0.00692f
C20312 VDD99.t202 VSS 0.00693f
C20313 VDD99.n335 VSS 0.00692f
C20314 VDD99.n336 VSS 0.00692f
C20315 VDD99.t425 VSS 0.0902f
C20316 VDD99.n337 VSS 0.043f
C20317 VDD99.t229 VSS 0.00693f
C20318 VDD99.n338 VSS 0.00692f
C20319 VDD99.t228 VSS 0.0835f
C20320 VDD99.t225 VSS 0.0915f
C20321 VDD99.n339 VSS 0.043f
C20322 VDD99.t386 VSS 0.00693f
C20323 VDD99.t381 VSS 0.00285f
C20324 VDD99.n340 VSS 0.00285f
C20325 VDD99.n341 VSS 0.00622f
C20326 VDD99.t385 VSS 0.0835f
C20327 VDD99.t380 VSS 0.102f
C20328 VDD99.t362 VSS 0.0474f
C20329 VDD99.n342 VSS 0.043f
C20330 VDD99.t291 VSS 0.00693f
C20331 VDD99.t422 VSS 0.00285f
C20332 VDD99.n343 VSS 0.00285f
C20333 VDD99.n344 VSS 0.00622f
C20334 VDD99.t290 VSS 0.0835f
C20335 VDD99.t421 VSS 0.102f
C20336 VDD99.t168 VSS 0.0474f
C20337 VDD99.t389 VSS 0.0833f
C20338 VDD99.n345 VSS 0.043f
C20339 VDD99.t390 VSS 0.00743f
C20340 VDD99.n346 VSS 0.0533f
C20341 VDD99.n347 VSS 0.0395f
C20342 VDD99.n348 VSS 0.0405f
C20343 VDD99.n349 VSS 0.0215f
C20344 VDD99.n350 VSS 0.0395f
C20345 VDD99.n351 VSS 0.0404f
C20346 VDD99.n352 VSS 0.0239f
C20347 VDD99.n353 VSS 0.0343f
C20348 VDD99.n354 VSS 0.0319f
C20349 VDD99.n355 VSS 0.0239f
C20350 VDD99.n356 VSS 0.0814f
C20351 VDD99.t180 VSS 0.0069f
C20352 VDD99.t400 VSS 0.00693f
C20353 VDD99.n357 VSS 0.0408f
C20354 VDD99.t179 VSS 0.0611f
C20355 VDD99.t165 VSS 0.0474f
C20356 VDD99.t327 VSS 0.00285f
C20357 VDD99.n358 VSS 0.00285f
C20358 VDD99.n359 VSS 0.00622f
C20359 VDD99.t402 VSS 0.00693f
C20360 VDD99.n360 VSS 0.00692f
C20361 VDD99.n361 VSS 0.0381f
C20362 VDD99.t211 VSS 0.0915f
C20363 VDD99.n362 VSS 0.00692f
C20364 VDD99.t272 VSS 0.00693f
C20365 VDD99.n363 VSS 0.00692f
C20366 VDD99.n364 VSS 0.00692f
C20367 VDD99.t258 VSS 0.0902f
C20368 VDD99.n365 VSS 0.043f
C20369 VDD99.t64 VSS 0.00693f
C20370 VDD99.n366 VSS 0.00692f
C20371 VDD99.t63 VSS 0.0835f
C20372 VDD99.t208 VSS 0.0915f
C20373 VDD99.n367 VSS 0.043f
C20374 VDD99.t218 VSS 0.00693f
C20375 VDD99.t506 VSS 0.00285f
C20376 VDD99.n368 VSS 0.00285f
C20377 VDD99.n369 VSS 0.00622f
C20378 VDD99.t217 VSS 0.0835f
C20379 VDD99.t505 VSS 0.102f
C20380 VDD99.t371 VSS 0.0474f
C20381 VDD99.n370 VSS 0.043f
C20382 VDD99.t7 VSS 0.00693f
C20383 VDD99.t265 VSS 0.00285f
C20384 VDD99.n371 VSS 0.00285f
C20385 VDD99.n372 VSS 0.00622f
C20386 VDD99.t6 VSS 0.0835f
C20387 VDD99.t264 VSS 0.102f
C20388 VDD99.t150 VSS 0.0474f
C20389 VDD99.t397 VSS 0.0833f
C20390 VDD99.n373 VSS 0.043f
C20391 VDD99.t398 VSS 0.00743f
C20392 VDD99.n374 VSS 0.0533f
C20393 VDD99.n375 VSS 0.0395f
C20394 VDD99.n376 VSS 0.0405f
C20395 VDD99.n377 VSS 0.0215f
C20396 VDD99.n378 VSS 0.0395f
C20397 VDD99.n379 VSS 0.0404f
C20398 VDD99.n380 VSS 0.0239f
C20399 VDD99.n381 VSS 0.0343f
C20400 VDD99.n382 VSS 0.0319f
C20401 VDD99.n383 VSS 0.0239f
C20402 VDD99.n384 VSS 0.0817f
C20403 VDD99.n385 VSS 0.0941f
C20404 VDD99.t323 VSS 0.0902f
C20405 VDD99.t271 VSS 0.0835f
C20406 VDD99.n386 VSS 0.043f
C20407 VDD99.n387 VSS 0.0256f
C20408 VDD99.n388 VSS 0.0353f
C20409 VDD99.n389 VSS 0.0381f
C20410 VDD99.t508 VSS 0.00693f
C20411 VDD99.n390 VSS 0.0353f
C20412 VDD99.n391 VSS 0.0256f
C20413 VDD99.n392 VSS 0.043f
C20414 VDD99.t507 VSS 0.0835f
C20415 VDD99.t214 VSS 0.0915f
C20416 VDD99.t326 VSS 0.102f
C20417 VDD99.t401 VSS 0.0835f
C20418 VDD99.n393 VSS 0.043f
C20419 VDD99.n394 VSS 0.0256f
C20420 VDD99.n395 VSS 0.0333f
C20421 VDD99.n396 VSS 0.0316f
C20422 VDD99.n397 VSS 0.0227f
C20423 VDD99.n398 VSS 0.043f
C20424 VDD99.t399 VSS 0.0474f
C20425 VDD99.n399 VSS 0.0643f
C20426 VDD99.n400 VSS 0.0387f
C20427 VDD99.n401 VSS 0.0432f
C20428 VDD99.n402 VSS 0.0386f
C20429 VDD99.t173 VSS 0.0902f
C20430 VDD99.t201 VSS 0.0835f
C20431 VDD99.n403 VSS 0.043f
C20432 VDD99.n404 VSS 0.0253f
C20433 VDD99.n405 VSS 0.0347f
C20434 VDD99.n406 VSS 0.0375f
C20435 VDD99.t379 VSS 0.00693f
C20436 VDD99.n407 VSS 0.0347f
C20437 VDD99.n408 VSS 0.0253f
C20438 VDD99.n409 VSS 0.043f
C20439 VDD99.t378 VSS 0.0835f
C20440 VDD99.t382 VSS 0.0915f
C20441 VDD99.t171 VSS 0.102f
C20442 VDD99.t238 VSS 0.0835f
C20443 VDD99.n410 VSS 0.043f
C20444 VDD99.n411 VSS 0.0253f
C20445 VDD99.n412 VSS 0.0328f
C20446 VDD99.n413 VSS 0.0311f
C20447 VDD99.n414 VSS 0.0225f
C20448 VDD99.n415 VSS 0.043f
C20449 VDD99.t387 VSS 0.0474f
C20450 VDD99.n416 VSS 0.0643f
C20451 VDD99.n417 VSS 0.0371f
C20452 VDD99.n418 VSS 0.0609f
C20453 VDD99.n419 VSS 0.037f
C20454 VDD99.t59 VSS 0.00693f
C20455 VDD99.n420 VSS 0.035f
C20456 VDD99.n421 VSS 0.0255f
C20457 VDD99.n422 VSS 0.043f
C20458 VDD99.t58 VSS 0.0835f
C20459 VDD99.t3 VSS 0.0915f
C20460 VDD99.t395 VSS 0.0835f
C20461 VDD99.n423 VSS 0.043f
C20462 VDD99.n424 VSS 0.0255f
C20463 VDD99.n425 VSS 0.035f
C20464 VDD99.n426 VSS 0.0378f
C20465 VDD99.t417 VSS 0.00693f
C20466 VDD99.n427 VSS 0.033f
C20467 VDD99.n428 VSS 0.0255f
C20468 VDD99.n429 VSS 0.043f
C20469 VDD99.t416 VSS 0.0835f
C20470 VDD99.t438 VSS 0.102f
C20471 VDD99.t187 VSS 0.0474f
C20472 VDD99.n430 VSS 0.043f
C20473 VDD99.t463 VSS 0.00693f
C20474 VDD99.t462 VSS 0.0474f
C20475 VDD99.t177 VSS 0.0611f
C20476 VDD99.n431 VSS 0.0643f
C20477 VDD99.t178 VSS 0.0069f
C20478 VDD99.n432 VSS 0.00692f
C20479 VDD99.t346 VSS 0.0902f
C20480 VDD99.n433 VSS 0.043f
C20481 VDD99.t252 VSS 0.00693f
C20482 VDD99.n434 VSS 0.00692f
C20483 VDD99.t251 VSS 0.0835f
C20484 VDD99.t248 VSS 0.0915f
C20485 VDD99.n435 VSS 0.043f
C20486 VDD99.t315 VSS 0.00693f
C20487 VDD99.t320 VSS 0.00285f
C20488 VDD99.n436 VSS 0.00285f
C20489 VDD99.n437 VSS 0.00622f
C20490 VDD99.t314 VSS 0.0835f
C20491 VDD99.t319 VSS 0.102f
C20492 VDD99.t365 VSS 0.0474f
C20493 VDD99.n438 VSS 0.043f
C20494 VDD99.t25 VSS 0.00693f
C20495 VDD99.t350 VSS 0.00285f
C20496 VDD99.n439 VSS 0.00285f
C20497 VDD99.n440 VSS 0.00622f
C20498 VDD99.t24 VSS 0.0835f
C20499 VDD99.t349 VSS 0.102f
C20500 VDD99.t184 VSS 0.0474f
C20501 VDD99.t22 VSS 0.0833f
C20502 VDD99.n441 VSS 0.043f
C20503 VDD99.t23 VSS 0.00743f
C20504 VDD99.n442 VSS 0.0533f
C20505 VDD99.n443 VSS 0.0395f
C20506 VDD99.n444 VSS 0.0405f
C20507 VDD99.n445 VSS 0.0215f
C20508 VDD99.n446 VSS 0.0395f
C20509 VDD99.n447 VSS 0.0404f
C20510 VDD99.n448 VSS 0.0239f
C20511 VDD99.n449 VSS 0.0343f
C20512 VDD99.n450 VSS 0.0319f
C20513 VDD99.n451 VSS 0.0239f
C20514 VDD99.n452 VSS 0.0601f
C20515 VDD99.n453 VSS 0.00692f
C20516 VDD99.t101 VSS 0.0902f
C20517 VDD99.n454 VSS 0.043f
C20518 VDD99.t357 VSS 0.00693f
C20519 VDD99.n455 VSS 0.00692f
C20520 VDD99.t356 VSS 0.0835f
C20521 VDD99.t245 VSS 0.0915f
C20522 VDD99.n456 VSS 0.043f
C20523 VDD99.t322 VSS 0.00693f
C20524 VDD99.n457 VSS 0.00692f
C20525 VDD99.t321 VSS 0.0835f
C20526 VDD99.t316 VSS 0.0915f
C20527 VDD99.n458 VSS 0.043f
C20528 VDD99.t17 VSS 0.00693f
C20529 VDD99.t105 VSS 0.00285f
C20530 VDD99.n459 VSS 0.00285f
C20531 VDD99.n460 VSS 0.00622f
C20532 VDD99.t16 VSS 0.0835f
C20533 VDD99.t104 VSS 0.102f
C20534 VDD99.t162 VSS 0.0474f
C20535 VDD99.n461 VSS 0.043f
C20536 VDD99.t21 VSS 0.00693f
C20537 VDD99.t20 VSS 0.0474f
C20538 VDD99.t160 VSS 0.0611f
C20539 VDD99.n462 VSS 0.0606f
C20540 VDD99.n463 VSS 0.0572f
C20541 VDD99.t161 VSS 0.0069f
C20542 VDD99.n464 VSS 0.0351f
C20543 VDD99.t39 VSS 0.0069f
C20544 VDD99.n465 VSS 0.00692f
C20545 VDD99.t38 VSS 0.0662f
C20546 VDD99.n466 VSS 0.0629f
C20547 VDD99.t428 VSS 0.0542f
C20548 VDD99.t266 VSS 0.0833f
C20549 VDD99.n467 VSS 0.043f
C20550 VDD99.t207 VSS 0.0069f
C20551 VDD99.n468 VSS 0.0226f
C20552 VDD99.n469 VSS 0.0741f
C20553 VDD99.t74 VSS 0.0165f
C20554 VDD99.t12 VSS 0.0069f
C20555 VDD99.t446 VSS 0.00285f
C20556 VDD99.n470 VSS 0.00285f
C20557 VDD99.n471 VSS 0.00622f
C20558 VDD99.n472 VSS 0.00692f
C20559 VDD99.n473 VSS 0.0519f
C20560 VDD99.t19 VSS 0.0069f
C20561 VDD99.t418 VSS 0.167f
C20562 VDD99.t420 VSS 0.00693f
C20563 VDD99.t419 VSS 0.00693f
C20564 VDD99.n474 VSS 0.0638f
C20565 VDD99.n475 VSS 0.0292f
C20566 VDD99.n476 VSS 0.086f
C20567 VDD99.t268 VSS 0.0947f
C20568 VDD99.t445 VSS 0.131f
C20569 VDD99.t73 VSS 0.0222f
C20570 VDD99.t18 VSS 0.0921f
C20571 VDD99.t206 VSS 0.0614f
C20572 VDD99.n478 VSS 0.0727f
C20573 VDD99.t205 VSS 0.0579f
C20574 VDD99.n479 VSS 0.0248f
C20575 VDD99.n480 VSS 0.0871f
C20576 VDD99.n481 VSS 0.0515f
C20577 VDD99.n482 VSS 0.0245f
C20578 VDD99.n483 VSS 0.0132f
C20579 VDD99.n484 VSS 0.072f
C20580 VDD99.t11 VSS 0.0849f
C20581 VDD99.n485 VSS 0.059f
C20582 VDD99.n486 VSS 0.0311f
C20583 VDD99.n487 VSS 0.0345f
C20584 VDD99.n488 VSS 0.0266f
C20585 VDD99.t267 VSS 0.00704f
C20586 VDD99.n489 VSS 0.0385f
C20587 VDD99.n490 VSS 0.0242f
C20588 VDD99.n491 VSS 0.034f
C20589 VDD99.n492 VSS 0.0319f
C20590 VDD99.n493 VSS 0.0285f
C20591 VDD99.n494 VSS 0.0355f
C20592 VDD99.n495 VSS 0.0225f
C20593 VDD99.n496 VSS 0.0311f
C20594 VDD99.n497 VSS 0.0328f
C20595 VDD99.n498 VSS 0.0253f
C20596 VDD99.n499 VSS 0.0375f
C20597 VDD99.n500 VSS 0.0347f
C20598 VDD99.n501 VSS 0.0253f
C20599 VDD99.n502 VSS 0.0375f
C20600 VDD99.n503 VSS 0.0347f
C20601 VDD99.n504 VSS 0.0253f
C20602 VDD99.n505 VSS 0.0367f
C20603 VDD99.n506 VSS 0.0616f
C20604 VDD99.n507 VSS 0.0385f
C20605 VDD99.n508 VSS 0.0404f
C20606 VDD99.n509 VSS 0.0226f
C20607 VDD99.n510 VSS 0.106f
C20608 VDD99.n511 VSS 1.3f
C20609 VDD99.n512 VSS 0.649f
C20610 VDD99.n513 VSS 0.613f
C20611 VDD99.n514 VSS 0.995f
C20612 VDD99.n515 VSS 0.00693f
C20613 VDD99.n516 VSS 0.00191f
C20614 VDD99.n517 VSS 0.0128f
C20615 VDD99.n518 VSS 2.67f
C20616 VDD99.n519 VSS 1.4f
C20617 VDD99.n520 VSS 1.4f
C20618 VDD99.n521 VSS 0.0721f
C20619 VDD99.n522 VSS 0.0975f
C20620 VDD99.n523 VSS 0.069f
C20621 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.t2 VSS 0.025f
C20622 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.t0 VSS 0.0206f
C20623 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.n0 VSS 0.0206f
C20624 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.n1 VSS 0.0494f
C20625 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.t8 VSS 0.0459f
C20626 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.t6 VSS 0.0302f
C20627 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.n2 VSS 0.0814f
C20628 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.t5 VSS 0.0329f
C20629 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.t7 VSS 0.0263f
C20630 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.n3 VSS 0.0764f
C20631 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.n4 VSS 0.606f
C20632 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.t4 VSS 0.0641f
C20633 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.t3 VSS 0.0199f
C20634 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.n5 VSS 0.0675f
C20635 CLK_div_90_mag_0.CLK_div_3_mag_0.Q0.n6 VSS 0.447f
C20636 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n0 VSS 0.651f
C20637 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n1 VSS 0.242f
C20638 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t9 VSS 0.0256f
C20639 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t6 VSS 0.0388f
C20640 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n2 VSS 0.0689f
C20641 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t14 VSS 0.0223f
C20642 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t12 VSS 0.0279f
C20643 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n3 VSS 0.0646f
C20644 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n4 VSS 0.499f
C20645 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t13 VSS 0.0223f
C20646 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t10 VSS 0.0279f
C20647 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n5 VSS 0.0726f
C20648 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t11 VSS 0.0223f
C20649 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t4 VSS 0.0279f
C20650 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n6 VSS 0.0661f
C20651 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n7 VSS 0.67f
C20652 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t3 VSS 0.0256f
C20653 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t15 VSS 0.0388f
C20654 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n8 VSS 0.0686f
C20655 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t7 VSS 0.0256f
C20656 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t5 VSS 0.0388f
C20657 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n9 VSS 0.0686f
C20658 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n10 VSS 0.276f
C20659 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t8 VSS 0.0321f
C20660 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.t2 VSS 0.0082f
C20661 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n11 VSS 0.0531f
C20662 CLK_div_93_mag_0.CLK_div_31_mag_0.Q3.n12 VSS 0.204f
C20663 VDD93.n0 VSS 0.0182f
C20664 VDD93.t247 VSS 0.0147f
C20665 VDD93.t249 VSS 0.00615f
C20666 VDD93.n1 VSS 0.0194f
C20667 VDD93.t248 VSS 0.0556f
C20668 VDD93.n2 VSS 0.286f
C20669 VDD93.n3 VSS 0.00616f
C20670 VDD93.t115 VSS 0.0487f
C20671 VDD93.t213 VSS 0.0743f
C20672 VDD93.n4 VSS 0.0384f
C20673 VDD93.t214 VSS 0.00616f
C20674 VDD93.n5 VSS 0.0168f
C20675 VDD93.t243 VSS 0.00254f
C20676 VDD93.n6 VSS 0.00254f
C20677 VDD93.n7 VSS 0.00555f
C20678 VDD93.t340 VSS 0.00618f
C20679 VDD93.n8 VSS 0.00618f
C20680 VDD93.n9 VSS 0.0306f
C20681 VDD93.t223 VSS 0.0816f
C20682 VDD93.n10 VSS 0.00618f
C20683 VDD93.t188 VSS 0.00618f
C20684 VDD93.n11 VSS 0.00618f
C20685 VDD93.n12 VSS 0.00618f
C20686 VDD93.t374 VSS 0.0805f
C20687 VDD93.n13 VSS 0.0384f
C20688 VDD93.t378 VSS 0.00618f
C20689 VDD93.n14 VSS 0.00618f
C20690 VDD93.t377 VSS 0.0745f
C20691 VDD93.t220 VSS 0.0816f
C20692 VDD93.n15 VSS 0.0384f
C20693 VDD93.t55 VSS 0.00618f
C20694 VDD93.t50 VSS 0.00254f
C20695 VDD93.n16 VSS 0.00254f
C20696 VDD93.n17 VSS 0.00555f
C20697 VDD93.t54 VSS 0.0745f
C20698 VDD93.t49 VSS 0.091f
C20699 VDD93.t403 VSS 0.0423f
C20700 VDD93.n18 VSS 0.0384f
C20701 VDD93.t312 VSS 0.00618f
C20702 VDD93.t372 VSS 0.00254f
C20703 VDD93.n19 VSS 0.00254f
C20704 VDD93.n20 VSS 0.00555f
C20705 VDD93.t311 VSS 0.0745f
C20706 VDD93.t371 VSS 0.091f
C20707 VDD93.t207 VSS 0.0423f
C20708 VDD93.t101 VSS 0.0743f
C20709 VDD93.n21 VSS 0.0384f
C20710 VDD93.t102 VSS 0.00663f
C20711 VDD93.n22 VSS 0.0476f
C20712 VDD93.n23 VSS 0.0352f
C20713 VDD93.n24 VSS 0.0361f
C20714 VDD93.n25 VSS 0.0192f
C20715 VDD93.n26 VSS 0.0352f
C20716 VDD93.n27 VSS 0.036f
C20717 VDD93.n28 VSS 0.0214f
C20718 VDD93.n29 VSS 0.0306f
C20719 VDD93.n30 VSS 0.0285f
C20720 VDD93.n31 VSS 0.0214f
C20721 VDD93.n32 VSS 0.0583f
C20722 VDD93.n33 VSS 0.0663f
C20723 VDD93.t239 VSS 0.0805f
C20724 VDD93.t187 VSS 0.0745f
C20725 VDD93.n34 VSS 0.0384f
C20726 VDD93.n35 VSS 0.0214f
C20727 VDD93.n36 VSS 0.0285f
C20728 VDD93.n37 VSS 0.0306f
C20729 VDD93.t48 VSS 0.00618f
C20730 VDD93.n38 VSS 0.0285f
C20731 VDD93.n39 VSS 0.0214f
C20732 VDD93.n40 VSS 0.0384f
C20733 VDD93.t47 VSS 0.0745f
C20734 VDD93.t51 VSS 0.0816f
C20735 VDD93.n41 VSS 0.0137f
C20736 VDD93.t111 VSS 0.00615f
C20737 VDD93.n42 VSS 0.0408f
C20738 VDD93.t216 VSS 0.00615f
C20739 VDD93.n43 VSS 0.315f
C20740 VDD93.n44 VSS 0.00618f
C20741 VDD93.t112 VSS 0.0805f
C20742 VDD93.n45 VSS 0.0384f
C20743 VDD93.t130 VSS 0.00618f
C20744 VDD93.n46 VSS 0.00618f
C20745 VDD93.t129 VSS 0.0745f
C20746 VDD93.t411 VSS 0.0816f
C20747 VDD93.n47 VSS 0.0384f
C20748 VDD93.t57 VSS 0.00618f
C20749 VDD93.t297 VSS 0.00254f
C20750 VDD93.n48 VSS 0.00254f
C20751 VDD93.n49 VSS 0.00555f
C20752 VDD93.t56 VSS 0.0745f
C20753 VDD93.t296 VSS 0.091f
C20754 VDD93.t394 VSS 0.0423f
C20755 VDD93.n50 VSS 0.0384f
C20756 VDD93.t121 VSS 0.00618f
C20757 VDD93.t119 VSS 0.00254f
C20758 VDD93.n51 VSS 0.00254f
C20759 VDD93.n52 VSS 0.00555f
C20760 VDD93.t120 VSS 0.0745f
C20761 VDD93.t118 VSS 0.091f
C20762 VDD93.t217 VSS 0.0423f
C20763 VDD93.t88 VSS 0.0743f
C20764 VDD93.n53 VSS 0.0384f
C20765 VDD93.t89 VSS 0.00577f
C20766 VDD93.t100 VSS 0.0053f
C20767 VDD93.t487 VSS 0.00402f
C20768 VDD93.n54 VSS 0.0104f
C20769 VDD93.n55 VSS 0.0581f
C20770 VDD93.n56 VSS 0.0759f
C20771 VDD93.n57 VSS 0.00136f
C20772 VDD93.t486 VSS 0.00401f
C20773 VDD93.n58 VSS 0.00543f
C20774 VDD93.t87 VSS 0.00515f
C20775 VDD93.n59 VSS 0.00508f
C20776 VDD93.n60 VSS 5.13e-20
C20777 VDD93.n61 VSS 0.0016f
C20778 VDD93.n62 VSS 7.36e-19
C20779 VDD93.n63 VSS 6.11e-19
C20780 VDD93.n64 VSS 0.0046f
C20781 VDD93.n65 VSS 0.0144f
C20782 VDD93.n66 VSS 0.0353f
C20783 VDD93.n67 VSS 0.0352f
C20784 VDD93.n68 VSS 0.0361f
C20785 VDD93.n69 VSS 0.0192f
C20786 VDD93.n70 VSS 0.0352f
C20787 VDD93.n71 VSS 0.036f
C20788 VDD93.n72 VSS 0.0214f
C20789 VDD93.n73 VSS 0.0306f
C20790 VDD93.n74 VSS 0.0285f
C20791 VDD93.n75 VSS 0.0214f
C20792 VDD93.n76 VSS 0.0533f
C20793 VDD93.n77 VSS 0.00614f
C20794 VDD93.t172 VSS 0.0649f
C20795 VDD93.t417 VSS 0.0593f
C20796 VDD93.n78 VSS 0.0331f
C20797 VDD93.t418 VSS 0.00615f
C20798 VDD93.n79 VSS 0.299f
C20799 VDD93.n80 VSS 0.00614f
C20800 VDD93.t414 VSS 0.0649f
C20801 VDD93.t298 VSS 0.0439f
C20802 VDD93.n81 VSS 0.0331f
C20803 VDD93.t299 VSS 0.00615f
C20804 VDD93.n82 VSS 0.00614f
C20805 VDD93.n83 VSS 0.309f
C20806 VDD93.n84 VSS 0.17f
C20807 VDD93.t58 VSS 0.0285f
C20808 VDD93.t24 VSS 0.0593f
C20809 VDD93.n85 VSS 0.0331f
C20810 VDD93.t25 VSS 0.00615f
C20811 VDD93.t171 VSS 0.00254f
C20812 VDD93.n86 VSS 0.00254f
C20813 VDD93.n87 VSS 0.00551f
C20814 VDD93.t170 VSS 0.0724f
C20815 VDD93.t210 VSS 0.0336f
C20816 VDD93.n88 VSS 0.0331f
C20817 VDD93.n89 VSS 0.0352f
C20818 VDD93.t434 VSS 0.00618f
C20819 VDD93.n90 VSS 0.0383f
C20820 VDD93.t141 VSS 0.0487f
C20821 VDD93.n91 VSS 0.00618f
C20822 VDD93.t436 VSS 0.00615f
C20823 VDD93.t461 VSS 0.0487f
C20824 VDD93.n92 VSS 0.00618f
C20825 VDD93.t182 VSS 0.00615f
C20826 VDD93.t360 VSS 0.0582f
C20827 VDD93.n93 VSS 0.0654f
C20828 VDD93.t361 VSS 0.00615f
C20829 VDD93.t358 VSS 0.0573f
C20830 VDD93.n94 VSS 0.066f
C20831 VDD93.t359 VSS 0.00615f
C20832 VDD93.n95 VSS 0.00618f
C20833 VDD93.t427 VSS 0.0813f
C20834 VDD93.n96 VSS 0.0384f
C20835 VDD93.t328 VSS 0.00618f
C20836 VDD93.t327 VSS 0.0725f
C20837 VDD93.t68 VSS 0.0544f
C20838 VDD93.n97 VSS 0.0593f
C20839 VDD93.t69 VSS 0.00615f
C20840 VDD93.n98 VSS 0.00618f
C20841 VDD93.t446 VSS 0.0487f
C20842 VDD93.n99 VSS 0.0384f
C20843 VDD93.t128 VSS 0.00623f
C20844 VDD93.t330 VSS 0.00619f
C20845 VDD93.n100 VSS 0.0441f
C20846 VDD93.t438 VSS 0.00618f
C20847 VDD93.t65 VSS 0.0805f
C20848 VDD93.n101 VSS 0.0225f
C20849 VDD93.n102 VSS 0.0418f
C20850 VDD93.t64 VSS 0.00254f
C20851 VDD93.n103 VSS 0.00254f
C20852 VDD93.n104 VSS 0.00555f
C20853 VDD93.t274 VSS 0.00618f
C20854 VDD93.t190 VSS 0.00618f
C20855 VDD93.n105 VSS 0.00618f
C20856 VDD93.n106 VSS 0.0316f
C20857 VDD93.n107 VSS 0.0392f
C20858 VDD93.t127 VSS 0.0738f
C20859 VDD93.t329 VSS 0.0526f
C20860 VDD93.n108 VSS 0.0571f
C20861 VDD93.t144 VSS 0.0487f
C20862 VDD93.n109 VSS 0.00618f
C20863 VDD93.n110 VSS 0.00618f
C20864 VDD93.n111 VSS 0.0402f
C20865 VDD93.n112 VSS 0.0394f
C20866 VDD93.n113 VSS 0.0319f
C20867 VDD93.n114 VSS 0.0384f
C20868 VDD93.t45 VSS 0.074f
C20869 VDD93.t43 VSS 0.0519f
C20870 VDD93.t44 VSS 0.0089f
C20871 VDD93.t310 VSS 0.00618f
C20872 VDD93.t46 VSS 0.00618f
C20873 VDD93.n115 VSS 0.032f
C20874 VDD93.n116 VSS 0.0564f
C20875 VDD93.n117 VSS 0.0119f
C20876 VDD93.n118 VSS 0.00618f
C20877 VDD93.n119 VSS 0.0405f
C20878 VDD93.n120 VSS 0.0567f
C20879 VDD93.t34 VSS 0.0487f
C20880 VDD93.t273 VSS 0.0743f
C20881 VDD93.n121 VSS 0.0384f
C20882 VDD93.n122 VSS 0.0411f
C20883 VDD93.n123 VSS 0.0405f
C20884 VDD93.n124 VSS 0.0454f
C20885 VDD93.n125 VSS 0.0279f
C20886 VDD93.t75 VSS 0.00618f
C20887 VDD93.n126 VSS 0.0616f
C20888 VDD93.t443 VSS 0.00615f
C20889 VDD93.n127 VSS 0.00618f
C20890 VDD93.t288 VSS 0.0805f
C20891 VDD93.n128 VSS 0.0384f
C20892 VDD93.t251 VSS 0.00618f
C20893 VDD93.n129 VSS 0.00618f
C20894 VDD93.t250 VSS 0.0745f
C20895 VDD93.t154 VSS 0.0816f
C20896 VDD93.n130 VSS 0.0384f
C20897 VDD93.t370 VSS 0.00618f
C20898 VDD93.t365 VSS 0.00254f
C20899 VDD93.n131 VSS 0.00254f
C20900 VDD93.n132 VSS 0.00555f
C20901 VDD93.t369 VSS 0.0745f
C20902 VDD93.t364 VSS 0.091f
C20903 VDD93.t397 VSS 0.0423f
C20904 VDD93.n133 VSS 0.0384f
C20905 VDD93.t314 VSS 0.00618f
C20906 VDD93.t445 VSS 0.00254f
C20907 VDD93.n134 VSS 0.00254f
C20908 VDD93.n135 VSS 0.00555f
C20909 VDD93.t313 VSS 0.0745f
C20910 VDD93.t444 VSS 0.091f
C20911 VDD93.t138 VSS 0.0423f
C20912 VDD93.t98 VSS 0.0743f
C20913 VDD93.n136 VSS 0.0384f
C20914 VDD93.t99 VSS 0.00618f
C20915 VDD93.t80 VSS 0.0053f
C20916 VDD93.t481 VSS 0.00402f
C20917 VDD93.n137 VSS 0.0104f
C20918 VDD93.n138 VSS 0.00975f
C20919 VDD93.t97 VSS 0.0053f
C20920 VDD93.t475 VSS 0.00402f
C20921 VDD93.n139 VSS 0.0104f
C20922 VDD93.n140 VSS 0.00783f
C20923 VDD93.n141 VSS 0.0408f
C20924 VDD93.n142 VSS 0.0288f
C20925 VDD93.n143 VSS 0.0192f
C20926 VDD93.n144 VSS 0.0352f
C20927 VDD93.n145 VSS 0.0361f
C20928 VDD93.n146 VSS 0.0192f
C20929 VDD93.n147 VSS 0.0352f
C20930 VDD93.n148 VSS 0.036f
C20931 VDD93.n149 VSS 0.0214f
C20932 VDD93.n150 VSS 0.0306f
C20933 VDD93.n151 VSS 0.0285f
C20934 VDD93.n152 VSS 0.0214f
C20935 VDD93.n153 VSS 0.055f
C20936 VDD93.t466 VSS 0.0547f
C20937 VDD93.n154 VSS 0.0574f
C20938 VDD93.n155 VSS 0.00776f
C20939 VDD93.n156 VSS 0.00618f
C20940 VDD93.t10 VSS 0.0805f
C20941 VDD93.n157 VSS 0.0384f
C20942 VDD93.n158 VSS 0.00618f
C20943 VDD93.t17 VSS 0.00618f
C20944 VDD93.t84 VSS 0.0424f
C20945 VDD93.n159 VSS 0.0384f
C20946 VDD93.n160 VSS 0.00618f
C20947 VDD93.t470 VSS 0.00254f
C20948 VDD93.n161 VSS 0.00254f
C20949 VDD93.n162 VSS 0.00555f
C20950 VDD93.t16 VSS 0.0745f
C20951 VDD93.t157 VSS 0.0816f
C20952 VDD93.n163 VSS 0.0384f
C20953 VDD93.t363 VSS 0.00618f
C20954 VDD93.n164 VSS 0.00618f
C20955 VDD93.n165 VSS 0.00618f
C20956 VDD93.t469 VSS 0.0421f
C20957 VDD93.t324 VSS 0.091f
C20958 VDD93.t331 VSS 0.0747f
C20959 VDD93.n166 VSS 0.0384f
C20960 VDD93.t362 VSS 0.0745f
C20961 VDD93.t366 VSS 0.0816f
C20962 VDD93.n167 VSS 0.0384f
C20963 VDD93.t123 VSS 0.00618f
C20964 VDD93.t316 VSS 0.00618f
C20965 VDD93.n168 VSS 0.00618f
C20966 VDD93.t122 VSS 0.0815f
C20967 VDD93.t352 VSS 0.0747f
C20968 VDD93.n169 VSS 0.0384f
C20969 VDD93.t9 VSS 0.00254f
C20970 VDD93.n170 VSS 0.00254f
C20971 VDD93.n171 VSS 0.00555f
C20972 VDD93.t346 VSS 0.00618f
C20973 VDD93.t315 VSS 0.0745f
C20974 VDD93.t8 VSS 0.091f
C20975 VDD93.t151 VSS 0.0423f
C20976 VDD93.n172 VSS 0.0384f
C20977 VDD93.n173 VSS 0.00618f
C20978 VDD93.t82 VSS 0.00618f
C20979 VDD93.t345 VSS 0.0815f
C20980 VDD93.t355 VSS 0.0747f
C20981 VDD93.t322 VSS 0.0803f
C20982 VDD93.n174 VSS 0.0384f
C20983 VDD93.t323 VSS 0.00618f
C20984 VDD93.t148 VSS 0.00777f
C20985 VDD93.t147 VSS 0.0545f
C20986 VDD93.t81 VSS 0.0423f
C20987 VDD93.n175 VSS 0.0574f
C20988 VDD93.n176 VSS 0.00618f
C20989 VDD93.t135 VSS 0.0805f
C20990 VDD93.n177 VSS 0.0384f
C20991 VDD93.t227 VSS 0.00618f
C20992 VDD93.n178 VSS 0.00618f
C20993 VDD93.t226 VSS 0.0745f
C20994 VDD93.t194 VSS 0.0816f
C20995 VDD93.n179 VSS 0.0384f
C20996 VDD93.t169 VSS 0.00618f
C20997 VDD93.t229 VSS 0.00254f
C20998 VDD93.n180 VSS 0.00254f
C20999 VDD93.n181 VSS 0.00555f
C21000 VDD93.t168 VSS 0.0745f
C21001 VDD93.t228 VSS 0.091f
C21002 VDD93.t406 VSS 0.0423f
C21003 VDD93.n182 VSS 0.0384f
C21004 VDD93.t62 VSS 0.00618f
C21005 VDD93.t150 VSS 0.00254f
C21006 VDD93.n183 VSS 0.00254f
C21007 VDD93.n184 VSS 0.00555f
C21008 VDD93.t61 VSS 0.0745f
C21009 VDD93.t149 VSS 0.091f
C21010 VDD93.t455 VSS 0.0423f
C21011 VDD93.t71 VSS 0.0743f
C21012 VDD93.n185 VSS 0.0384f
C21013 VDD93.t72 VSS 0.00618f
C21014 VDD93.t94 VSS 0.0053f
C21015 VDD93.t477 VSS 0.00402f
C21016 VDD93.n186 VSS 0.0104f
C21017 VDD93.n187 VSS 0.00861f
C21018 VDD93.t70 VSS 0.0053f
C21019 VDD93.t485 VSS 0.00402f
C21020 VDD93.n188 VSS 0.0104f
C21021 VDD93.n189 VSS 0.00828f
C21022 VDD93.n190 VSS 0.0424f
C21023 VDD93.n191 VSS 0.0288f
C21024 VDD93.n192 VSS 0.0192f
C21025 VDD93.n193 VSS 0.0352f
C21026 VDD93.n194 VSS 0.0361f
C21027 VDD93.n195 VSS 0.0192f
C21028 VDD93.n196 VSS 0.0352f
C21029 VDD93.n197 VSS 0.036f
C21030 VDD93.n198 VSS 0.0214f
C21031 VDD93.n199 VSS 0.0306f
C21032 VDD93.n200 VSS 0.0285f
C21033 VDD93.n201 VSS 0.0214f
C21034 VDD93.n202 VSS 0.0558f
C21035 VDD93.t279 VSS 0.0547f
C21036 VDD93.n203 VSS 0.0574f
C21037 VDD93.n204 VSS 0.00776f
C21038 VDD93.n205 VSS 0.00618f
C21039 VDD93.t160 VSS 0.0649f
C21040 VDD93.n206 VSS 0.0331f
C21041 VDD93.n207 VSS 0.00618f
C21042 VDD93.t233 VSS 0.00618f
C21043 VDD93.t91 VSS 0.0424f
C21044 VDD93.n208 VSS 0.0384f
C21045 VDD93.n209 VSS 0.00618f
C21046 VDD93.t270 VSS 0.00254f
C21047 VDD93.n210 VSS 0.00254f
C21048 VDD93.n211 VSS 0.00555f
C21049 VDD93.t232 VSS 0.0593f
C21050 VDD93.t197 VSS 0.0649f
C21051 VDD93.n212 VSS 0.0331f
C21052 VDD93.t231 VSS 0.00618f
C21053 VDD93.n213 VSS 0.00618f
C21054 VDD93.n214 VSS 0.00618f
C21055 VDD93.t269 VSS 0.0421f
C21056 VDD93.t236 VSS 0.091f
C21057 VDD93.t382 VSS 0.0747f
C21058 VDD93.n215 VSS 0.0384f
C21059 VDD93.n216 VSS 0.0331f
C21060 VDD93.t266 VSS 0.00618f
C21061 VDD93.t342 VSS 0.00618f
C21062 VDD93.n217 VSS 0.00618f
C21063 VDD93.t265 VSS 0.0815f
C21064 VDD93.t259 VSS 0.0747f
C21065 VDD93.n218 VSS 0.0384f
C21066 VDD93.t164 VSS 0.00254f
C21067 VDD93.n219 VSS 0.00254f
C21068 VDD93.n220 VSS 0.00555f
C21069 VDD93.t386 VSS 0.00618f
C21070 VDD93.t341 VSS 0.0593f
C21071 VDD93.t163 VSS 0.0724f
C21072 VDD93.t302 VSS 0.0336f
C21073 VDD93.n221 VSS 0.0331f
C21074 VDD93.n222 VSS 0.00618f
C21075 VDD93.t96 VSS 0.00618f
C21076 VDD93.t385 VSS 0.0815f
C21077 VDD93.t291 VSS 0.0747f
C21078 VDD93.t234 VSS 0.0803f
C21079 VDD93.n223 VSS 0.0384f
C21080 VDD93.t235 VSS 0.00618f
C21081 VDD93.t301 VSS 0.00777f
C21082 VDD93.t95 VSS 0.0336f
C21083 VDD93.t230 VSS 0.0439f
C21084 VDD93.t165 VSS 0.0285f
C21085 VDD93.n224 VSS 0.171f
C21086 VDD93.n225 VSS 0.0947f
C21087 VDD93.t300 VSS 0.0681f
C21088 VDD93.t306 VSS 0.00618f
C21089 VDD93.t262 VSS 0.0747f
C21090 VDD93.n226 VSS 0.00618f
C21091 VDD93.t410 VSS 0.00254f
C21092 VDD93.n227 VSS 0.00254f
C21093 VDD93.n228 VSS 0.00555f
C21094 VDD93.n229 VSS 0.00618f
C21095 VDD93.n230 VSS 0.0361f
C21096 VDD93.t77 VSS 0.0745f
C21097 VDD93.n231 VSS 0.00618f
C21098 VDD93.t480 VSS 0.00402f
C21099 VDD93.t76 VSS 0.0053f
C21100 VDD93.n232 VSS 0.0104f
C21101 VDD93.t476 VSS 0.00402f
C21102 VDD93.t90 VSS 0.0053f
C21103 VDD93.n233 VSS 0.0104f
C21104 VDD93.n234 VSS 0.00158f
C21105 VDD93.n235 VSS 0.00938f
C21106 VDD93.n236 VSS 0.0512f
C21107 VDD93.n237 VSS 0.0288f
C21108 VDD93.t276 VSS 0.00254f
C21109 VDD93.n238 VSS 0.00254f
C21110 VDD93.n239 VSS 0.00555f
C21111 VDD93.n240 VSS 0.0353f
C21112 VDD93.n241 VSS 0.0191f
C21113 VDD93.n242 VSS 0.0384f
C21114 VDD93.t275 VSS 0.0421f
C21115 VDD93.t458 VSS 0.091f
C21116 VDD93.t18 VSS 0.0747f
C21117 VDD93.t256 VSS 0.091f
C21118 VDD93.t409 VSS 0.0421f
C21119 VDD93.n243 VSS 0.0384f
C21120 VDD93.n244 VSS 0.0191f
C21121 VDD93.n245 VSS 0.0353f
C21122 VDD93.n246 VSS 0.036f
C21123 VDD93.t388 VSS 0.00618f
C21124 VDD93.n247 VSS 0.00618f
C21125 VDD93.n248 VSS 0.0284f
C21126 VDD93.n249 VSS 0.0306f
C21127 VDD93.n250 VSS 0.0214f
C21128 VDD93.n251 VSS 0.0384f
C21129 VDD93.t387 VSS 0.0815f
C21130 VDD93.t389 VSS 0.0747f
C21131 VDD93.t305 VSS 0.0803f
C21132 VDD93.n252 VSS 0.0384f
C21133 VDD93.n253 VSS 0.0214f
C21134 VDD93.n254 VSS 0.0577f
C21135 VDD93.n255 VSS 0.0139f
C21136 VDD93.n256 VSS 0.0368f
C21137 VDD93.n257 VSS 0.038f
C21138 VDD93.n258 VSS 0.0289f
C21139 VDD93.n259 VSS 0.0293f
C21140 VDD93.n260 VSS 0.0305f
C21141 VDD93.n261 VSS 0.0352f
C21142 VDD93.n262 VSS 0.0326f
C21143 VDD93.n263 VSS 0.0282f
C21144 VDD93.n264 VSS 0.0391f
C21145 VDD93.n265 VSS 0.0435f
C21146 VDD93.n266 VSS 0.0289f
C21147 VDD93.n267 VSS 0.0313f
C21148 VDD93.n268 VSS 0.0314f
C21149 VDD93.n269 VSS 0.0288f
C21150 VDD93.n270 VSS 0.0435f
C21151 VDD93.n271 VSS 0.0393f
C21152 VDD93.n272 VSS 0.028f
C21153 VDD93.n273 VSS 0.0326f
C21154 VDD93.n274 VSS 0.0353f
C21155 VDD93.n275 VSS 0.0304f
C21156 VDD93.n276 VSS 0.0293f
C21157 VDD93.n277 VSS 0.0291f
C21158 VDD93.n278 VSS 0.0378f
C21159 VDD93.n279 VSS 0.037f
C21160 VDD93.n280 VSS 0.0141f
C21161 VDD93.n281 VSS 0.0667f
C21162 VDD93.t272 VSS 0.00618f
C21163 VDD93.t124 VSS 0.0747f
C21164 VDD93.n282 VSS 0.00618f
C21165 VDD93.t393 VSS 0.00254f
C21166 VDD93.n283 VSS 0.00254f
C21167 VDD93.n284 VSS 0.00555f
C21168 VDD93.n285 VSS 0.00618f
C21169 VDD93.n286 VSS 0.0361f
C21170 VDD93.t107 VSS 0.0745f
C21171 VDD93.n287 VSS 0.00618f
C21172 VDD93.t483 VSS 0.00402f
C21173 VDD93.t106 VSS 0.0053f
C21174 VDD93.n288 VSS 0.0104f
C21175 VDD93.n289 VSS 0.0029f
C21176 VDD93.t478 VSS 0.00402f
C21177 VDD93.t83 VSS 0.0053f
C21178 VDD93.n290 VSS 0.0104f
C21179 VDD93.n291 VSS 0.00847f
C21180 VDD93.n292 VSS 0.0462f
C21181 VDD93.n293 VSS 0.0288f
C21182 VDD93.t465 VSS 0.00254f
C21183 VDD93.n294 VSS 0.00254f
C21184 VDD93.n295 VSS 0.00555f
C21185 VDD93.n296 VSS 0.0353f
C21186 VDD93.n297 VSS 0.0191f
C21187 VDD93.n298 VSS 0.0384f
C21188 VDD93.t464 VSS 0.0421f
C21189 VDD93.t282 VSS 0.091f
C21190 VDD93.t319 VSS 0.0747f
C21191 VDD93.t349 VSS 0.091f
C21192 VDD93.t392 VSS 0.0421f
C21193 VDD93.n299 VSS 0.0384f
C21194 VDD93.n300 VSS 0.0191f
C21195 VDD93.n301 VSS 0.0353f
C21196 VDD93.n302 VSS 0.036f
C21197 VDD93.t348 VSS 0.00618f
C21198 VDD93.n303 VSS 0.00618f
C21199 VDD93.n304 VSS 0.0284f
C21200 VDD93.n305 VSS 0.0306f
C21201 VDD93.n306 VSS 0.0214f
C21202 VDD93.n307 VSS 0.0384f
C21203 VDD93.t347 VSS 0.0815f
C21204 VDD93.t191 VSS 0.0747f
C21205 VDD93.t271 VSS 0.0803f
C21206 VDD93.n308 VSS 0.0384f
C21207 VDD93.n309 VSS 0.0214f
C21208 VDD93.n310 VSS 0.0549f
C21209 VDD93.n311 VSS 0.0636f
C21210 VDD93.n312 VSS 0.0163f
C21211 VDD93.n313 VSS 0.0386f
C21212 VDD93.n314 VSS 0.0374f
C21213 VDD93.n315 VSS 0.0285f
C21214 VDD93.n316 VSS 0.0289f
C21215 VDD93.n317 VSS 0.0277f
C21216 VDD93.n318 VSS 0.0346f
C21217 VDD93.n319 VSS 0.032f
C21218 VDD93.n320 VSS 0.0302f
C21219 VDD93.n321 VSS 0.0385f
C21220 VDD93.n322 VSS 0.0427f
C21221 VDD93.n323 VSS 0.0285f
C21222 VDD93.n324 VSS 0.0333f
C21223 VDD93.n325 VSS 0.0334f
C21224 VDD93.n326 VSS 0.0284f
C21225 VDD93.n327 VSS 0.0427f
C21226 VDD93.n328 VSS 0.0386f
C21227 VDD93.n329 VSS 0.0301f
C21228 VDD93.n330 VSS 0.032f
C21229 VDD93.n331 VSS 0.0348f
C21230 VDD93.n332 VSS 0.0276f
C21231 VDD93.n333 VSS 0.0289f
C21232 VDD93.n334 VSS 0.0286f
C21233 VDD93.n335 VSS 0.0373f
C21234 VDD93.n336 VSS 0.0388f
C21235 VDD93.n337 VSS 0.0164f
C21236 VDD93.n338 VSS 0.0655f
C21237 VDD93.n339 VSS 0.0595f
C21238 VDD93.t442 VSS 0.0545f
C21239 VDD93.n340 VSS 0.0574f
C21240 VDD93.t74 VSS 0.0423f
C21241 VDD93.n341 VSS 0.0384f
C21242 VDD93.t439 VSS 0.0423f
C21243 VDD93.t63 VSS 0.091f
C21244 VDD93.t189 VSS 0.0745f
C21245 VDD93.n342 VSS 0.0384f
C21246 VDD93.t334 VSS 0.0816f
C21247 VDD93.t309 VSS 0.0745f
C21248 VDD93.n343 VSS 0.0384f
C21249 VDD93.t422 VSS 0.0816f
C21250 VDD93.t437 VSS 0.0745f
C21251 VDD93.n344 VSS 0.0384f
C21252 VDD93.n345 VSS 0.0182f
C21253 VDD93.n346 VSS 0.017f
C21254 VDD93.n347 VSS 0.00588f
C21255 VDD93.n348 VSS 0.00902f
C21256 VDD93.t253 VSS 0.00616f
C21257 VDD93.n349 VSS 0.00616f
C21258 VDD93.n350 VSS 0.0339f
C21259 VDD93.t2 VSS 0.0847f
C21260 VDD93.n351 VSS 0.00616f
C21261 VDD93.t201 VSS 0.00616f
C21262 VDD93.n352 VSS 0.00616f
C21263 VDD93.n353 VSS 0.0337f
C21264 VDD93.t200 VSS 0.103f
C21265 VDD93.n354 VSS 0.0422f
C21266 VDD93.t21 VSS 0.103f
C21267 VDD93.n355 VSS 0.0882f
C21268 VDD93.n356 VSS 0.0886f
C21269 VDD93.n357 VSS 0.00616f
C21270 VDD93.t184 VSS 0.0112f
C21271 VDD93.n358 VSS 0.00753f
C21272 VDD93.t175 VSS 0.159f
C21273 VDD93.n359 VSS 0.00616f
C21274 VDD93.t186 VSS 0.0112f
C21275 VDD93.n360 VSS 0.00743f
C21276 VDD93.t13 VSS 0.159f
C21277 VDD93.n361 VSS 0.00616f
C21278 VDD93.t27 VSS 0.0112f
C21279 VDD93.n362 VSS 0.00743f
C21280 VDD93.t430 VSS 0.159f
C21281 VDD93.n363 VSS 0.00616f
C21282 VDD93.t380 VSS 0.0112f
C21283 VDD93.n364 VSS 0.00751f
C21284 VDD93.t40 VSS 0.129f
C21285 VDD93.n365 VSS 0.00651f
C21286 VDD93.n366 VSS 0.0308f
C21287 VDD93.n367 VSS 0.016f
C21288 VDD93.t379 VSS 0.159f
C21289 VDD93.n368 VSS 0.016f
C21290 VDD93.n369 VSS 0.0215f
C21291 VDD93.n370 VSS 0.0276f
C21292 VDD93.n371 VSS 0.016f
C21293 VDD93.t26 VSS 0.159f
C21294 VDD93.n372 VSS 0.016f
C21295 VDD93.n373 VSS 0.0215f
C21296 VDD93.n374 VSS 0.0276f
C21297 VDD93.n375 VSS 0.016f
C21298 VDD93.t185 VSS 0.159f
C21299 VDD93.n376 VSS 0.016f
C21300 VDD93.n377 VSS 0.0215f
C21301 VDD93.n378 VSS 0.0276f
C21302 VDD93.n379 VSS 0.016f
C21303 VDD93.t183 VSS 0.0756f
C21304 VDD93.n380 VSS 0.016f
C21305 VDD93.n381 VSS 0.0312f
C21306 VDD93.t178 VSS 0.102f
C21307 VDD93.n382 VSS 0.0559f
C21308 VDD93.t295 VSS 0.00616f
C21309 VDD93.n383 VSS 0.0379f
C21310 VDD93.t294 VSS 0.102f
C21311 VDD93.n384 VSS 0.0516f
C21312 VDD93.n385 VSS 0.0277f
C21313 VDD93.n386 VSS 0.0439f
C21314 VDD93.n387 VSS 0.0416f
C21315 VDD93.n388 VSS 0.034f
C21316 VDD93.n389 VSS 0.0324f
C21317 VDD93.t255 VSS 0.00616f
C21318 VDD93.n390 VSS 0.0324f
C21319 VDD93.n391 VSS 0.0335f
C21320 VDD93.t254 VSS 0.147f
C21321 VDD93.t5 VSS 0.141f
C21322 VDD93.t252 VSS 0.117f
C21323 VDD93.n392 VSS 0.0354f
C21324 VDD93.n393 VSS 0.0499f
C21325 VDD93.n394 VSS 0.00618f
C21326 VDD93.t37 VSS 0.0805f
C21327 VDD93.n395 VSS 0.0384f
C21328 VDD93.t132 VSS 0.00618f
C21329 VDD93.n396 VSS 0.00618f
C21330 VDD93.t131 VSS 0.0745f
C21331 VDD93.t419 VSS 0.0816f
C21332 VDD93.n397 VSS 0.0384f
C21333 VDD93.t338 VSS 0.00618f
C21334 VDD93.t308 VSS 0.00254f
C21335 VDD93.n398 VSS 0.00254f
C21336 VDD93.n399 VSS 0.00555f
C21337 VDD93.t337 VSS 0.0745f
C21338 VDD93.t307 VSS 0.091f
C21339 VDD93.t400 VSS 0.0423f
C21340 VDD93.n400 VSS 0.0384f
C21341 VDD93.t426 VSS 0.00618f
C21342 VDD93.t33 VSS 0.00254f
C21343 VDD93.n401 VSS 0.00254f
C21344 VDD93.n402 VSS 0.00555f
C21345 VDD93.t425 VSS 0.0745f
C21346 VDD93.t32 VSS 0.091f
C21347 VDD93.t452 VSS 0.0423f
C21348 VDD93.t104 VSS 0.0743f
C21349 VDD93.n403 VSS 0.0384f
C21350 VDD93.t105 VSS 0.00618f
C21351 VDD93.t73 VSS 0.0053f
C21352 VDD93.t484 VSS 0.00402f
C21353 VDD93.n404 VSS 0.0104f
C21354 VDD93.n405 VSS 0.00959f
C21355 VDD93.t103 VSS 0.0053f
C21356 VDD93.t474 VSS 0.00402f
C21357 VDD93.n406 VSS 0.0104f
C21358 VDD93.n407 VSS 0.00777f
C21359 VDD93.n408 VSS 0.0496f
C21360 VDD93.n409 VSS 0.0288f
C21361 VDD93.n410 VSS 0.0192f
C21362 VDD93.n411 VSS 0.0352f
C21363 VDD93.n412 VSS 0.0361f
C21364 VDD93.n413 VSS 0.0192f
C21365 VDD93.n414 VSS 0.0352f
C21366 VDD93.n415 VSS 0.036f
C21367 VDD93.n416 VSS 0.0214f
C21368 VDD93.n417 VSS 0.0306f
C21369 VDD93.n418 VSS 0.0285f
C21370 VDD93.n419 VSS 0.0214f
C21371 VDD93.n420 VSS 0.0227f
C21372 VDD93.n421 VSS 0.0505f
C21373 VDD93.n422 VSS 0.0463f
C21374 VDD93.n423 VSS 0.0595f
C21375 VDD93.n424 VSS 0.017f
C21376 VDD93.n425 VSS 0.0255f
C21377 VDD93.n426 VSS 0.0399f
C21378 VDD93.n427 VSS 0.0348f
C21379 VDD93.n428 VSS 0.041f
C21380 VDD93.n429 VSS 0.0253f
C21381 VDD93.n430 VSS 0.0385f
C21382 VDD93.n431 VSS 0.0337f
C21383 VDD93.n432 VSS 0.0349f
C21384 VDD93.t31 VSS 0.0148f
C21385 VDD93.t472 VSS 0.00615f
C21386 VDD93.n433 VSS 0.033f
C21387 VDD93.t471 VSS 0.0548f
C21388 VDD93.n434 VSS 0.0649f
C21389 VDD93.t381 VSS 0.0583f
C21390 VDD93.t30 VSS 0.0946f
C21391 VDD93.n435 VSS 0.0455f
C21392 VDD93.n436 VSS 0.0329f
C21393 VDD93.n437 VSS 0.0275f
C21394 VDD93.n438 VSS 0.108f
C21395 VDD93.n439 VSS 0.156f
C21396 VDD93.t181 VSS 0.0551f
C21397 VDD93.n440 VSS 0.057f
C21398 VDD93.n441 VSS 0.0337f
C21399 VDD93.n442 VSS 0.0385f
C21400 VDD93.t134 VSS 0.00618f
C21401 VDD93.n443 VSS 0.0402f
C21402 VDD93.n444 VSS 0.0253f
C21403 VDD93.n445 VSS 0.0384f
C21404 VDD93.t133 VSS 0.0726f
C21405 VDD93.t435 VSS 0.0543f
C21406 VDD93.n446 VSS 0.0593f
C21407 VDD93.n447 VSS 0.0348f
C21408 VDD93.n448 VSS 0.0399f
C21409 VDD93.n449 VSS 0.026f
C21410 VDD93.n450 VSS 0.0384f
C21411 VDD93.t433 VSS 0.0738f
C21412 VDD93.t267 VSS 0.0525f
C21413 VDD93.n451 VSS 0.0571f
C21414 VDD93.t268 VSS 0.00615f
C21415 VDD93.n452 VSS 0.00618f
C21416 VDD93.t285 VSS 0.0487f
C21417 VDD93.n453 VSS 0.0384f
C21418 VDD93.t344 VSS 0.00618f
C21419 VDD93.t343 VSS 0.074f
C21420 VDD93.t0 VSS 0.0518f
C21421 VDD93.n454 VSS 0.0567f
C21422 VDD93.t1 VSS 0.00615f
C21423 VDD93.n455 VSS 0.00618f
C21424 VDD93.t449 VSS 0.0487f
C21425 VDD93.t277 VSS 0.0743f
C21426 VDD93.n456 VSS 0.0384f
C21427 VDD93.t278 VSS 0.00655f
C21428 VDD93.n457 VSS 0.025f
C21429 VDD93.n458 VSS 0.0378f
C21430 VDD93.n459 VSS 0.0332f
C21431 VDD93.n460 VSS 0.0387f
C21432 VDD93.n461 VSS 0.0253f
C21433 VDD93.n462 VSS 0.0385f
C21434 VDD93.n463 VSS 0.0337f
C21435 VDD93.n464 VSS 0.033f
C21436 VDD93.n465 VSS 0.187f
C21437 VDD93.n466 VSS 0.236f
C21438 VDD93.n467 VSS 0.399f
C21439 VDD93.n468 VSS 0.00123f
C21440 VDD93.n469 VSS 0.00618f
C21441 VDD93.n470 VSS 0.0242f
C21442 VDD93.n471 VSS 0.432f
C21443 VDD93.n472 VSS 0.386f
C21444 VDD93.t245 VSS 0.00615f
C21445 VDD93.t244 VSS 0.0336f
C21446 VDD93.n473 VSS 0.0946f
C21447 VDD93.t205 VSS 0.0681f
C21448 VDD93.t206 VSS 0.00637f
C21449 VDD93.n474 VSS 0.04f
C21450 VDD93.n475 VSS 0.153f
C21451 VDD93.n476 VSS 0.0145f
C21452 VDD93.n477 VSS 0.0327f
C21453 VDD93.n478 VSS 0.0338f
C21454 VDD93.n479 VSS 0.0181f
C21455 VDD93.n480 VSS 0.157f
C21456 VDD93.n481 VSS 0.0338f
C21457 VDD93.n482 VSS 0.036f
C21458 VDD93.n483 VSS 0.0252f
C21459 VDD93.n484 VSS 0.0289f
C21460 VDD93.n485 VSS 0.162f
C21461 VDD93.n486 VSS 0.0297f
C21462 VDD93.n487 VSS 0.0252f
C21463 VDD93.n488 VSS 0.0382f
C21464 VDD93.n489 VSS 0.0427f
C21465 VDD93.n490 VSS 0.161f
C21466 VDD93.n491 VSS 0.0298f
C21467 VDD93.t215 VSS 0.0545f
C21468 VDD93.n492 VSS 0.0574f
C21469 VDD93.t110 VSS 0.0423f
C21470 VDD93.n493 VSS 0.0384f
C21471 VDD93.t202 VSS 0.0423f
C21472 VDD93.t242 VSS 0.091f
C21473 VDD93.t339 VSS 0.0745f
C21474 VDD93.n494 VSS 0.0384f
C21475 VDD93.n495 VSS 0.0214f
C21476 VDD93.n496 VSS 0.0269f
C21477 VDD93.n497 VSS 0.0234f
C21478 VDD93.n498 VSS 0.024f
C21479 VDD93.n499 VSS 0.0418f
C21480 VDD93.n500 VSS 0.0341f
C21481 VDD93.n501 VSS 0.141f
C21482 VDD93.n502 VSS 0.0235f
C21483 VDD93.n503 VSS 0.0231f
C21484 VDD93.n504 VSS 0.0301f
C21485 VDD93.n505 VSS 0.14f
C21486 VDD93.n506 VSS 0.872f
C21487 VDD93.n507 VSS 0.182f
C21488 VDD93.t318 VSS 0.00618f
C21489 VDD93.t317 VSS 0.0548f
C21490 VDD93.n508 VSS 0.0635f
C21491 VDD93.t373 VSS 0.0553f
C21492 VDD93.n509 VSS 0.0373f
C21493 VDD93.t246 VSS 0.0525f
C21494 VDD93.n510 VSS 0.0963f
C21495 VDD93.n511 VSS 0.0425f
C21496 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.t7 VSS 0.0156f
C21497 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.t3 VSS 0.0237f
C21498 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.n0 VSS 0.0421f
C21499 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.t2 VSS 0.0136f
C21500 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.t8 VSS 0.0171f
C21501 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.n1 VSS 0.0395f
C21502 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.n2 VSS 0.308f
C21503 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.t9 VSS 0.0389f
C21504 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.t5 VSS 0.00562f
C21505 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.n3 VSS 0.0323f
C21506 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.t6 VSS 0.0136f
C21507 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.t4 VSS 0.0171f
C21508 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.n4 VSS 0.0404f
C21509 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.n5 VSS 1.36f
C21510 CLK_div_93_mag_0.CLK_div_31_mag_0.Q4.n6 VSS 0.186f
C21511 VDD96.t49 VSS 0.0551f
C21512 VDD96.n0 VSS 0.0639f
C21513 VDD96.t50 VSS 0.00619f
C21514 VDD96.t313 VSS 0.0557f
C21515 VDD96.n1 VSS 0.0375f
C21516 VDD96.t257 VSS 0.0149f
C21517 VDD96.t256 VSS 0.0529f
C21518 VDD96.t34 VSS 0.056f
C21519 VDD96.n2 VSS 0.0969f
C21520 VDD96.t35 VSS 0.00619f
C21521 VDD96.n3 VSS 0.00621f
C21522 VDD96.t362 VSS 0.049f
C21523 VDD96.t71 VSS 0.0748f
C21524 VDD96.n4 VSS 0.0386f
C21525 VDD96.t72 VSS 0.00622f
C21526 VDD96.t361 VSS 0.00622f
C21527 VDD96.n5 VSS 0.0311f
C21528 VDD96.t330 VSS 0.00256f
C21529 VDD96.n6 VSS 0.00256f
C21530 VDD96.n7 VSS 0.00558f
C21531 VDD96.n8 VSS 0.0201f
C21532 VDD96.t133 VSS 0.0821f
C21533 VDD96.n9 VSS 0.00621f
C21534 VDD96.t273 VSS 0.00622f
C21535 VDD96.n10 VSS 0.00621f
C21536 VDD96.n11 VSS 0.0308f
C21537 VDD96.t333 VSS 0.081f
C21538 VDD96.n12 VSS 0.00621f
C21539 VDD96.n13 VSS 0.00621f
C21540 VDD96.t310 VSS 0.081f
C21541 VDD96.n14 VSS 0.0386f
C21542 VDD96.t197 VSS 0.00622f
C21543 VDD96.n15 VSS 0.00621f
C21544 VDD96.t196 VSS 0.075f
C21545 VDD96.t139 VSS 0.0821f
C21546 VDD96.n16 VSS 0.0386f
C21547 VDD96.t132 VSS 0.00622f
C21548 VDD96.t271 VSS 0.00256f
C21549 VDD96.n17 VSS 0.00256f
C21550 VDD96.n18 VSS 0.00558f
C21551 VDD96.t131 VSS 0.075f
C21552 VDD96.t270 VSS 0.0915f
C21553 VDD96.t294 VSS 0.0425f
C21554 VDD96.n19 VSS 0.0386f
C21555 VDD96.t199 VSS 0.00622f
C21556 VDD96.t309 VSS 0.00256f
C21557 VDD96.n20 VSS 0.00256f
C21558 VDD96.n21 VSS 0.00558f
C21559 VDD96.t198 VSS 0.075f
C21560 VDD96.t308 VSS 0.0915f
C21561 VDD96.t68 VSS 0.0425f
C21562 VDD96.t176 VSS 0.0748f
C21563 VDD96.n22 VSS 0.0386f
C21564 VDD96.t177 VSS 0.00667f
C21565 VDD96.n23 VSS 0.0479f
C21566 VDD96.n24 VSS 0.0354f
C21567 VDD96.n25 VSS 0.0364f
C21568 VDD96.n26 VSS 0.0193f
C21569 VDD96.n27 VSS 0.0354f
C21570 VDD96.n28 VSS 0.0363f
C21571 VDD96.n29 VSS 0.0215f
C21572 VDD96.n30 VSS 0.0308f
C21573 VDD96.n31 VSS 0.0286f
C21574 VDD96.n32 VSS 0.0215f
C21575 VDD96.n33 VSS 0.0586f
C21576 VDD96.n34 VSS 0.0667f
C21577 VDD96.t143 VSS 0.00622f
C21578 VDD96.n35 VSS 0.0286f
C21579 VDD96.n36 VSS 0.0215f
C21580 VDD96.n37 VSS 0.0386f
C21581 VDD96.t142 VSS 0.075f
C21582 VDD96.t136 VSS 0.0821f
C21583 VDD96.t272 VSS 0.075f
C21584 VDD96.n38 VSS 0.0386f
C21585 VDD96.n39 VSS 0.0215f
C21586 VDD96.n40 VSS 0.0286f
C21587 VDD96.n41 VSS 0.0308f
C21588 VDD96.t84 VSS 0.00622f
C21589 VDD96.n42 VSS 0.0271f
C21590 VDD96.n43 VSS 0.0215f
C21591 VDD96.n44 VSS 0.0386f
C21592 VDD96.t83 VSS 0.075f
C21593 VDD96.t329 VSS 0.0915f
C21594 VDD96.t73 VSS 0.0425f
C21595 VDD96.n45 VSS 0.0909f
C21596 VDD96.t57 VSS 0.00619f
C21597 VDD96.t357 VSS 0.0506f
C21598 VDD96.t350 VSS 0.0836f
C21599 VDD96.n46 VSS 0.0655f
C21600 VDD96.n47 VSS 0.00622f
C21601 VDD96.t145 VSS 0.00622f
C21602 VDD96.t144 VSS 0.0499f
C21603 VDD96.t160 VSS 0.0502f
C21604 VDD96.n48 VSS 0.0655f
C21605 VDD96.n49 VSS 0.00621f
C21606 VDD96.t354 VSS 0.00256f
C21607 VDD96.n50 VSS 0.00256f
C21608 VDD96.n51 VSS 0.00558f
C21609 VDD96.t353 VSS 0.0833f
C21610 VDD96.t102 VSS 0.0529f
C21611 VDD96.t46 VSS 0.0337f
C21612 VDD96.n52 VSS 0.0625f
C21613 VDD96.t12 VSS 0.00622f
C21614 VDD96.n53 VSS 0.00622f
C21615 VDD96.t11 VSS 0.103f
C21616 VDD96.t22 VSS 0.103f
C21617 VDD96.n54 VSS 0.0625f
C21618 VDD96.n55 VSS 0.00621f
C21619 VDD96.t93 VSS 0.00621f
C21620 VDD96.t15 VSS 0.0334f
C21621 VDD96.t92 VSS 0.0337f
C21622 VDD96.n56 VSS 0.0625f
C21623 VDD96.t33 VSS 0.00622f
C21624 VDD96.n57 VSS 0.00622f
C21625 VDD96.t32 VSS 0.103f
C21626 VDD96.t193 VSS 0.103f
C21627 VDD96.n58 VSS 0.0625f
C21628 VDD96.t349 VSS 0.00256f
C21629 VDD96.n59 VSS 0.00256f
C21630 VDD96.n60 VSS 0.00558f
C21631 VDD96.t28 VSS 0.00621f
C21632 VDD96.t348 VSS 0.0334f
C21633 VDD96.t27 VSS 0.0529f
C21634 VDD96.t53 VSS 0.0836f
C21635 VDD96.n61 VSS 0.0655f
C21636 VDD96.n62 VSS 0.00622f
C21637 VDD96.t332 VSS 0.00622f
C21638 VDD96.t331 VSS 0.0499f
C21639 VDD96.t29 VSS 0.0502f
C21640 VDD96.n63 VSS 0.0655f
C21641 VDD96.t45 VSS 0.00621f
C21642 VDD96.t339 VSS 0.00621f
C21643 VDD96.t94 VSS 0.0751f
C21644 VDD96.n64 VSS 0.00622f
C21645 VDD96.t287 VSS 0.00256f
C21646 VDD96.n65 VSS 0.00256f
C21647 VDD96.n66 VSS 0.00558f
C21648 VDD96.n67 VSS 0.00622f
C21649 VDD96.n68 VSS 0.0364f
C21650 VDD96.t156 VSS 0.0749f
C21651 VDD96.n69 VSS 0.00622f
C21652 VDD96.t384 VSS 0.00404f
C21653 VDD96.t155 VSS 0.00533f
C21654 VDD96.n70 VSS 0.0105f
C21655 VDD96.n71 VSS 0.00809f
C21656 VDD96.t379 VSS 0.00404f
C21657 VDD96.t159 VSS 0.00533f
C21658 VDD96.n72 VSS 0.0105f
C21659 VDD96.n73 VSS 0.043f
C21660 VDD96.n74 VSS 0.029f
C21661 VDD96.t356 VSS 0.00256f
C21662 VDD96.n75 VSS 0.00256f
C21663 VDD96.n76 VSS 0.00558f
C21664 VDD96.n77 VSS 0.0355f
C21665 VDD96.n78 VSS 0.0192f
C21666 VDD96.n79 VSS 0.0386f
C21667 VDD96.t355 VSS 0.0424f
C21668 VDD96.t340 VSS 0.0915f
C21669 VDD96.t89 VSS 0.0751f
C21670 VDD96.t190 VSS 0.0915f
C21671 VDD96.t286 VSS 0.0424f
C21672 VDD96.n80 VSS 0.0386f
C21673 VDD96.n81 VSS 0.0192f
C21674 VDD96.n82 VSS 0.0355f
C21675 VDD96.n83 VSS 0.0362f
C21676 VDD96.t26 VSS 0.00621f
C21677 VDD96.n84 VSS 0.00622f
C21678 VDD96.n85 VSS 0.0286f
C21679 VDD96.n86 VSS 0.0308f
C21680 VDD96.n87 VSS 0.0215f
C21681 VDD96.n88 VSS 0.0386f
C21682 VDD96.t25 VSS 0.082f
C21683 VDD96.t97 VSS 0.0751f
C21684 VDD96.t338 VSS 0.0808f
C21685 VDD96.n89 VSS 0.0386f
C21686 VDD96.n90 VSS 0.0215f
C21687 VDD96.n91 VSS 0.053f
C21688 VDD96.n92 VSS 0.0594f
C21689 VDD96.t44 VSS 0.0833f
C21690 VDD96.t60 VSS 0.138f
C21691 VDD96.t61 VSS 0.00622f
C21692 VDD96.n93 VSS 0.0241f
C21693 VDD96.n94 VSS 0.018f
C21694 VDD96.n95 VSS 0.0243f
C21695 VDD96.n96 VSS 0.0246f
C21696 VDD96.n97 VSS 0.0201f
C21697 VDD96.n98 VSS 0.0289f
C21698 VDD96.n99 VSS 0.0262f
C21699 VDD96.n100 VSS 0.0301f
C21700 VDD96.n101 VSS 0.0319f
C21701 VDD96.n102 VSS 0.0339f
C21702 VDD96.n103 VSS 0.0138f
C21703 VDD96.n104 VSS 0.0291f
C21704 VDD96.n105 VSS 0.0291f
C21705 VDD96.n106 VSS 0.0139f
C21706 VDD96.n107 VSS 0.0338f
C21707 VDD96.n108 VSS 0.032f
C21708 VDD96.n109 VSS 0.03f
C21709 VDD96.n110 VSS 0.0262f
C21710 VDD96.n111 VSS 0.029f
C21711 VDD96.n112 VSS 0.02f
C21712 VDD96.n113 VSS 0.0246f
C21713 VDD96.n114 VSS 0.0244f
C21714 VDD96.n115 VSS 0.018f
C21715 VDD96.n116 VSS 0.00648f
C21716 VDD96.n117 VSS 0.0411f
C21717 VDD96.n118 VSS 0.00657f
C21718 VDD96.n119 VSS 0.0419f
C21719 VDD96.n120 VSS 0.00621f
C21720 VDD96.t365 VSS 0.081f
C21721 VDD96.n121 VSS 0.0386f
C21722 VDD96.t109 VSS 0.00622f
C21723 VDD96.n122 VSS 0.00621f
C21724 VDD96.t108 VSS 0.075f
C21725 VDD96.t105 VSS 0.0821f
C21726 VDD96.n123 VSS 0.0386f
C21727 VDD96.t19 VSS 0.00622f
C21728 VDD96.t14 VSS 0.00256f
C21729 VDD96.n124 VSS 0.00256f
C21730 VDD96.n125 VSS 0.00558f
C21731 VDD96.t18 VSS 0.075f
C21732 VDD96.t13 VSS 0.0915f
C21733 VDD96.t291 VSS 0.0425f
C21734 VDD96.n126 VSS 0.0386f
C21735 VDD96.t101 VSS 0.00622f
C21736 VDD96.t369 VSS 0.00256f
C21737 VDD96.n127 VSS 0.00256f
C21738 VDD96.n128 VSS 0.00558f
C21739 VDD96.t100 VSS 0.075f
C21740 VDD96.t368 VSS 0.0915f
C21741 VDD96.t62 VSS 0.0425f
C21742 VDD96.t170 VSS 0.0748f
C21743 VDD96.n129 VSS 0.0386f
C21744 VDD96.t171 VSS 0.00581f
C21745 VDD96.n130 VSS 0.00161f
C21746 VDD96.t169 VSS 0.00518f
C21747 VDD96.n131 VSS 0.00512f
C21748 VDD96.t344 VSS 0.00256f
C21749 VDD96.n132 VSS 0.00256f
C21750 VDD96.n133 VSS 0.00558f
C21751 VDD96.n134 VSS 0.0333f
C21752 VDD96.t151 VSS 0.00622f
C21753 VDD96.t306 VSS 0.0442f
C21754 VDD96.n135 VSS 0.00621f
C21755 VDD96.t307 VSS 0.00622f
C21756 VDD96.n136 VSS 0.00621f
C21757 VDD96.n137 VSS 0.0308f
C21758 VDD96.t345 VSS 0.0653f
C21759 VDD96.n138 VSS 0.00621f
C21760 VDD96.n139 VSS 0.00621f
C21761 VDD96.t326 VSS 0.081f
C21762 VDD96.n140 VSS 0.0386f
C21763 VDD96.t242 VSS 0.00622f
C21764 VDD96.n141 VSS 0.00621f
C21765 VDD96.t241 VSS 0.075f
C21766 VDD96.t238 VSS 0.0821f
C21767 VDD96.n142 VSS 0.0386f
C21768 VDD96.t300 VSS 0.00622f
C21769 VDD96.t305 VSS 0.00256f
C21770 VDD96.n143 VSS 0.00256f
C21771 VDD96.n144 VSS 0.00558f
C21772 VDD96.t299 VSS 0.075f
C21773 VDD96.t304 VSS 0.0915f
C21774 VDD96.t288 VSS 0.0425f
C21775 VDD96.n145 VSS 0.0386f
C21776 VDD96.t5 VSS 0.00622f
C21777 VDD96.t320 VSS 0.00256f
C21778 VDD96.n146 VSS 0.00256f
C21779 VDD96.n147 VSS 0.00558f
C21780 VDD96.t4 VSS 0.075f
C21781 VDD96.t319 VSS 0.0915f
C21782 VDD96.t222 VSS 0.0425f
C21783 VDD96.t167 VSS 0.0748f
C21784 VDD96.n148 VSS 0.0386f
C21785 VDD96.t168 VSS 0.00622f
C21786 VDD96.t149 VSS 0.00533f
C21787 VDD96.t382 VSS 0.00404f
C21788 VDD96.n149 VSS 0.0105f
C21789 VDD96.t166 VSS 0.00533f
C21790 VDD96.t378 VSS 0.00404f
C21791 VDD96.n150 VSS 0.0105f
C21792 VDD96.n151 VSS 0.00872f
C21793 VDD96.n152 VSS 0.0456f
C21794 VDD96.n153 VSS 0.0289f
C21795 VDD96.n154 VSS 0.0193f
C21796 VDD96.n155 VSS 0.0354f
C21797 VDD96.n156 VSS 0.0364f
C21798 VDD96.n157 VSS 0.0193f
C21799 VDD96.n158 VSS 0.0354f
C21800 VDD96.n159 VSS 0.0363f
C21801 VDD96.n160 VSS 0.0215f
C21802 VDD96.n161 VSS 0.0308f
C21803 VDD96.n162 VSS 0.0286f
C21804 VDD96.n163 VSS 0.0215f
C21805 VDD96.n164 VSS 0.0538f
C21806 VDD96.t322 VSS 0.00619f
C21807 VDD96.t148 VSS 0.00622f
C21808 VDD96.n165 VSS 0.033f
C21809 VDD96.t321 VSS 0.0549f
C21810 VDD96.t323 VSS 0.0425f
C21811 VDD96.t80 VSS 0.00256f
C21812 VDD96.n166 VSS 0.00256f
C21813 VDD96.n167 VSS 0.00558f
C21814 VDD96.t82 VSS 0.00622f
C21815 VDD96.n168 VSS 0.00621f
C21816 VDD96.n169 VSS 0.0308f
C21817 VDD96.t258 VSS 0.0821f
C21818 VDD96.n170 VSS 0.00621f
C21819 VDD96.t1 VSS 0.00622f
C21820 VDD96.n171 VSS 0.00621f
C21821 VDD96.n172 VSS 0.00621f
C21822 VDD96.t65 VSS 0.081f
C21823 VDD96.n173 VSS 0.0386f
C21824 VDD96.t52 VSS 0.00622f
C21825 VDD96.n174 VSS 0.00621f
C21826 VDD96.t51 VSS 0.075f
C21827 VDD96.t261 VSS 0.0821f
C21828 VDD96.n175 VSS 0.0386f
C21829 VDD96.t208 VSS 0.00622f
C21830 VDD96.t203 VSS 0.00256f
C21831 VDD96.n176 VSS 0.00256f
C21832 VDD96.n177 VSS 0.00558f
C21833 VDD96.t207 VSS 0.075f
C21834 VDD96.t202 VSS 0.0915f
C21835 VDD96.t280 VSS 0.0425f
C21836 VDD96.n178 VSS 0.0386f
C21837 VDD96.t88 VSS 0.00622f
C21838 VDD96.t59 VSS 0.00256f
C21839 VDD96.n179 VSS 0.00256f
C21840 VDD96.n180 VSS 0.00558f
C21841 VDD96.t87 VSS 0.075f
C21842 VDD96.t58 VSS 0.0915f
C21843 VDD96.t316 VSS 0.0425f
C21844 VDD96.t173 VSS 0.0748f
C21845 VDD96.n181 VSS 0.0386f
C21846 VDD96.t174 VSS 0.00622f
C21847 VDD96.t146 VSS 0.00533f
C21848 VDD96.t385 VSS 0.00404f
C21849 VDD96.n182 VSS 0.0105f
C21850 VDD96.t172 VSS 0.00533f
C21851 VDD96.t375 VSS 0.00404f
C21852 VDD96.n183 VSS 0.0105f
C21853 VDD96.n184 VSS 0.00796f
C21854 VDD96.n185 VSS 0.0434f
C21855 VDD96.n186 VSS 0.0289f
C21856 VDD96.n187 VSS 0.0193f
C21857 VDD96.n188 VSS 0.0354f
C21858 VDD96.n189 VSS 0.0364f
C21859 VDD96.n190 VSS 0.0193f
C21860 VDD96.n191 VSS 0.0354f
C21861 VDD96.n192 VSS 0.0363f
C21862 VDD96.n193 VSS 0.0215f
C21863 VDD96.n194 VSS 0.0308f
C21864 VDD96.n195 VSS 0.0286f
C21865 VDD96.n196 VSS 0.0215f
C21866 VDD96.n197 VSS 0.0586f
C21867 VDD96.n198 VSS 0.0667f
C21868 VDD96.t76 VSS 0.081f
C21869 VDD96.t0 VSS 0.075f
C21870 VDD96.n199 VSS 0.0386f
C21871 VDD96.n200 VSS 0.0215f
C21872 VDD96.n201 VSS 0.0286f
C21873 VDD96.n202 VSS 0.0308f
C21874 VDD96.t201 VSS 0.00622f
C21875 VDD96.n203 VSS 0.0286f
C21876 VDD96.n204 VSS 0.0215f
C21877 VDD96.n205 VSS 0.0386f
C21878 VDD96.t200 VSS 0.075f
C21879 VDD96.t204 VSS 0.0821f
C21880 VDD96.t79 VSS 0.0915f
C21881 VDD96.t81 VSS 0.075f
C21882 VDD96.n206 VSS 0.0386f
C21883 VDD96.n207 VSS 0.0215f
C21884 VDD96.n208 VSS 0.0271f
C21885 VDD96.n209 VSS 0.0254f
C21886 VDD96.n210 VSS 0.0193f
C21887 VDD96.n211 VSS 0.0386f
C21888 VDD96.t147 VSS 0.0425f
C21889 VDD96.n212 VSS 0.0577f
C21890 VDD96.n213 VSS 0.0305f
C21891 VDD96.n214 VSS 0.0516f
C21892 VDD96.n215 VSS 0.0301f
C21893 VDD96.t315 VSS 0.00622f
C21894 VDD96.n216 VSS 0.0286f
C21895 VDD96.n217 VSS 0.0215f
C21896 VDD96.n218 VSS 0.0333f
C21897 VDD96.t314 VSS 0.0596f
C21898 VDD96.t235 VSS 0.0653f
C21899 VDD96.n219 VSS 0.0333f
C21900 VDD96.n220 VSS 0.0215f
C21901 VDD96.n221 VSS 0.0286f
C21902 VDD96.n222 VSS 0.0308f
C21903 VDD96.t234 VSS 0.00622f
C21904 VDD96.n223 VSS 0.0271f
C21905 VDD96.n224 VSS 0.0215f
C21906 VDD96.t230 VSS 0.0338f
C21907 VDD96.t343 VSS 0.0728f
C21908 VDD96.t233 VSS 0.0596f
C21909 VDD96.n225 VSS 0.0333f
C21910 VDD96.t301 VSS 0.0287f
C21911 VDD96.n226 VSS 0.172f
C21912 VDD96.t150 VSS 0.0338f
C21913 VDD96.n227 VSS 0.0953f
C21914 VDD96.t225 VSS 0.0685f
C21915 VDD96.t226 VSS 0.00619f
C21916 VDD96.n228 VSS 0.00619f
C21917 VDD96.t123 VSS 0.0313f
C21918 VDD96.n229 VSS 0.00618f
C21919 VDD96.t38 VSS 0.0821f
C21920 VDD96.n230 VSS 0.0646f
C21921 VDD96.n231 VSS 0.00619f
C21922 VDD96.t86 VSS 0.00618f
C21923 VDD96.t85 VSS 0.049f
C21924 VDD96.t179 VSS 0.0493f
C21925 VDD96.n232 VSS 0.0646f
C21926 VDD96.n233 VSS 0.00618f
C21927 VDD96.t337 VSS 0.00256f
C21928 VDD96.n234 VSS 0.00256f
C21929 VDD96.n235 VSS 0.00554f
C21930 VDD96.t336 VSS 0.0818f
C21931 VDD96.t209 VSS 0.0519f
C21932 VDD96.t6 VSS 0.0331f
C21933 VDD96.n236 VSS 0.0616f
C21934 VDD96.t275 VSS 0.00618f
C21935 VDD96.n237 VSS 0.00619f
C21936 VDD96.t274 VSS 0.101f
C21937 VDD96.t128 VSS 0.101f
C21938 VDD96.n238 VSS 0.0616f
C21939 VDD96.n239 VSS 0.00618f
C21940 VDD96.t252 VSS 0.00618f
C21941 VDD96.t245 VSS 0.0328f
C21942 VDD96.t251 VSS 0.0331f
C21943 VDD96.n240 VSS 0.0616f
C21944 VDD96.t3 VSS 0.00618f
C21945 VDD96.n241 VSS 0.00619f
C21946 VDD96.t2 VSS 0.101f
C21947 VDD96.t267 VSS 0.101f
C21948 VDD96.n242 VSS 0.0616f
C21949 VDD96.t37 VSS 0.00256f
C21950 VDD96.n243 VSS 0.00256f
C21951 VDD96.n244 VSS 0.00554f
C21952 VDD96.t189 VSS 0.00618f
C21953 VDD96.t36 VSS 0.0328f
C21954 VDD96.t188 VSS 0.0519f
C21955 VDD96.t120 VSS 0.0821f
C21956 VDD96.n245 VSS 0.0646f
C21957 VDD96.n246 VSS 0.00619f
C21958 VDD96.t165 VSS 0.00618f
C21959 VDD96.t164 VSS 0.049f
C21960 VDD96.t217 VSS 0.0493f
C21961 VDD96.n247 VSS 0.0646f
C21962 VDD96.t10 VSS 0.00618f
C21963 VDD96.t9 VSS 0.0818f
C21964 VDD96.t113 VSS 0.0314f
C21965 VDD96.t114 VSS 0.00619f
C21966 VDD96.t116 VSS 0.00621f
C21967 VDD96.t253 VSS 0.0751f
C21968 VDD96.n248 VSS 0.00622f
C21969 VDD96.t285 VSS 0.00256f
C21970 VDD96.n249 VSS 0.00256f
C21971 VDD96.n250 VSS 0.00558f
C21972 VDD96.n251 VSS 0.00622f
C21973 VDD96.n252 VSS 0.0364f
C21974 VDD96.t183 VSS 0.0749f
C21975 VDD96.n253 VSS 0.00622f
C21976 VDD96.t374 VSS 0.00404f
C21977 VDD96.t182 VSS 0.00533f
C21978 VDD96.n254 VSS 0.0105f
C21979 VDD96.n255 VSS 0.00774f
C21980 VDD96.t370 VSS 0.00404f
C21981 VDD96.t178 VSS 0.00533f
C21982 VDD96.n256 VSS 0.0105f
C21983 VDD96.n257 VSS 0.0047f
C21984 VDD96.n258 VSS 0.00376f
C21985 VDD96.n259 VSS 0.0381f
C21986 VDD96.n260 VSS 0.029f
C21987 VDD96.t127 VSS 0.00256f
C21988 VDD96.n261 VSS 0.00256f
C21989 VDD96.n262 VSS 0.00558f
C21990 VDD96.n263 VSS 0.0355f
C21991 VDD96.n264 VSS 0.0192f
C21992 VDD96.n265 VSS 0.0386f
C21993 VDD96.t126 VSS 0.0424f
C21994 VDD96.t117 VSS 0.0915f
C21995 VDD96.t248 VSS 0.0751f
C21996 VDD96.t264 VSS 0.0915f
C21997 VDD96.t284 VSS 0.0424f
C21998 VDD96.n266 VSS 0.0386f
C21999 VDD96.n267 VSS 0.0192f
C22000 VDD96.n268 VSS 0.0355f
C22001 VDD96.n269 VSS 0.0362f
C22002 VDD96.t187 VSS 0.00621f
C22003 VDD96.n270 VSS 0.00622f
C22004 VDD96.n271 VSS 0.0286f
C22005 VDD96.n272 VSS 0.0308f
C22006 VDD96.n273 VSS 0.0215f
C22007 VDD96.n274 VSS 0.0386f
C22008 VDD96.t186 VSS 0.082f
C22009 VDD96.t41 VSS 0.0751f
C22010 VDD96.t115 VSS 0.0808f
C22011 VDD96.n275 VSS 0.0386f
C22012 VDD96.n276 VSS 0.0215f
C22013 VDD96.n277 VSS 0.0544f
C22014 VDD96.n278 VSS 0.0689f
C22015 VDD96.n279 VSS 0.036f
C22016 VDD96.n280 VSS 0.0316f
C22017 VDD96.n281 VSS 0.024f
C22018 VDD96.n282 VSS 0.0243f
C22019 VDD96.n283 VSS 0.0202f
C22020 VDD96.n284 VSS 0.0287f
C22021 VDD96.n285 VSS 0.026f
C22022 VDD96.n286 VSS 0.0302f
C22023 VDD96.n287 VSS 0.0317f
C22024 VDD96.n288 VSS 0.0337f
C22025 VDD96.n289 VSS 0.0138f
C22026 VDD96.n290 VSS 0.0289f
C22027 VDD96.n291 VSS 0.0289f
C22028 VDD96.n292 VSS 0.0139f
C22029 VDD96.n293 VSS 0.0336f
C22030 VDD96.n294 VSS 0.0317f
C22031 VDD96.n295 VSS 0.0301f
C22032 VDD96.n296 VSS 0.026f
C22033 VDD96.n297 VSS 0.0288f
C22034 VDD96.n298 VSS 0.02f
C22035 VDD96.n299 VSS 0.0243f
C22036 VDD96.n300 VSS 0.0241f
C22037 VDD96.n301 VSS 0.0315f
C22038 VDD96.n302 VSS 0.0361f
C22039 VDD96.n303 VSS 0.038f
C22040 VDD96.n304 VSS 0.00621f
C22041 VDD96.t227 VSS 0.081f
C22042 VDD96.n305 VSS 0.0386f
C22043 VDD96.t216 VSS 0.00622f
C22044 VDD96.n306 VSS 0.00621f
C22045 VDD96.t215 VSS 0.075f
C22046 VDD96.t212 VSS 0.0821f
C22047 VDD96.n307 VSS 0.0386f
C22048 VDD96.t244 VSS 0.00622f
C22049 VDD96.t277 VSS 0.00256f
C22050 VDD96.n308 VSS 0.00256f
C22051 VDD96.n309 VSS 0.00558f
C22052 VDD96.t243 VSS 0.075f
C22053 VDD96.t276 VSS 0.0915f
C22054 VDD96.t278 VSS 0.0425f
C22055 VDD96.n310 VSS 0.0386f
C22056 VDD96.t298 VSS 0.00622f
C22057 VDD96.t221 VSS 0.00256f
C22058 VDD96.n311 VSS 0.00256f
C22059 VDD96.n312 VSS 0.00558f
C22060 VDD96.t297 VSS 0.075f
C22061 VDD96.t220 VSS 0.0915f
C22062 VDD96.t110 VSS 0.0425f
C22063 VDD96.t153 VSS 0.0748f
C22064 VDD96.n313 VSS 0.0386f
C22065 VDD96.t154 VSS 0.00622f
C22066 VDD96.t163 VSS 0.00533f
C22067 VDD96.t372 VSS 0.00404f
C22068 VDD96.n314 VSS 0.0105f
C22069 VDD96.n315 VSS 0.00965f
C22070 VDD96.t152 VSS 0.00533f
C22071 VDD96.t380 VSS 0.00404f
C22072 VDD96.n316 VSS 0.0104f
C22073 VDD96.n317 VSS 0.00417f
C22074 VDD96.n318 VSS 4.32e-19
C22075 VDD96.n319 VSS 0.00277f
C22076 VDD96.n320 VSS 0.0438f
C22077 VDD96.n321 VSS 0.0289f
C22078 VDD96.n322 VSS 0.0193f
C22079 VDD96.n323 VSS 0.0354f
C22080 VDD96.n324 VSS 0.0364f
C22081 VDD96.n325 VSS 0.0193f
C22082 VDD96.n326 VSS 0.0354f
C22083 VDD96.n327 VSS 0.0363f
C22084 VDD96.n328 VSS 0.0215f
C22085 VDD96.n329 VSS 0.0308f
C22086 VDD96.n330 VSS 0.0286f
C22087 VDD96.n331 VSS 0.0215f
C22088 VDD96.n332 VSS 0.0542f
C22089 VDD96.n333 VSS 0.0489f
C22090 VDD96.n334 VSS 0.0343f
C22091 VDD96.n335 VSS 0.0329f
C22092 VDD96.n336 VSS 0.0193f
C22093 VDD96.n337 VSS 0.0232f
C22094 VDD96.n338 VSS 0.0105f
C22095 VDD96.t175 VSS 0.00533f
C22096 VDD96.t371 VSS 0.00404f
C22097 VDD96.n339 VSS 0.0104f
C22098 VDD96.n340 VSS 0.0442f
C22099 VDD96.n341 VSS 0.0854f
C22100 VDD96.n342 VSS 0.0173f
C22101 VDD96.n343 VSS 5.16e-20
C22102 VDD96.n344 VSS 0.00136f
C22103 VDD96.t377 VSS 0.00403f
C22104 VDD96.n345 VSS 0.00547f
C22105 VDD96.n346 VSS 7.4e-19
C22106 VDD96.n347 VSS 6.15e-19
C22107 VDD96.n348 VSS 0.00462f
C22108 VDD96.n349 VSS 0.0145f
C22109 VDD96.n350 VSS 0.0355f
C22110 VDD96.n351 VSS 0.0354f
C22111 VDD96.n352 VSS 0.0364f
C22112 VDD96.n353 VSS 0.0193f
C22113 VDD96.n354 VSS 0.0354f
C22114 VDD96.n355 VSS 0.0363f
C22115 VDD96.n356 VSS 0.0215f
C22116 VDD96.n357 VSS 0.0308f
C22117 VDD96.n358 VSS 0.0286f
C22118 VDD96.n359 VSS 0.0215f
C22119 VDD96.n360 VSS 0.0551f
C22120 VDD96.n361 VSS 0.0457f
C22121 VDD96.n362 VSS 0.0245f
C22122 VDD96.n363 VSS 0.0829f
C22123 VDD96.t56 VSS 0.0629f
C22124 VDD96.n364 VSS 0.054f
C22125 VDD96.t360 VSS 0.0377f
C22126 VDD96.n365 VSS 0.0386f
C22127 VDD96.n366 VSS 0.0143f
C22128 VDD96.n367 VSS 0.0485f
C22129 VDD96.n368 VSS 0.0517f
C22130 VDD96.n369 VSS 0.0241f
C22131 VDD96.n370 VSS 0.0357f
C22132 VDD96.n371 VSS 0.0316f
C22133 VDD96.n372 VSS 0.0452f
C22134 VDD96.n373 VSS 0.037f
C22135 VDD96.n374 VSS 0.0593f
C22136 VDD96.n375 VSS 0.00183f
C22137 VDD96.n376 VSS 0.0062f
C22138 VDD96.n377 VSS 0.0156f
C22139 RST.n0 VSS 0.116f
C22140 RST.n1 VSS 7.03e-19
C22141 RST.n2 VSS 6.62e-19
C22142 RST.t27 VSS 0.00542f
C22143 RST.n3 VSS 0.00496f
C22144 RST.n4 VSS 0.00191f
C22145 RST.t41 VSS 0.00861f
C22146 RST.n5 VSS 0.0106f
C22147 RST.n6 VSS 8.34e-20
C22148 RST.n7 VSS 7e-19
C22149 RST.n8 VSS 0.00439f
C22150 RST.n9 VSS 0.00351f
C22151 RST.t114 VSS 0.00568f
C22152 RST.t122 VSS 0.00863f
C22153 RST.n10 VSS 0.0153f
C22154 RST.n11 VSS 0.00822f
C22155 RST.t82 VSS 0.00568f
C22156 RST.t104 VSS 0.00863f
C22157 RST.n12 VSS 0.0153f
C22158 RST.n13 VSS 0.0832f
C22159 RST.n14 VSS 0.259f
C22160 RST.n15 VSS 0.162f
C22161 RST.t42 VSS 0.00568f
C22162 RST.t53 VSS 0.00863f
C22163 RST.n16 VSS 0.0153f
C22164 RST.n17 VSS 0.00795f
C22165 RST.n18 VSS 0.307f
C22166 RST.n19 VSS 8.9e-19
C22167 RST.n20 VSS 0.00267f
C22168 RST.t29 VSS 0.00863f
C22169 RST.t120 VSS 0.00568f
C22170 RST.n21 VSS 0.0152f
C22171 RST.n22 VSS 0.00199f
C22172 RST.n23 VSS 7.14e-19
C22173 RST.n24 VSS 0.0566f
C22174 RST.n25 VSS 0.00248f
C22175 RST.t26 VSS 0.00872f
C22176 RST.t116 VSS 0.00552f
C22177 RST.n26 VSS 0.0153f
C22178 RST.n27 VSS 0.00199f
C22179 RST.n28 VSS 0.00132f
C22180 RST.n29 VSS 7.02e-19
C22181 RST.n30 VSS 0.034f
C22182 RST.n31 VSS 0.398f
C22183 RST.n32 VSS 8.9e-19
C22184 RST.n33 VSS 0.00267f
C22185 RST.t6 VSS 0.00863f
C22186 RST.t101 VSS 0.00568f
C22187 RST.n34 VSS 0.0152f
C22188 RST.n35 VSS 0.00199f
C22189 RST.n36 VSS 7.14e-19
C22190 RST.n37 VSS 0.0566f
C22191 RST.n38 VSS 0.35f
C22192 RST.n39 VSS 0.24f
C22193 RST.t49 VSS 0.00552f
C22194 RST.t93 VSS 0.00872f
C22195 RST.n40 VSS 0.0153f
C22196 RST.n41 VSS 0.00199f
C22197 RST.n42 VSS 0.00132f
C22198 RST.n43 VSS 7.02e-19
C22199 RST.n44 VSS 0.00248f
C22200 RST.n45 VSS 0.021f
C22201 RST.n46 VSS 0.114f
C22202 RST.n47 VSS 0.289f
C22203 RST.n48 VSS 0.142f
C22204 RST.n49 VSS 0.245f
C22205 RST.n50 VSS 0.0103f
C22206 RST.n51 VSS 0.131f
C22207 RST.n52 VSS 0.0147f
C22208 RST.t45 VSS 0.00568f
C22209 RST.t23 VSS 0.00863f
C22210 RST.n53 VSS 0.0152f
C22211 RST.n54 VSS 0.00267f
C22212 RST.n55 VSS 0.00196f
C22213 RST.n56 VSS 9.12e-19
C22214 RST.n57 VSS 7.14e-19
C22215 RST.n58 VSS 0.0568f
C22216 RST.n59 VSS 0.00256f
C22217 RST.n60 VSS 0.00132f
C22218 RST.t110 VSS 0.0087f
C22219 RST.t2 VSS 0.00554f
C22220 RST.n61 VSS 0.0153f
C22221 RST.n62 VSS 0.00196f
C22222 RST.n63 VSS 7.02e-19
C22223 RST.n64 VSS 0.032f
C22224 RST.n65 VSS 0.00249f
C22225 RST.n66 VSS 0.0013f
C22226 RST.t88 VSS 0.00568f
C22227 RST.t66 VSS 0.00863f
C22228 RST.n67 VSS 0.0152f
C22229 RST.n68 VSS 0.00202f
C22230 RST.n69 VSS 7.02e-19
C22231 RST.n70 VSS 0.00108f
C22232 RST.n71 VSS 0.004f
C22233 RST.n72 VSS 0.0749f
C22234 RST.t86 VSS 0.00863f
C22235 RST.t85 VSS 0.00568f
C22236 RST.n73 VSS 0.0153f
C22237 RST.n74 VSS 0.0882f
C22238 RST.n75 VSS 0.136f
C22239 RST.n76 VSS 9.45e-19
C22240 RST.t89 VSS 0.00568f
C22241 RST.t34 VSS 0.00863f
C22242 RST.n77 VSS 0.0152f
C22243 RST.n78 VSS 0.00253f
C22244 RST.n79 VSS 7.02e-19
C22245 RST.n80 VSS 0.00196f
C22246 RST.n81 VSS 0.00265f
C22247 RST.n82 VSS 0.00111f
C22248 RST.n83 VSS 0.00269f
C22249 RST.n84 VSS 0.149f
C22250 RST.n85 VSS 0.143f
C22251 RST.n86 VSS 0.00269f
C22252 RST.n87 VSS 0.00127f
C22253 RST.t60 VSS 0.00568f
C22254 RST.t44 VSS 0.00863f
C22255 RST.n88 VSS 0.0152f
C22256 RST.n89 VSS 0.00202f
C22257 RST.n90 VSS 7.56e-19
C22258 RST.n91 VSS 9.93e-19
C22259 RST.n92 VSS 0.00363f
C22260 RST.n93 VSS 2.07e-19
C22261 RST.n94 VSS 0.00147f
C22262 RST.n95 VSS 0.00143f
C22263 RST.n96 VSS 0.0692f
C22264 RST.n97 VSS 0.23f
C22265 RST.n98 VSS 0.407f
C22266 RST.n99 VSS 0.00215f
C22267 RST.t87 VSS 0.00863f
C22268 RST.t77 VSS 0.00568f
C22269 RST.n100 VSS 0.0152f
C22270 RST.n101 VSS 0.00199f
C22271 RST.n102 VSS 0.00132f
C22272 RST.n103 VSS 7.02e-19
C22273 RST.n104 VSS 9.32e-19
C22274 RST.n105 VSS 0.00385f
C22275 RST.n106 VSS 0.224f
C22276 RST.n107 VSS 0.00245f
C22277 RST.n108 VSS 0.101f
C22278 RST.n109 VSS 0.362f
C22279 RST.n110 VSS 0.041f
C22280 RST.n111 VSS 0.22f
C22281 RST.t80 VSS 0.00863f
C22282 RST.t119 VSS 0.00568f
C22283 RST.n112 VSS 0.0152f
C22284 RST.n113 VSS 0.00207f
C22285 RST.n114 VSS 0.00127f
C22286 RST.n115 VSS 7.02e-19
C22287 RST.n116 VSS 0.00155f
C22288 RST.n117 VSS 9.55e-19
C22289 RST.n118 VSS 0.00389f
C22290 RST.n119 VSS 0.0663f
C22291 RST.n120 VSS 0.00282f
C22292 RST.n121 VSS 0.00101f
C22293 RST.n122 VSS 7.83e-19
C22294 RST.t106 VSS 0.00863f
C22295 RST.t14 VSS 0.00568f
C22296 RST.n123 VSS 0.0152f
C22297 RST.n124 VSS 0.0021f
C22298 RST.n125 VSS 0.00265f
C22299 RST.n126 VSS 0.00122f
C22300 RST.n127 VSS 0.00109f
C22301 RST.n128 VSS 8.38e-20
C22302 RST.n129 VSS 0.0038f
C22303 RST.n130 VSS 8.38e-20
C22304 RST.n131 VSS 0.0557f
C22305 RST.n132 VSS 0.177f
C22306 RST.t79 VSS 0.00568f
C22307 RST.t58 VSS 0.00863f
C22308 RST.n133 VSS 0.0152f
C22309 RST.n134 VSS 0.00267f
C22310 RST.n135 VSS 0.00102f
C22311 RST.n136 VSS 0.00314f
C22312 RST.n137 VSS 0.00374f
C22313 RST.t74 VSS 0.00568f
C22314 RST.t54 VSS 0.00863f
C22315 RST.n138 VSS 0.0153f
C22316 RST.n139 VSS 0.0841f
C22317 RST.n140 VSS 0.148f
C22318 RST.n141 VSS 0.052f
C22319 RST.t31 VSS 0.00568f
C22320 RST.t15 VSS 0.00863f
C22321 RST.n142 VSS 0.0153f
C22322 RST.n143 VSS 0.0407f
C22323 RST.n144 VSS 0.19f
C22324 RST.n145 VSS 0.00256f
C22325 RST.n146 VSS 0.00132f
C22326 RST.t46 VSS 0.0087f
C22327 RST.t32 VSS 0.00554f
C22328 RST.n147 VSS 0.0153f
C22329 RST.n148 VSS 0.00196f
C22330 RST.n149 VSS 7.02e-19
C22331 RST.n150 VSS 0.0464f
C22332 RST.t90 VSS 0.00568f
C22333 RST.t69 VSS 0.00863f
C22334 RST.n151 VSS 0.0152f
C22335 RST.n152 VSS 0.00267f
C22336 RST.n153 VSS 0.00196f
C22337 RST.n154 VSS 9.12e-19
C22338 RST.n155 VSS 7.14e-19
C22339 RST.n156 VSS 0.0495f
C22340 RST.n157 VSS 0.278f
C22341 RST.n158 VSS 0.0572f
C22342 RST.n159 VSS 0.00585f
C22343 RST.n160 VSS 0.00291f
C22344 RST.n161 VSS 0.00968f
C22345 RST.n162 VSS 0.0334f
C22346 RST.n163 VSS 0.00621f
C22347 RST.n164 VSS 0.0029f
C22348 RST.n165 VSS 0.0355f
C22349 RST.n166 VSS 0.675f
C22350 RST.n167 VSS 0.757f
C22351 RST.n168 VSS 0.394f
C22352 RST.n169 VSS 0.0795f
C22353 RST.n170 VSS 0.0918f
C22354 RST.n171 VSS 4.13e-19
C22355 RST.n172 VSS 3.6e-19
C22356 RST.n173 VSS 0.00242f
C22357 RST.n174 VSS 0.00117f
C22358 RST.n175 VSS 5.4e-19
C22359 RST.n176 VSS 0.00332f
C22360 RST.n177 VSS 0.00523f
C22361 RST.n178 VSS 0.0108f
C22362 RST.n179 VSS 3.6e-19
C22363 RST.n180 VSS 0.00117f
C22364 RST.n181 VSS 0.00314f
C22365 RST.n182 VSS 0.00117f
C22366 RST.n183 VSS 8.37e-19
C22367 RST.t25 VSS 0.00568f
C22368 RST.t107 VSS 0.00863f
C22369 RST.n184 VSS 0.0152f
C22370 RST.n185 VSS 0.00215f
C22371 RST.n186 VSS 0.00409f
C22372 RST.n187 VSS 0.217f
C22373 RST.t92 VSS 0.00568f
C22374 RST.t36 VSS 0.00863f
C22375 RST.n188 VSS 0.0152f
C22376 RST.n189 VSS 0.00279f
C22377 RST.n190 VSS 9.43e-19
C22378 RST.n191 VSS 0.00344f
C22379 RST.n192 VSS 0.217f
C22380 RST.n193 VSS 0.214f
C22381 RST.n194 VSS 0.214f
C22382 RST.n195 VSS 6.21e-19
C22383 RST.n196 VSS 0.00329f
C22384 RST.n197 VSS 6.02e-19
C22385 RST.t28 VSS 0.00568f
C22386 RST.t111 VSS 0.00863f
C22387 RST.n198 VSS 0.0152f
C22388 RST.n199 VSS 0.00228f
C22389 RST.n200 VSS 2.43e-19
C22390 RST.n201 VSS 0.00113f
C22391 RST.n202 VSS 0.213f
C22392 RST.n203 VSS 0.213f
C22393 RST.n204 VSS 0.00234f
C22394 RST.n205 VSS 9.92e-19
C22395 RST.n206 VSS 0.0032f
C22396 RST.n207 VSS 0.00122f
C22397 RST.n208 VSS 7.29e-19
C22398 RST.t57 VSS 0.00568f
C22399 RST.t8 VSS 0.00863f
C22400 RST.n209 VSS 0.0152f
C22401 RST.n210 VSS 0.00212f
C22402 RST.n211 VSS 0.00366f
C22403 RST.n212 VSS 0.0277f
C22404 RST.n213 VSS 0.0374f
C22405 RST.n214 VSS 0.00248f
C22406 RST.t43 VSS 0.00872f
C22407 RST.t95 VSS 0.00552f
C22408 RST.n215 VSS 0.0153f
C22409 RST.n216 VSS 0.00199f
C22410 RST.n217 VSS 0.00132f
C22411 RST.n218 VSS 7.02e-19
C22412 RST.n219 VSS 0.0295f
C22413 RST.n220 VSS 8.9e-19
C22414 RST.n221 VSS 0.00267f
C22415 RST.t102 VSS 0.00863f
C22416 RST.t10 VSS 0.00568f
C22417 RST.n222 VSS 0.0152f
C22418 RST.n223 VSS 0.00199f
C22419 RST.n224 VSS 7.14e-19
C22420 RST.n225 VSS 0.0566f
C22421 RST.n226 VSS 0.00248f
C22422 RST.t94 VSS 0.00872f
C22423 RST.t7 VSS 0.00552f
C22424 RST.n227 VSS 0.0153f
C22425 RST.n228 VSS 0.00199f
C22426 RST.n229 VSS 0.00132f
C22427 RST.n230 VSS 7.02e-19
C22428 RST.n231 VSS 0.034f
C22429 RST.n232 VSS 0.425f
C22430 RST.n233 VSS 8.9e-19
C22431 RST.n234 VSS 0.00267f
C22432 RST.t62 VSS 0.00863f
C22433 RST.t109 VSS 0.00568f
C22434 RST.n235 VSS 0.0152f
C22435 RST.n236 VSS 0.00199f
C22436 RST.n237 VSS 7.14e-19
C22437 RST.n238 VSS 0.0566f
C22438 RST.n239 VSS 0.381f
C22439 RST.n240 VSS 0.0703f
C22440 RST.n241 VSS 0.146f
C22441 RST.n242 VSS 8.35f
C22442 RST.n243 VSS 0.215f
C22443 RST.n244 VSS 1.24f
C22444 RST.n245 VSS 8.9e-19
C22445 RST.n246 VSS 0.00267f
C22446 RST.t59 VSS 0.00568f
C22447 RST.t55 VSS 0.00863f
C22448 RST.n247 VSS 0.0152f
C22449 RST.n248 VSS 0.00199f
C22450 RST.n249 VSS 7.14e-19
C22451 RST.n250 VSS 0.0495f
C22452 RST.n251 VSS 0.00256f
C22453 RST.t35 VSS 0.0087f
C22454 RST.t16 VSS 0.00554f
C22455 RST.n252 VSS 0.0153f
C22456 RST.n253 VSS 0.00199f
C22457 RST.n254 VSS 0.00132f
C22458 RST.n255 VSS 7.02e-19
C22459 RST.n256 VSS 0.021f
C22460 RST.n257 VSS 8.9e-19
C22461 RST.n258 VSS 0.00267f
C22462 RST.t30 VSS 0.00568f
C22463 RST.t22 VSS 0.00863f
C22464 RST.n259 VSS 0.0152f
C22465 RST.n260 VSS 0.00199f
C22466 RST.n261 VSS 7.14e-19
C22467 RST.n262 VSS 0.0495f
C22468 RST.n263 VSS 0.00248f
C22469 RST.n264 VSS 0.00132f
C22470 RST.t125 VSS 0.00552f
C22471 RST.t118 VSS 0.00872f
C22472 RST.n265 VSS 0.0153f
C22473 RST.n266 VSS 0.00196f
C22474 RST.n267 VSS 7.02e-19
C22475 RST.n268 VSS 0.0386f
C22476 RST.t73 VSS 0.00863f
C22477 RST.t81 VSS 0.00568f
C22478 RST.n269 VSS 0.0152f
C22479 RST.n270 VSS 0.00267f
C22480 RST.n271 VSS 0.00196f
C22481 RST.n272 VSS 9.12e-19
C22482 RST.n273 VSS 7.14e-19
C22483 RST.n274 VSS 0.0533f
C22484 RST.n275 VSS 0.213f
C22485 RST.n276 VSS 0.00256f
C22486 RST.t48 VSS 0.0087f
C22487 RST.t83 VSS 0.00554f
C22488 RST.n277 VSS 0.0153f
C22489 RST.n278 VSS 0.00199f
C22490 RST.n279 VSS 0.00132f
C22491 RST.n280 VSS 7.02e-19
C22492 RST.n281 VSS 0.021f
C22493 RST.n282 VSS 0.0867f
C22494 RST.n283 VSS 0.168f
C22495 RST.n284 VSS 0.155f
C22496 RST.n285 VSS 0.153f
C22497 RST.t112 VSS 0.00568f
C22498 RST.t96 VSS 0.00863f
C22499 RST.n286 VSS 0.0153f
C22500 RST.n287 VSS 0.0461f
C22501 RST.n288 VSS 0.00265f
C22502 RST.n289 VSS 0.00329f
C22503 RST.n290 VSS 0.00116f
C22504 RST.t113 VSS 0.00568f
C22505 RST.t97 VSS 0.00863f
C22506 RST.n291 VSS 0.0152f
C22507 RST.n292 VSS 0.00216f
C22508 RST.n293 VSS 8.37e-19
C22509 RST.n294 VSS 4.3e-19
C22510 RST.n295 VSS 8.99e-19
C22511 RST.n296 VSS 0.00511f
C22512 RST.n297 VSS 0.0444f
C22513 RST.n298 VSS 0.231f
C22514 RST.n299 VSS 0.154f
C22515 RST.n300 VSS 0.169f
C22516 RST.n301 VSS 0.00329f
C22517 RST.n302 VSS 6.21e-19
C22518 RST.t19 VSS 0.00568f
C22519 RST.t105 VSS 0.00863f
C22520 RST.n303 VSS 0.0152f
C22521 RST.n304 VSS 0.00228f
C22522 RST.n305 VSS 0.00117f
C22523 RST.n306 VSS 5.4e-19
C22524 RST.n307 VSS 2.43e-19
C22525 RST.n308 VSS 0.00113f
C22526 RST.n309 VSS 6.02e-19
C22527 RST.n310 VSS 0.00332f
C22528 RST.n311 VSS 0.00446f
C22529 RST.n312 VSS 7.03e-19
C22530 RST.n313 VSS 6.62e-19
C22531 RST.n314 VSS 7.06e-19
C22532 RST.n315 VSS 7.89e-20
C22533 RST.t98 VSS 0.00863f
C22534 RST.n316 VSS 0.0107f
C22535 RST.t108 VSS 0.00517f
C22536 RST.n317 VSS 0.00508f
C22537 RST.n318 VSS 0.00191f
C22538 RST.n319 VSS 0.00344f
C22539 RST.t5 VSS 0.00863f
C22540 RST.t17 VSS 0.00568f
C22541 RST.n320 VSS 0.0153f
C22542 RST.n321 VSS 0.00822f
C22543 RST.t18 VSS 0.00863f
C22544 RST.t37 VSS 0.00568f
C22545 RST.n322 VSS 0.0153f
C22546 RST.n323 VSS 0.0832f
C22547 RST.n324 VSS 0.259f
C22548 RST.n325 VSS 0.215f
C22549 RST.t71 VSS 0.00863f
C22550 RST.t91 VSS 0.00568f
C22551 RST.n326 VSS 0.0153f
C22552 RST.n327 VSS 0.00778f
C22553 RST.n328 VSS 0.0158f
C22554 RST.n329 VSS 0.104f
C22555 RST.n330 VSS 0.0642f
C22556 RST.n331 VSS 0.0276f
C22557 RST.n332 VSS 4.13e-19
C22558 RST.n333 VSS 0.0032f
C22559 RST.n334 VSS 0.00366f
C22560 RST.n335 VSS 0.00122f
C22561 RST.t50 VSS 0.00568f
C22562 RST.t4 VSS 0.00863f
C22563 RST.n336 VSS 0.0152f
C22564 RST.n337 VSS 0.00212f
C22565 RST.n338 VSS 7.29e-19
C22566 RST.n339 VSS 3.6e-19
C22567 RST.n340 VSS 9.92e-19
C22568 RST.n341 VSS 0.00234f
C22569 RST.n342 VSS 0.213f
C22570 RST.n343 VSS 0.213f
C22571 RST.n344 VSS 0.00242f
C22572 RST.n345 VSS 0.214f
C22573 RST.t123 VSS 0.00568f
C22574 RST.t72 VSS 0.00863f
C22575 RST.n346 VSS 0.0152f
C22576 RST.n347 VSS 0.00279f
C22577 RST.n348 VSS 9.43e-19
C22578 RST.n349 VSS 0.00344f
C22579 RST.n350 VSS 0.00523f
C22580 RST.n351 VSS 0.214f
C22581 RST.n352 VSS 0.217f
C22582 RST.n353 VSS 0.217f
C22583 RST.n354 VSS 0.00311f
C22584 RST.n355 VSS 0.00116f
C22585 RST.t117 VSS 0.00568f
C22586 RST.t67 VSS 0.00863f
C22587 RST.n356 VSS 0.0152f
C22588 RST.n357 VSS 0.00215f
C22589 RST.n358 VSS 8.37e-19
C22590 RST.n359 VSS 0.00117f
C22591 RST.n360 VSS 0.00409f
C22592 RST.n361 VSS 3.6e-19
C22593 RST.n362 VSS 0.00248f
C22594 RST.n363 VSS 0.00248f
C22595 RST.n364 VSS 1.78f
C22596 RST.n365 VSS 9.22f
C22597 RST.n366 VSS 1.93f
C22598 RST.n367 VSS 0.0921f
C22599 RST.n368 VSS 0.0044f
C22600 RST.t3 VSS 0.00863f
C22601 RST.t9 VSS 0.00568f
C22602 RST.n369 VSS 0.0152f
C22603 RST.n370 VSS 0.00196f
C22604 RST.n371 VSS 7.15e-19
C22605 RST.n372 VSS 5.92e-19
C22606 RST.n373 VSS 5.13e-19
C22607 RST.n374 VSS 6.77e-19
C22608 RST.n375 VSS 0.0034f
C22609 RST.n376 VSS 0.00446f
C22610 RST.t76 VSS 0.00863f
C22611 RST.t99 VSS 0.00568f
C22612 RST.n377 VSS 0.0152f
C22613 RST.n378 VSS 0.00196f
C22614 RST.n379 VSS 7.15e-19
C22615 RST.n380 VSS 7.03e-19
C22616 RST.n381 VSS 6.77e-19
C22617 RST.n382 VSS 0.00344f
C22618 RST.t47 VSS 0.00872f
C22619 RST.t64 VSS 0.00552f
C22620 RST.n383 VSS 0.0153f
C22621 RST.n384 VSS 0.00823f
C22622 RST.t121 VSS 0.00863f
C22623 RST.t61 VSS 0.00568f
C22624 RST.n385 VSS 0.0153f
C22625 RST.n386 VSS 0.00793f
C22626 RST.n387 VSS 0.218f
C22627 RST.n388 VSS 0.216f
C22628 RST.n389 VSS 0.228f
C22629 RST.t56 VSS 0.00568f
C22630 RST.t68 VSS 0.00863f
C22631 RST.n390 VSS 0.0153f
C22632 RST.n391 VSS 0.00779f
C22633 RST.n392 VSS 0.123f
C22634 RST.n393 VSS 7.03e-19
C22635 RST.n394 VSS 6.62e-19
C22636 RST.t12 VSS 0.00542f
C22637 RST.n395 VSS 0.00496f
C22638 RST.n396 VSS 0.00191f
C22639 RST.t21 VSS 0.00861f
C22640 RST.n397 VSS 0.0106f
C22641 RST.n398 VSS 8.34e-20
C22642 RST.n399 VSS 7e-19
C22643 RST.n400 VSS 0.00439f
C22644 RST.n401 VSS 0.00351f
C22645 RST.n402 VSS 0.215f
C22646 RST.t115 VSS 0.00568f
C22647 RST.t124 VSS 0.00863f
C22648 RST.n403 VSS 0.0153f
C22649 RST.n404 VSS 0.00822f
C22650 RST.n405 VSS 0.219f
C22651 RST.t65 VSS 0.00568f
C22652 RST.t78 VSS 0.00863f
C22653 RST.n406 VSS 0.0153f
C22654 RST.n407 VSS 0.00816f
C22655 RST.n408 VSS 1.08f
C22656 RST.n409 VSS 0.0044f
C22657 RST.t52 VSS 0.00863f
C22658 RST.t51 VSS 0.00568f
C22659 RST.n410 VSS 0.0152f
C22660 RST.n411 VSS 0.00196f
C22661 RST.n412 VSS 7.15e-19
C22662 RST.n413 VSS 5.92e-19
C22663 RST.n414 VSS 5.13e-19
C22664 RST.n415 VSS 6.77e-19
C22665 RST.n416 VSS 0.0034f
C22666 RST.n417 VSS 0.00446f
C22667 RST.t40 VSS 0.00863f
C22668 RST.t39 VSS 0.00568f
C22669 RST.n418 VSS 0.0152f
C22670 RST.n419 VSS 0.00196f
C22671 RST.n420 VSS 7.15e-19
C22672 RST.n421 VSS 7.03e-19
C22673 RST.n422 VSS 6.77e-19
C22674 RST.n423 VSS 0.00344f
C22675 RST.t13 VSS 0.00872f
C22676 RST.t11 VSS 0.00552f
C22677 RST.n424 VSS 0.0153f
C22678 RST.n425 VSS 0.00823f
C22679 RST.t103 VSS 0.00863f
C22680 RST.t100 VSS 0.00568f
C22681 RST.n426 VSS 0.0153f
C22682 RST.n427 VSS 0.00793f
C22683 RST.n428 VSS 0.218f
C22684 RST.n429 VSS 0.216f
C22685 RST.n430 VSS 0.228f
C22686 RST.t75 VSS 0.00568f
C22687 RST.t63 VSS 0.00863f
C22688 RST.n431 VSS 0.0153f
C22689 RST.n432 VSS 0.00779f
C22690 RST.n433 VSS 0.123f
C22691 RST.n434 VSS 7.03e-19
C22692 RST.n435 VSS 6.62e-19
C22693 RST.t33 VSS 0.00542f
C22694 RST.n436 VSS 0.00496f
C22695 RST.n437 VSS 0.00191f
C22696 RST.t20 VSS 0.00861f
C22697 RST.n438 VSS 0.0106f
C22698 RST.n439 VSS 8.34e-20
C22699 RST.n440 VSS 7e-19
C22700 RST.n441 VSS 0.00439f
C22701 RST.n442 VSS 0.00351f
C22702 RST.n443 VSS 0.215f
C22703 RST.t38 VSS 0.00568f
C22704 RST.t24 VSS 0.00863f
C22705 RST.n444 VSS 0.0153f
C22706 RST.n445 VSS 0.00822f
C22707 RST.n446 VSS 0.219f
C22708 RST.t84 VSS 0.00568f
C22709 RST.t70 VSS 0.00863f
C22710 RST.n447 VSS 0.0153f
C22711 RST.n448 VSS 0.00816f
C22712 RST.n449 VSS 0.357f
C22713 RST.n450 VSS 7.75f
C22714 RST.n451 VSS 0.821f
C22715 RST.n452 VSS 0.355f
C22716 RST.n453 VSS 0.189f
C22717 RST.n454 VSS 0.0243f
C22718 RST.n455 VSS 7.74f
C22719 RST.n456 VSS 10.8f
C22720 RST.n457 VSS 2.51f
C22721 RST.n458 VSS 0.124f
C22722 RST.n459 VSS 2.82f
C22723 RST.n460 VSS 2.85f
C22724 RST.n461 VSS 0.0452f
C22725 Vdiv.n0 VSS 0.146f
C22726 Vdiv.n1 VSS 0.00333f
C22727 Vdiv.t1 VSS 0.00274f
C22728 Vdiv.n2 VSS 0.00274f
C22729 Vdiv.n3 VSS 0.00757f
C22730 Vdiv.n4 VSS 0.00899f
C22731 VDD.t185 VSS 0.00463f
C22732 VDD.n0 VSS 0.00347f
C22733 VDD.n1 VSS 0.126f
C22734 VDD.t79 VSS 0.0047f
C22735 VDD.n2 VSS 0.133f
C22736 VDD.n3 VSS 0.113f
C22737 VDD.t8 VSS 0.0019f
C22738 VDD.n4 VSS 0.0019f
C22739 VDD.n5 VSS 0.00431f
C22740 VDD.n6 VSS 0.136f
C22741 VDD.n7 VSS 0.124f
C22742 VDD.n8 VSS 0.124f
C22743 VDD.t23 VSS 0.00462f
C22744 VDD.n9 VSS 0.0151f
C22745 VDD.t34 VSS 0.00489f
C22746 VDD.n10 VSS 0.00871f
C22747 VDD.n11 VSS 0.00982f
C22748 VDD.n12 VSS 0.0224f
C22749 VDD.t33 VSS 2.41e-19
C22750 VDD.n13 VSS 0.0944f
C22751 VDD.t9 VSS 0.068f
C22752 VDD.t101 VSS 0.0316f
C22753 VDD.t10 VSS 0.0019f
C22754 VDD.n14 VSS 0.0019f
C22755 VDD.n15 VSS 0.00418f
C22756 VDD.n16 VSS 0.014f
C22757 VDD.n17 VSS 0.00951f
C22758 VDD.n18 VSS 0.0286f
C22759 VDD.t78 VSS 0.0553f
C22760 VDD.n19 VSS 0.0124f
C22761 VDD.t60 VSS 0.00463f
C22762 VDD.n20 VSS 0.0117f
C22763 VDD.n21 VSS 0.00891f
C22764 VDD.n22 VSS 0.00603f
C22765 VDD.n23 VSS 0.0543f
C22766 VDD.t59 VSS 0.0488f
C22767 VDD.t7 VSS 0.0679f
C22768 VDD.t83 VSS 0.0316f
C22769 VDD.t44 VSS 0.00463f
C22770 VDD.n24 VSS 0.0181f
C22771 VDD.n25 VSS 0.00951f
C22772 VDD.n26 VSS 0.0286f
C22773 VDD.t43 VSS 0.0553f
C22774 VDD.t16 VSS 0.00466f
C22775 VDD.n27 VSS 0.0225f
C22776 VDD.n28 VSS 0.00892f
C22777 VDD.n29 VSS 0.0543f
C22778 VDD.t15 VSS 0.0488f
C22779 VDD.t13 VSS 0.0679f
C22780 VDD.t95 VSS 0.0316f
C22781 VDD.t14 VSS 0.0019f
C22782 VDD.n30 VSS 0.0019f
C22783 VDD.n31 VSS 0.00417f
C22784 VDD.n32 VSS 0.0161f
C22785 VDD.n33 VSS 0.00951f
C22786 VDD.n34 VSS 0.0286f
C22787 VDD.t22 VSS 0.0553f
C22788 VDD.n35 VSS 0.0543f
C22789 VDD.t27 VSS 0.00464f
C22790 VDD.t12 VSS 0.0019f
C22791 VDD.n36 VSS 0.0019f
C22792 VDD.n37 VSS 0.00415f
C22793 VDD.t26 VSS 0.0488f
C22794 VDD.t11 VSS 0.0679f
C22795 VDD.t47 VSS 0.0316f
C22796 VDD.n38 VSS 0.0286f
C22797 VDD.t21 VSS 0.00462f
C22798 VDD.t20 VSS 0.0553f
C22799 VDD.t71 VSS 0.0486f
C22800 VDD.n39 VSS 0.0543f
C22801 VDD.t72 VSS 0.00481f
C22802 VDD.n40 VSS 0.0288f
C22803 VDD.n41 VSS 0.0241f
C22804 VDD.n42 VSS 0.00951f
C22805 VDD.n43 VSS 0.0262f
C22806 VDD.n44 VSS 0.0262f
C22807 VDD.n45 VSS 0.00892f
C22808 VDD.n46 VSS 0.178f
C22809 VDD.n47 VSS 2.57f
C22810 VDD.n48 VSS 0.37f
C22811 VDD.n49 VSS 0.493f
C22812 VDD.n50 VSS 0.445f
C22813 VDD.n51 VSS 0.449f
C22814 VDD.n52 VSS 2.99f
C22815 VDD.n53 VSS 0.202f
C22816 VDD.t184 VSS 0.0823f
C22817 VDD.n54 VSS 0.0308f
C22818 VDD.n55 VSS 0.00307f
C22819 VDD.n56 VSS 0.023f
C22820 VDD.n57 VSS 0.0125f
C22821 VDD.t58 VSS 0.00463f
C22822 VDD.t170 VSS 0.0019f
C22823 VDD.n58 VSS 0.0019f
C22824 VDD.n59 VSS 0.00415f
C22825 VDD.n60 VSS 0.0506f
C22826 VDD.t57 VSS 0.0508f
C22827 VDD.t169 VSS 0.0679f
C22828 VDD.t98 VSS 0.0316f
C22829 VDD.n61 VSS 0.0286f
C22830 VDD.t77 VSS 0.00462f
C22831 VDD.n62 VSS 0.0165f
C22832 VDD.n63 VSS 0.00463f
C22833 VDD.t123 VSS 0.0601f
C22834 VDD.n64 VSS 0.0286f
C22835 VDD.t149 VSS 0.00379f
C22836 VDD.n65 VSS 0.0321f
C22837 VDD.n66 VSS 0.00461f
C22838 VDD.t148 VSS 0.0555f
C22839 VDD.t73 VSS 0.0608f
C22840 VDD.n67 VSS 0.0286f
C22841 VDD.t146 VSS 0.00462f
C22842 VDD.n68 VSS 0.00461f
C22843 VDD.t145 VSS 0.0554f
C22844 VDD.t0 VSS 0.0607f
C22845 VDD.n69 VSS 0.0286f
C22846 VDD.t4 VSS 0.00379f
C22847 VDD.n70 VSS 0.0322f
C22848 VDD.n71 VSS 0.00461f
C22849 VDD.t3 VSS 0.0555f
C22850 VDD.t104 VSS 0.0608f
C22851 VDD.n72 VSS 0.0286f
C22852 VDD.t154 VSS 0.00462f
C22853 VDD.n73 VSS 0.00461f
C22854 VDD.t153 VSS 0.0555f
C22855 VDD.t150 VSS 0.0608f
C22856 VDD.n74 VSS 0.0286f
C22857 VDD.t144 VSS 0.00379f
C22858 VDD.n75 VSS 0.0322f
C22859 VDD.n76 VSS 0.00461f
C22860 VDD.t143 VSS 0.0555f
C22861 VDD.t181 VSS 0.0608f
C22862 VDD.n77 VSS 0.0286f
C22863 VDD.t39 VSS 0.00462f
C22864 VDD.n78 VSS 0.00461f
C22865 VDD.t38 VSS 0.0555f
C22866 VDD.t114 VSS 0.0608f
C22867 VDD.n79 VSS 0.0286f
C22868 VDD.t130 VSS 0.00379f
C22869 VDD.n80 VSS 0.0286f
C22870 VDD.t186 VSS 0.0519f
C22871 VDD.t155 VSS 0.12f
C22872 VDD.n81 VSS 0.0573f
C22873 VDD.t112 VSS 0.0629f
C22874 VDD.n82 VSS 0.0496f
C22875 VDD.t65 VSS 0.0518f
C22876 VDD.t66 VSS 0.00481f
C22877 VDD.n84 VSS 0.058f
C22878 VDD.n85 VSS 0.0515f
C22879 VDD.t187 VSS 0.00481f
C22880 VDD.n86 VSS 0.0579f
C22881 VDD.n87 VSS 0.0142f
C22882 VDD.t147 VSS 0.00349f
C22883 VDD.n88 VSS 0.0143f
C22884 VDD.n89 VSS 0.00461f
C22885 VDD.t171 VSS 0.0608f
C22886 VDD.n90 VSS 0.00461f
C22887 VDD.t140 VSS 0.00379f
C22888 VDD.n91 VSS 0.0321f
C22889 VDD.n92 VSS 0.00461f
C22890 VDD.t142 VSS 0.00462f
C22891 VDD.t133 VSS 0.0601f
C22892 VDD.n93 VSS 0.00507f
C22893 VDD.n94 VSS 0.00461f
C22894 VDD.n95 VSS 0.0185f
C22895 VDD.t132 VSS 0.00379f
C22896 VDD.t126 VSS 0.00349f
C22897 VDD.n96 VSS 0.029f
C22898 VDD.n97 VSS 0.00461f
C22899 VDD.n98 VSS 0.00461f
C22900 VDD.t87 VSS 0.00472f
C22901 VDD.t86 VSS 0.0519f
C22902 VDD.t136 VSS 0.0601f
C22903 VDD.n99 VSS 0.00507f
C22904 VDD.t128 VSS 0.00349f
C22905 VDD.n100 VSS 0.0291f
C22906 VDD.n101 VSS 0.0167f
C22907 VDD.n102 VSS 0.0143f
C22908 VDD.n103 VSS 0.0286f
C22909 VDD.t127 VSS 0.0316f
C22910 VDD.n104 VSS 0.0504f
C22911 VDD.n105 VSS 0.0356f
C22912 VDD.n106 VSS 0.0441f
C22913 VDD.n107 VSS 0.0455f
C22914 VDD.n108 VSS 0.0286f
C22915 VDD.t91 VSS 0.00463f
C22916 VDD.t89 VSS 0.00463f
C22917 VDD.t54 VSS 0.12f
C22918 VDD.n109 VSS 0.0573f
C22919 VDD.t52 VSS 0.0629f
C22920 VDD.n110 VSS 0.0496f
C22921 VDD.t90 VSS 0.0518f
C22922 VDD.t88 VSS 0.0519f
C22923 VDD.n112 VSS 0.0515f
C22924 VDD.n113 VSS 0.038f
C22925 VDD.n114 VSS 0.0276f
C22926 VDD.n115 VSS 0.00461f
C22927 VDD.n116 VSS 0.00461f
C22928 VDD.t28 VSS 0.12f
C22929 VDD.n117 VSS 0.0573f
C22930 VDD.t35 VSS 0.00349f
C22931 VDD.n118 VSS 0.029f
C22932 VDD.t32 VSS 0.00349f
C22933 VDD.n119 VSS 0.029f
C22934 VDD.t180 VSS 0.00463f
C22935 VDD.t64 VSS 0.00463f
C22936 VDD.t179 VSS 0.0518f
C22937 VDD.t31 VSS 0.0629f
C22938 VDD.n120 VSS 0.0496f
C22939 VDD.t63 VSS 0.0519f
C22940 VDD.n122 VSS 0.0515f
C22941 VDD.n123 VSS 0.038f
C22942 VDD.n124 VSS 0.0218f
C22943 VDD.n125 VSS 0.00461f
C22944 VDD.n126 VSS 0.00461f
C22945 VDD.n127 VSS 0.0366f
C22946 VDD.n128 VSS 0.0512f
C22947 VDD.n129 VSS 0.0218f
C22948 VDD.n130 VSS 0.0381f
C22949 VDD.n131 VSS 0.0142f
C22950 VDD.n132 VSS 0.0195f
C22951 VDD.n133 VSS 0.0286f
C22952 VDD.n134 VSS 0.0356f
C22953 VDD.n135 VSS 0.0456f
C22954 VDD.n136 VSS 0.0221f
C22955 VDD.n137 VSS 0.0381f
C22956 VDD.n138 VSS 0.0136f
C22957 VDD.n139 VSS 0.02f
C22958 VDD.t53 VSS 0.00349f
C22959 VDD.n140 VSS 0.029f
C22960 VDD.n141 VSS 0.0322f
C22961 VDD.n142 VSS 0.0113f
C22962 VDD.n143 VSS 0.0143f
C22963 VDD.n144 VSS 0.0286f
C22964 VDD.t131 VSS 0.0555f
C22965 VDD.t107 VSS 0.0608f
C22966 VDD.t188 VSS 0.0608f
C22967 VDD.t141 VSS 0.0555f
C22968 VDD.n145 VSS 0.0286f
C22969 VDD.n146 VSS 0.0143f
C22970 VDD.n147 VSS 0.0212f
C22971 VDD.n148 VSS 0.0228f
C22972 VDD.t139 VSS 0.0555f
C22973 VDD.n149 VSS 0.0286f
C22974 VDD.n150 VSS 0.0143f
C22975 VDD.n151 VSS 0.0113f
C22976 VDD.n152 VSS 0.0185f
C22977 VDD.t163 VSS 0.00462f
C22978 VDD.n153 VSS 0.00461f
C22979 VDD.n154 VSS 0.0228f
C22980 VDD.n155 VSS 0.0211f
C22981 VDD.n156 VSS 0.00951f
C22982 VDD.n157 VSS 0.0286f
C22983 VDD.t162 VSS 0.0555f
C22984 VDD.t40 VSS 0.0608f
C22985 VDD.n158 VSS 0.0286f
C22986 VDD.t119 VSS 0.0555f
C22987 VDD.t176 VSS 0.0608f
C22988 VDD.t160 VSS 0.0555f
C22989 VDD.n159 VSS 0.0286f
C22990 VDD.t161 VSS 0.00495f
C22991 VDD.n160 VSS 0.0354f
C22992 VDD.n161 VSS 0.0185f
C22993 VDD.n162 VSS 0.0113f
C22994 VDD.t120 VSS 0.00379f
C22995 VDD.n163 VSS 0.0322f
C22996 VDD.n164 VSS 0.029f
C22997 VDD.n165 VSS 0.0195f
C22998 VDD.t113 VSS 0.00349f
C22999 VDD.n166 VSS 0.029f
C23000 VDD.n167 VSS 0.0322f
C23001 VDD.n168 VSS 0.00461f
C23002 VDD.t129 VSS 0.0555f
C23003 VDD.t166 VSS 0.0608f
C23004 VDD.t164 VSS 0.0555f
C23005 VDD.n169 VSS 0.0286f
C23006 VDD.t165 VSS 0.00495f
C23007 VDD.n170 VSS 0.0354f
C23008 VDD.n171 VSS 0.0185f
C23009 VDD.n172 VSS 0.0113f
C23010 VDD.n173 VSS 0.0143f
C23011 VDD.n174 VSS 0.0228f
C23012 VDD.n175 VSS 0.0211f
C23013 VDD.n176 VSS 0.00951f
C23014 VDD.n177 VSS 0.0185f
C23015 VDD.n178 VSS 0.0113f
C23016 VDD.n179 VSS 0.0143f
C23017 VDD.n180 VSS 0.0228f
C23018 VDD.n181 VSS 0.0212f
C23019 VDD.n182 VSS 0.0143f
C23020 VDD.n183 VSS 0.0185f
C23021 VDD.n184 VSS 0.0113f
C23022 VDD.n185 VSS 0.0143f
C23023 VDD.n186 VSS 0.0228f
C23024 VDD.n187 VSS 0.0211f
C23025 VDD.n188 VSS 0.0143f
C23026 VDD.n189 VSS 0.0185f
C23027 VDD.n190 VSS 0.0118f
C23028 VDD.t76 VSS 0.0443f
C23029 VDD.n191 VSS 0.0483f
C23030 VDD.n192 VSS 0.00432f
C23031 VDD.n193 VSS 0.0165f
C23032 VDD.n194 VSS 0.00227f
C23033 VDD.t36 VSS 0.00161f
C23034 VDD.n195 VSS 0.0111f
C23035 VDD.n196 VSS 0.00227f
C23036 VDD.n197 VSS 0.00177f
C23037 VDD.t37 VSS 0.00463f
C23038 VDD.t175 VSS 0.0019f
C23039 VDD.n198 VSS 0.0019f
C23040 VDD.n199 VSS 0.00415f
C23041 VDD.n200 VSS 0.0242f
C23042 VDD.n201 VSS 0.00951f
C23043 VDD.t46 VSS 0.00462f
C23044 VDD.n202 VSS 0.0241f
C23045 VDD.n203 VSS 0.00892f
C23046 VDD.t62 VSS 0.0019f
C23047 VDD.n204 VSS 0.0019f
C23048 VDD.n205 VSS 0.00415f
C23049 VDD.t118 VSS 0.00463f
C23050 VDD.n206 VSS 0.0258f
C23051 VDD.n207 VSS 0.0262f
C23052 VDD.n208 VSS 0.00951f
C23053 VDD.t25 VSS 0.00462f
C23054 VDD.n209 VSS 0.0241f
C23055 VDD.n210 VSS 0.00892f
C23056 VDD.t68 VSS 0.0019f
C23057 VDD.n211 VSS 0.0019f
C23058 VDD.n212 VSS 0.00415f
C23059 VDD.t6 VSS 0.00463f
C23060 VDD.n213 VSS 0.0258f
C23061 VDD.n214 VSS 0.0262f
C23062 VDD.n215 VSS 0.00951f
C23063 VDD.t110 VSS 0.0447f
C23064 VDD.t51 VSS 0.00462f
C23065 VDD.n216 VSS 0.0241f
C23066 VDD.t111 VSS 0.00481f
C23067 VDD.n217 VSS 0.0288f
C23068 VDD.n218 VSS 0.0543f
C23069 VDD.t50 VSS 0.0553f
C23070 VDD.n219 VSS 0.0286f
C23071 VDD.t17 VSS 0.0316f
C23072 VDD.t67 VSS 0.0679f
C23073 VDD.t5 VSS 0.0447f
C23074 VDD.n220 VSS 0.0543f
C23075 VDD.t24 VSS 0.0553f
C23076 VDD.n221 VSS 0.0286f
C23077 VDD.t92 VSS 0.0316f
C23078 VDD.t61 VSS 0.0679f
C23079 VDD.t117 VSS 0.0447f
C23080 VDD.n222 VSS 0.0543f
C23081 VDD.t45 VSS 0.0553f
C23082 VDD.n223 VSS 0.0286f
C23083 VDD.t80 VSS 0.0316f
C23084 VDD.t174 VSS 0.0514f
C23085 VDD.n224 VSS 0.0431f
C23086 VDD.n225 VSS 0.00284f
C23087 VDD.n226 VSS 0.0146f
C23088 VDD.n227 VSS 0.0115f
C23089 VDD.n228 VSS 0.159f
C23090 VDD.n229 VSS 0.127f
C23091 VDD.n230 VSS 0.00953f
C23092 VDD.n231 VSS 0.0143f
C23093 VDD.n232 VSS 0.161f
C23094 VDD.n233 VSS 0.143f
C23095 VDD.n234 VSS 0.00951f
C23096 VDD.n235 VSS 0.0262f
C23097 VDD.n236 VSS 0.0258f
C23098 VDD.n237 VSS 0.00307f
C23099 VDD90.t453 VSS 0.00244f
C23100 VDD90.n0 VSS 0.00244f
C23101 VDD90.n1 VSS 0.00544f
C23102 VDD90.n2 VSS 0.105f
C23103 VDD90.t379 VSS 0.15f
C23104 VDD90.t408 VSS 0.048f
C23105 VDD90.n3 VSS 0.0557f
C23106 VDD90.t397 VSS 0.023f
C23107 VDD90.t139 VSS 0.006f
C23108 VDD90.n4 VSS 0.11f
C23109 VDD90.n5 VSS 0.0857f
C23110 VDD90.n6 VSS 0.00593f
C23111 VDD90.t454 VSS 0.0714f
C23112 VDD90.n7 VSS 0.0368f
C23113 VDD90.t175 VSS 0.00592f
C23114 VDD90.n8 VSS 0.0059f
C23115 VDD90.n9 VSS 0.0142f
C23116 VDD90.n10 VSS 0.0576f
C23117 VDD90.t174 VSS 0.0465f
C23118 VDD90.t146 VSS 0.0534f
C23119 VDD90.n11 VSS 0.0429f
C23120 VDD90.t37 VSS 0.0526f
C23121 VDD90.n12 VSS 0.0059f
C23122 VDD90.n13 VSS 0.174f
C23123 VDD90.n14 VSS 0.014f
C23124 VDD90.t71 VSS 0.00593f
C23125 VDD90.n15 VSS 0.164f
C23126 VDD90.t42 VSS 0.0273f
C23127 VDD90.n16 VSS 0.00592f
C23128 VDD90.t48 VSS 0.00593f
C23129 VDD90.n17 VSS 0.00592f
C23130 VDD90.n18 VSS 0.0293f
C23131 VDD90.t87 VSS 0.0622f
C23132 VDD90.n19 VSS 0.00592f
C23133 VDD90.t352 VSS 0.0059f
C23134 VDD90.t468 VSS 0.00593f
C23135 VDD90.n20 VSS 0.028f
C23136 VDD90.t351 VSS 0.0523f
C23137 VDD90.t348 VSS 0.0405f
C23138 VDD90.t229 VSS 0.00244f
C23139 VDD90.n21 VSS 0.00244f
C23140 VDD90.n22 VSS 0.00532f
C23141 VDD90.t470 VSS 0.00593f
C23142 VDD90.n23 VSS 0.00592f
C23143 VDD90.n24 VSS 0.0293f
C23144 VDD90.t211 VSS 0.0782f
C23145 VDD90.n25 VSS 0.00592f
C23146 VDD90.t395 VSS 0.00593f
C23147 VDD90.n26 VSS 0.00592f
C23148 VDD90.n27 VSS 0.00592f
C23149 VDD90.t380 VSS 0.0771f
C23150 VDD90.n28 VSS 0.0368f
C23151 VDD90.t438 VSS 0.00593f
C23152 VDD90.n29 VSS 0.00592f
C23153 VDD90.t437 VSS 0.0714f
C23154 VDD90.t214 VSS 0.0782f
C23155 VDD90.n30 VSS 0.0368f
C23156 VDD90.t127 VSS 0.00593f
C23157 VDD90.t132 VSS 0.00244f
C23158 VDD90.n31 VSS 0.00244f
C23159 VDD90.n32 VSS 0.00532f
C23160 VDD90.t126 VSS 0.0714f
C23161 VDD90.t131 VSS 0.0872f
C23162 VDD90.t203 VSS 0.0405f
C23163 VDD90.n33 VSS 0.0368f
C23164 VDD90.t183 VSS 0.00593f
C23165 VDD90.t384 VSS 0.00244f
C23166 VDD90.n34 VSS 0.00244f
C23167 VDD90.n35 VSS 0.00532f
C23168 VDD90.t182 VSS 0.0714f
C23169 VDD90.t383 VSS 0.0872f
C23170 VDD90.t353 VSS 0.0405f
C23171 VDD90.t50 VSS 0.0712f
C23172 VDD90.n36 VSS 0.0368f
C23173 VDD90.t51 VSS 0.00553f
C23174 VDD90.t49 VSS 0.00508f
C23175 VDD90.t472 VSS 0.00385f
C23176 VDD90.n37 VSS 0.00993f
C23177 VDD90.n38 VSS 0.00176f
C23178 VDD90.t66 VSS 0.00508f
C23179 VDD90.t478 VSS 0.00385f
C23180 VDD90.n39 VSS 0.00993f
C23181 VDD90.n40 VSS 0.00233f
C23182 VDD90.n41 VSS 0.00121f
C23183 VDD90.n42 VSS 6.09e-19
C23184 VDD90.n43 VSS 0.00543f
C23185 VDD90.n44 VSS 5.86e-19
C23186 VDD90.t63 VSS 0.00494f
C23187 VDD90.n45 VSS 0.00487f
C23188 VDD90.t481 VSS 0.00384f
C23189 VDD90.n46 VSS 0.00165f
C23190 VDD90.n47 VSS 0.00521f
C23191 VDD90.n48 VSS 0.00179f
C23192 VDD90.n49 VSS 0.00148f
C23193 VDD90.t56 VSS 0.00505f
C23194 VDD90.t484 VSS 0.00386f
C23195 VDD90.n50 VSS 0.00996f
C23196 VDD90.n51 VSS 0.00187f
C23197 VDD90.n52 VSS 0.00158f
C23198 VDD90.n53 VSS 6.09e-19
C23199 VDD90.n54 VSS 0.0192f
C23200 VDD90.n55 VSS 0.0744f
C23201 VDD90.n56 VSS 0.109f
C23202 VDD90.t476 VSS 0.00393f
C23203 VDD90.t72 VSS 0.00499f
C23204 VDD90.n57 VSS 0.00994f
C23205 VDD90.n58 VSS 0.00362f
C23206 VDD90.n59 VSS 0.00148f
C23207 VDD90.t477 VSS 0.00386f
C23208 VDD90.t69 VSS 0.00505f
C23209 VDD90.n60 VSS 0.00996f
C23210 VDD90.n61 VSS 0.00194f
C23211 VDD90.n62 VSS 0.00153f
C23212 VDD90.n63 VSS 6.09e-19
C23213 VDD90.n64 VSS 0.0192f
C23214 VDD90.n65 VSS 0.0251f
C23215 VDD90.n66 VSS 0.121f
C23216 VDD90.n67 VSS 0.0507f
C23217 VDD90.n68 VSS 5.75e-19
C23218 VDD90.n69 VSS 0.00476f
C23219 VDD90.n70 VSS 0.0138f
C23220 VDD90.n71 VSS 0.0338f
C23221 VDD90.n72 VSS 0.0337f
C23222 VDD90.n73 VSS 0.0346f
C23223 VDD90.n74 VSS 0.0184f
C23224 VDD90.n75 VSS 0.0337f
C23225 VDD90.n76 VSS 0.0345f
C23226 VDD90.n77 VSS 0.0205f
C23227 VDD90.n78 VSS 0.0293f
C23228 VDD90.n79 VSS 0.0273f
C23229 VDD90.n80 VSS 0.0205f
C23230 VDD90.n81 VSS 0.0559f
C23231 VDD90.n82 VSS 0.0635f
C23232 VDD90.t232 VSS 0.0771f
C23233 VDD90.t394 VSS 0.0714f
C23234 VDD90.n83 VSS 0.0368f
C23235 VDD90.n84 VSS 0.0205f
C23236 VDD90.n85 VSS 0.0273f
C23237 VDD90.n86 VSS 0.0293f
C23238 VDD90.t134 VSS 0.00593f
C23239 VDD90.n87 VSS 0.0273f
C23240 VDD90.n88 VSS 0.0205f
C23241 VDD90.n89 VSS 0.0368f
C23242 VDD90.t133 VSS 0.0714f
C23243 VDD90.t128 VSS 0.0782f
C23244 VDD90.t228 VSS 0.0872f
C23245 VDD90.t469 VSS 0.0714f
C23246 VDD90.n90 VSS 0.0368f
C23247 VDD90.n91 VSS 0.0205f
C23248 VDD90.n92 VSS 0.0258f
C23249 VDD90.n93 VSS 0.0242f
C23250 VDD90.n94 VSS 0.0184f
C23251 VDD90.n95 VSS 0.0368f
C23252 VDD90.t467 VSS 0.0405f
C23253 VDD90.n96 VSS 0.055f
C23254 VDD90.n97 VSS 0.0186f
C23255 VDD90.n98 VSS 0.00592f
C23256 VDD90.t295 VSS 0.0771f
C23257 VDD90.n99 VSS 0.0368f
C23258 VDD90.t410 VSS 0.00593f
C23259 VDD90.n100 VSS 0.00592f
C23260 VDD90.t409 VSS 0.0714f
C23261 VDD90.t95 VSS 0.0782f
C23262 VDD90.n101 VSS 0.0368f
C23263 VDD90.t41 VSS 0.00593f
C23264 VDD90.t46 VSS 0.00244f
C23265 VDD90.n102 VSS 0.00244f
C23266 VDD90.n103 VSS 0.00532f
C23267 VDD90.t40 VSS 0.0714f
C23268 VDD90.t45 VSS 0.0872f
C23269 VDD90.t225 VSS 0.0405f
C23270 VDD90.n104 VSS 0.0368f
C23271 VDD90.t344 VSS 0.00593f
C23272 VDD90.t298 VSS 0.00244f
C23273 VDD90.n105 VSS 0.00244f
C23274 VDD90.n106 VSS 0.00532f
C23275 VDD90.t343 VSS 0.0714f
C23276 VDD90.t297 VSS 0.0872f
C23277 VDD90.t429 VSS 0.0405f
C23278 VDD90.t73 VSS 0.0712f
C23279 VDD90.n107 VSS 0.0368f
C23280 VDD90.t74 VSS 0.00635f
C23281 VDD90.n108 VSS 0.0456f
C23282 VDD90.n109 VSS 0.0337f
C23283 VDD90.n110 VSS 0.0346f
C23284 VDD90.n111 VSS 0.0184f
C23285 VDD90.n112 VSS 0.0337f
C23286 VDD90.n113 VSS 0.0345f
C23287 VDD90.n114 VSS 0.0205f
C23288 VDD90.n115 VSS 0.0293f
C23289 VDD90.n116 VSS 0.0273f
C23290 VDD90.n117 VSS 0.0205f
C23291 VDD90.n118 VSS 0.0525f
C23292 VDD90.n119 VSS 0.0419f
C23293 VDD90.n120 VSS 0.03f
C23294 VDD90.t99 VSS 0.00593f
C23295 VDD90.n121 VSS 0.0273f
C23296 VDD90.n122 VSS 0.0205f
C23297 VDD90.n123 VSS 0.0317f
C23298 VDD90.t98 VSS 0.0568f
C23299 VDD90.t92 VSS 0.0622f
C23300 VDD90.t47 VSS 0.0421f
C23301 VDD90.n124 VSS 0.0317f
C23302 VDD90.n125 VSS 0.0205f
C23303 VDD90.n126 VSS 0.0273f
C23304 VDD90.n127 VSS 0.0293f
C23305 VDD90.t91 VSS 0.00593f
C23306 VDD90.t86 VSS 0.00244f
C23307 VDD90.n128 VSS 0.00244f
C23308 VDD90.n129 VSS 0.00532f
C23309 VDD90.n130 VSS 0.0242f
C23310 VDD90.t433 VSS 0.00593f
C23311 VDD90.n131 VSS 0.00592f
C23312 VDD90.n132 VSS 0.0291f
C23313 VDD90.t293 VSS 0.0405f
C23314 VDD90.t294 VSS 0.00593f
C23315 VDD90.n133 VSS 0.00592f
C23316 VDD90.n134 VSS 0.0291f
C23317 VDD90.t362 VSS 0.0405f
C23318 VDD90.t363 VSS 0.00593f
C23319 VDD90.n135 VSS 0.00592f
C23320 VDD90.n136 VSS 0.0291f
C23321 VDD90.t115 VSS 0.0059f
C23322 VDD90.n137 VSS 0.0209f
C23323 VDD90.t396 VSS 0.153f
C23324 VDD90.n138 VSS 0.0718f
C23325 VDD90.t83 VSS 0.0757f
C23326 VDD90.t84 VSS 0.0059f
C23327 VDD90.n139 VSS 0.028f
C23328 VDD90.t117 VSS 0.00601f
C23329 VDD90.n140 VSS 0.0322f
C23330 VDD90.n141 VSS 0.0195f
C23331 VDD90.n142 VSS 0.0835f
C23332 VDD90.t116 VSS 0.0493f
C23333 VDD90.t114 VSS 0.0837f
C23334 VDD90.n143 VSS 0.0546f
C23335 VDD90.t303 VSS 0.0467f
C23336 VDD90.n144 VSS 0.0368f
C23337 VDD90.n145 VSS 0.0207f
C23338 VDD90.n146 VSS 0.0276f
C23339 VDD90.t193 VSS 0.0059f
C23340 VDD90.n147 VSS 0.0209f
C23341 VDD90.t192 VSS 0.0525f
C23342 VDD90.n148 VSS 0.0861f
C23343 VDD90.t434 VSS 0.0467f
C23344 VDD90.n149 VSS 0.0368f
C23345 VDD90.n150 VSS 0.0207f
C23346 VDD90.n151 VSS 0.0276f
C23347 VDD90.t407 VSS 0.0059f
C23348 VDD90.n152 VSS 0.0209f
C23349 VDD90.t406 VSS 0.0525f
C23350 VDD90.n153 VSS 0.0861f
C23351 VDD90.t300 VSS 0.0467f
C23352 VDD90.t432 VSS 0.0712f
C23353 VDD90.n154 VSS 0.0368f
C23354 VDD90.n155 VSS 0.0207f
C23355 VDD90.n156 VSS 0.0746f
C23356 VDD90.n157 VSS 0.0627f
C23357 VDD90.n158 VSS 0.0194f
C23358 VDD90.n159 VSS 0.0205f
C23359 VDD90.n160 VSS 0.0317f
C23360 VDD90.t90 VSS 0.0568f
C23361 VDD90.t85 VSS 0.0694f
C23362 VDD90.t422 VSS 0.0322f
C23363 VDD90.n161 VSS 0.0317f
C23364 VDD90.t70 VSS 0.0322f
C23365 VDD90.n162 VSS 0.0908f
C23366 VDD90.t427 VSS 0.0653f
C23367 VDD90.t428 VSS 0.0059f
C23368 VDD90.t32 VSS 0.0622f
C23369 VDD90.n163 VSS 0.0317f
C23370 VDD90.t12 VSS 0.00593f
C23371 VDD90.n164 VSS 0.00592f
C23372 VDD90.t11 VSS 0.0568f
C23373 VDD90.t24 VSS 0.0622f
C23374 VDD90.n165 VSS 0.0317f
C23375 VDD90.n166 VSS 0.124f
C23376 VDD90.t317 VSS 0.00593f
C23377 VDD90.n167 VSS 0.00592f
C23378 VDD90.n168 VSS 0.0317f
C23379 VDD90.n169 VSS 0.137f
C23380 VDD90.n170 VSS 0.00601f
C23381 VDD90.n171 VSS 0.108f
C23382 VDD90.n172 VSS 0.0846f
C23383 VDD90.n173 VSS 0.00592f
C23384 VDD90.n174 VSS 0.00592f
C23385 VDD90.t356 VSS 0.0771f
C23386 VDD90.n175 VSS 0.0368f
C23387 VDD90.t418 VSS 0.00593f
C23388 VDD90.n176 VSS 0.00592f
C23389 VDD90.t417 VSS 0.0714f
C23390 VDD90.t414 VSS 0.0782f
C23391 VDD90.n177 VSS 0.0368f
C23392 VDD90.t188 VSS 0.00593f
C23393 VDD90.t197 VSS 0.00244f
C23394 VDD90.n178 VSS 0.00244f
C23395 VDD90.n179 VSS 0.00532f
C23396 VDD90.t187 VSS 0.0714f
C23397 VDD90.t196 VSS 0.0872f
C23398 VDD90.t272 VSS 0.0405f
C23399 VDD90.n180 VSS 0.0368f
C23400 VDD90.t218 VSS 0.00593f
C23401 VDD90.t365 VSS 0.00244f
C23402 VDD90.n181 VSS 0.00244f
C23403 VDD90.n182 VSS 0.00532f
C23404 VDD90.t217 VSS 0.0714f
C23405 VDD90.t364 VSS 0.0872f
C23406 VDD90.t18 VSS 0.0405f
C23407 VDD90.t64 VSS 0.0712f
C23408 VDD90.n183 VSS 0.0368f
C23409 VDD90.t65 VSS 0.00635f
C23410 VDD90.n184 VSS 0.0456f
C23411 VDD90.n185 VSS 0.0337f
C23412 VDD90.n186 VSS 0.0346f
C23413 VDD90.n187 VSS 0.0184f
C23414 VDD90.n188 VSS 0.0337f
C23415 VDD90.n189 VSS 0.0345f
C23416 VDD90.n190 VSS 0.0205f
C23417 VDD90.n191 VSS 0.0293f
C23418 VDD90.n192 VSS 0.0273f
C23419 VDD90.n193 VSS 0.0205f
C23420 VDD90.n194 VSS 0.0525f
C23421 VDD90.t367 VSS 0.0059f
C23422 VDD90.t316 VSS 0.0421f
C23423 VDD90.t320 VSS 0.0273f
C23424 VDD90.n195 VSS 0.164f
C23425 VDD90.t277 VSS 0.0568f
C23426 VDD90.t35 VSS 0.0694f
C23427 VDD90.t359 VSS 0.0322f
C23428 VDD90.t36 VSS 0.00244f
C23429 VDD90.n196 VSS 0.00244f
C23430 VDD90.n197 VSS 0.00532f
C23431 VDD90.n198 VSS 0.0242f
C23432 VDD90.t231 VSS 0.00593f
C23433 VDD90.n199 VSS 0.0193f
C23434 VDD90.n200 VSS 0.0184f
C23435 VDD90.n201 VSS 0.0317f
C23436 VDD90.t230 VSS 0.0322f
C23437 VDD90.n202 VSS 0.0908f
C23438 VDD90.t366 VSS 0.0653f
C23439 VDD90.n203 VSS 0.0182f
C23440 VDD90.n204 VSS 0.0372f
C23441 VDD90.n205 VSS 0.0429f
C23442 VDD90.n206 VSS 0.0753f
C23443 VDD90.n207 VSS 0.00593f
C23444 VDD90.t259 VSS 0.0714f
C23445 VDD90.n208 VSS 0.0368f
C23446 VDD90.t241 VSS 0.00592f
C23447 VDD90.t195 VSS 0.00603f
C23448 VDD90.n209 VSS 0.099f
C23449 VDD90.t240 VSS 0.0465f
C23450 VDD90.t8 VSS 0.0534f
C23451 VDD90.n210 VSS 0.0923f
C23452 VDD90.n211 VSS 0.00743f
C23453 VDD90.n212 VSS 0.0142f
C23454 VDD90.n213 VSS 0.0197f
C23455 VDD90.t202 VSS 0.00603f
C23456 VDD90.n214 VSS 0.00592f
C23457 VDD90.n215 VSS 0.0249f
C23458 VDD90.t184 VSS 0.0273f
C23459 VDD90.t210 VSS 0.00244f
C23460 VDD90.n216 VSS 0.00244f
C23461 VDD90.n217 VSS 0.00532f
C23462 VDD90.n218 VSS 0.0242f
C23463 VDD90.n219 VSS 0.015f
C23464 VDD90.t411 VSS 0.0622f
C23465 VDD90.n220 VSS 0.00592f
C23466 VDD90.t121 VSS 0.00593f
C23467 VDD90.t206 VSS 0.0622f
C23468 VDD90.t120 VSS 0.0568f
C23469 VDD90.n221 VSS 0.0317f
C23470 VDD90.n222 VSS 0.0242f
C23471 VDD90.n223 VSS 0.0251f
C23472 VDD90.n224 VSS 0.0293f
C23473 VDD90.n225 VSS 0.0205f
C23474 VDD90.n226 VSS 0.0317f
C23475 VDD90.t194 VSS 0.0421f
C23476 VDD90.n227 VSS 0.164f
C23477 VDD90.n228 VSS 0.0059f
C23478 VDD90.n229 VSS 0.0267f
C23479 VDD90.t158 VSS 0.0504f
C23480 VDD90.t103 VSS 0.0526f
C23481 VDD90.n230 VSS 0.0609f
C23482 VDD90.t439 VSS 0.053f
C23483 VDD90.n231 VSS 0.0358f
C23484 VDD90.n232 VSS 0.0172f
C23485 VDD90.n233 VSS 0.159f
C23486 VDD90.t58 VSS 0.00603f
C23487 VDD90.n234 VSS 0.129f
C23488 VDD90.t17 VSS 0.00618f
C23489 VDD90.t16 VSS 0.0653f
C23490 VDD90.n235 VSS 0.0908f
C23491 VDD90.t57 VSS 0.0322f
C23492 VDD90.n236 VSS 0.0317f
C23493 VDD90.t13 VSS 0.0322f
C23494 VDD90.t209 VSS 0.0694f
C23495 VDD90.t201 VSS 0.0568f
C23496 VDD90.n237 VSS 0.0317f
C23497 VDD90.n238 VSS 0.0205f
C23498 VDD90.n239 VSS 0.0976f
C23499 VDD90.n240 VSS 0.0924f
C23500 VDD90.n241 VSS 0.0347f
C23501 VDD90.n242 VSS 0.0297f
C23502 VDD90.n243 VSS 0.0999f
C23503 VDD90.n244 VSS 0.0351f
C23504 VDD90.n245 VSS 0.029f
C23505 VDD90.n246 VSS 0.0324f
C23506 VDD90.t256 VSS 0.00244f
C23507 VDD90.n247 VSS 0.00244f
C23508 VDD90.n248 VSS 0.00532f
C23509 VDD90.n249 VSS 0.0191f
C23510 VDD90.n250 VSS 0.00593f
C23511 VDD90.n251 VSS 0.0261f
C23512 VDD90.t252 VSS 0.0524f
C23513 VDD90.n252 VSS 0.0059f
C23514 VDD90.t239 VSS 0.00592f
C23515 VDD90.t108 VSS 0.0716f
C23516 VDD90.n253 VSS 0.00593f
C23517 VDD90.t444 VSS 0.00244f
C23518 VDD90.n254 VSS 0.00244f
C23519 VDD90.n255 VSS 0.00532f
C23520 VDD90.n256 VSS 0.00593f
C23521 VDD90.n257 VSS 0.0346f
C23522 VDD90.t76 VSS 0.0714f
C23523 VDD90.n258 VSS 7.98e-19
C23524 VDD90.t480 VSS 0.00385f
C23525 VDD90.n259 VSS 0.00529f
C23526 VDD90.t75 VSS 0.00498f
C23527 VDD90.n260 VSS 0.00474f
C23528 VDD90.t473 VSS 0.00385f
C23529 VDD90.t52 VSS 0.00508f
C23530 VDD90.n261 VSS 0.00992f
C23531 VDD90.n262 VSS 0.066f
C23532 VDD90.n263 VSS 0.0648f
C23533 VDD90.n264 VSS 0.00286f
C23534 VDD90.n265 VSS 0.00553f
C23535 VDD90.n266 VSS 0.0156f
C23536 VDD90.t258 VSS 0.00244f
C23537 VDD90.n267 VSS 0.00244f
C23538 VDD90.n268 VSS 0.00532f
C23539 VDD90.n269 VSS 0.0338f
C23540 VDD90.n270 VSS 0.0338f
C23541 VDD90.n271 VSS 0.0368f
C23542 VDD90.t257 VSS 0.0404f
C23543 VDD90.t242 VSS 0.0872f
C23544 VDD90.t385 VSS 0.0716f
C23545 VDD90.t391 VSS 0.0872f
C23546 VDD90.t443 VSS 0.0404f
C23547 VDD90.n272 VSS 0.0368f
C23548 VDD90.n273 VSS 0.0183f
C23549 VDD90.n274 VSS 0.0338f
C23550 VDD90.n275 VSS 0.0345f
C23551 VDD90.t125 VSS 0.00592f
C23552 VDD90.n276 VSS 0.00593f
C23553 VDD90.n277 VSS 0.0272f
C23554 VDD90.n278 VSS 0.0293f
C23555 VDD90.n279 VSS 0.0205f
C23556 VDD90.n280 VSS 0.0368f
C23557 VDD90.t124 VSS 0.0781f
C23558 VDD90.t111 VSS 0.0716f
C23559 VDD90.t238 VSS 0.077f
C23560 VDD90.n281 VSS 0.0368f
C23561 VDD90.n282 VSS 0.0205f
C23562 VDD90.n283 VSS 0.0524f
C23563 VDD90.t307 VSS 0.00592f
C23564 VDD90.t388 VSS 0.0716f
C23565 VDD90.n284 VSS 0.00593f
C23566 VDD90.t400 VSS 0.0407f
C23567 VDD90.n285 VSS 0.00593f
C23568 VDD90.n286 VSS 0.00618f
C23569 VDD90.t262 VSS 0.0524f
C23570 VDD90.n287 VSS 0.055f
C23571 VDD90.n288 VSS 0.028f
C23572 VDD90.t266 VSS 0.00244f
C23573 VDD90.n289 VSS 0.00244f
C23574 VDD90.n290 VSS 0.00544f
C23575 VDD90.n291 VSS 0.142f
C23576 VDD90.n292 VSS 0.00593f
C23577 VDD90.n293 VSS 0.0258f
C23578 VDD90.n294 VSS 0.105f
C23579 VDD90.n295 VSS 0.0183f
C23580 VDD90.n296 VSS 0.0368f
C23581 VDD90.t265 VSS 0.0404f
C23582 VDD90.t308 VSS 0.0872f
C23583 VDD90.t249 VSS 0.0716f
C23584 VDD90.t106 VSS 0.0781f
C23585 VDD90.n297 VSS 0.0368f
C23586 VDD90.n298 VSS 0.0178f
C23587 VDD90.t107 VSS 0.006f
C23588 VDD90.n299 VSS 0.11f
C23589 VDD90.n300 VSS 0.0182f
C23590 VDD90.t123 VSS 0.00592f
C23591 VDD90.n301 VSS 0.0231f
C23592 VDD90.n302 VSS 0.0205f
C23593 VDD90.n303 VSS 0.0368f
C23594 VDD90.t122 VSS 0.0781f
C23595 VDD90.t340 VSS 0.0716f
C23596 VDD90.t306 VSS 0.077f
C23597 VDD90.n304 VSS 0.0368f
C23598 VDD90.n305 VSS 0.0205f
C23599 VDD90.n306 VSS 0.0301f
C23600 VDD90.n307 VSS 0.0418f
C23601 VDD90.n308 VSS 0.0186f
C23602 VDD90.n309 VSS 0.055f
C23603 VDD90.t235 VSS 0.0407f
C23604 VDD90.t285 VSS 0.0781f
C23605 VDD90.n310 VSS 0.00593f
C23606 VDD90.n311 VSS 0.0258f
C23607 VDD90.t286 VSS 0.00592f
C23608 VDD90.n312 VSS 0.00593f
C23609 VDD90.t287 VSS 0.0716f
C23610 VDD90.n313 VSS 0.0368f
C23611 VDD90.t153 VSS 0.00592f
C23612 VDD90.n314 VSS 0.00593f
C23613 VDD90.t152 VSS 0.0781f
C23614 VDD90.t269 VSS 0.0716f
C23615 VDD90.t398 VSS 0.077f
C23616 VDD90.n315 VSS 0.0368f
C23617 VDD90.t399 VSS 0.00592f
C23618 VDD90.t449 VSS 0.00592f
C23619 VDD90.t282 VSS 0.0716f
C23620 VDD90.n316 VSS 0.00593f
C23621 VDD90.t276 VSS 0.00244f
C23622 VDD90.n317 VSS 0.00244f
C23623 VDD90.n318 VSS 0.00532f
C23624 VDD90.n319 VSS 0.00593f
C23625 VDD90.n320 VSS 0.0346f
C23626 VDD90.t53 VSS 0.0714f
C23627 VDD90.n321 VSS 0.00635f
C23628 VDD90.t268 VSS 0.00244f
C23629 VDD90.n322 VSS 0.00244f
C23630 VDD90.n323 VSS 0.00532f
C23631 VDD90.n324 VSS 0.0338f
C23632 VDD90.n325 VSS 0.0456f
C23633 VDD90.n326 VSS 0.0368f
C23634 VDD90.t267 VSS 0.0404f
C23635 VDD90.t445 VSS 0.0872f
C23636 VDD90.t149 VSS 0.0716f
C23637 VDD90.t290 VSS 0.0872f
C23638 VDD90.t275 VSS 0.0404f
C23639 VDD90.n327 VSS 0.0368f
C23640 VDD90.n328 VSS 0.0183f
C23641 VDD90.n329 VSS 0.0338f
C23642 VDD90.n330 VSS 0.0345f
C23643 VDD90.t155 VSS 0.00592f
C23644 VDD90.n331 VSS 0.00593f
C23645 VDD90.n332 VSS 0.0272f
C23646 VDD90.n333 VSS 0.0293f
C23647 VDD90.n334 VSS 0.0205f
C23648 VDD90.n335 VSS 0.0368f
C23649 VDD90.t154 VSS 0.0781f
C23650 VDD90.t373 VSS 0.0716f
C23651 VDD90.t448 VSS 0.077f
C23652 VDD90.n336 VSS 0.0368f
C23653 VDD90.n337 VSS 0.0205f
C23654 VDD90.n338 VSS 0.0558f
C23655 VDD90.n339 VSS 0.0634f
C23656 VDD90.n340 VSS 0.0205f
C23657 VDD90.n341 VSS 0.0272f
C23658 VDD90.n342 VSS 0.0293f
C23659 VDD90.n343 VSS 0.0205f
C23660 VDD90.n344 VSS 0.0272f
C23661 VDD90.n345 VSS 0.0293f
C23662 VDD90.n346 VSS 0.0205f
C23663 VDD90.n347 VSS 0.0368f
C23664 VDD90.t27 VSS 0.0716f
C23665 VDD90.t403 VSS 0.0872f
C23666 VDD90.t255 VSS 0.0404f
C23667 VDD90.n348 VSS 0.0368f
C23668 VDD90.n349 VSS 0.0137f
C23669 VDD90.n350 VSS 0.0462f
C23670 VDD90.n351 VSS 0.0524f
C23671 VDD90.n352 VSS 0.0969f
C23672 VDD90.n353 VSS 0.167f
C23673 VDD90.n354 VSS 0.143f
C23674 VDD90.n355 VSS 0.127f
C23675 VDD90.t278 VSS 0.00603f
C23676 VDD90.n356 VSS 0.0976f
C23677 VDD90.n357 VSS 0.0205f
C23678 VDD90.n358 VSS 0.0293f
C23679 VDD90.n359 VSS 0.0265f
C23680 VDD90.n360 VSS 0.0737f
C23681 VDD90.n361 VSS 0.0205f
C23682 VDD90.n362 VSS 0.0293f
C23683 VDD90.n363 VSS 0.0273f
C23684 VDD90.n364 VSS 0.0179f
C23685 VDD90.n365 VSS 0.00602f
C23686 VDD90.n366 VSS 0.102f
C23687 VDD90.n367 VSS 0.00592f
C23688 VDD90.t419 VSS 0.0771f
C23689 VDD90.n368 VSS 0.0368f
C23690 VDD90.t31 VSS 0.00593f
C23691 VDD90.n369 VSS 0.00592f
C23692 VDD90.t30 VSS 0.0714f
C23693 VDD90.t21 VSS 0.0782f
C23694 VDD90.n370 VSS 0.0368f
C23695 VDD90.t319 VSS 0.00593f
C23696 VDD90.t315 VSS 0.00244f
C23697 VDD90.n371 VSS 0.00244f
C23698 VDD90.n372 VSS 0.00532f
C23699 VDD90.t318 VSS 0.0714f
C23700 VDD90.t314 VSS 0.0872f
C23701 VDD90.t440 VSS 0.0405f
C23702 VDD90.n373 VSS 0.0368f
C23703 VDD90.t157 VSS 0.00593f
C23704 VDD90.t426 VSS 0.00244f
C23705 VDD90.n374 VSS 0.00244f
C23706 VDD90.n375 VSS 0.00532f
C23707 VDD90.t156 VSS 0.0714f
C23708 VDD90.t425 VSS 0.0872f
C23709 VDD90.t345 VSS 0.0405f
C23710 VDD90.t67 VSS 0.0712f
C23711 VDD90.n376 VSS 0.0368f
C23712 VDD90.t68 VSS 0.00635f
C23713 VDD90.n377 VSS 0.0456f
C23714 VDD90.n378 VSS 0.0337f
C23715 VDD90.n379 VSS 0.0346f
C23716 VDD90.n380 VSS 0.0184f
C23717 VDD90.n381 VSS 0.0337f
C23718 VDD90.n382 VSS 0.0345f
C23719 VDD90.n383 VSS 0.0205f
C23720 VDD90.n384 VSS 0.0293f
C23721 VDD90.n385 VSS 0.0273f
C23722 VDD90.n386 VSS 0.0205f
C23723 VDD90.n387 VSS 0.0525f
C23724 VDD90.n388 VSS 0.0351f
C23725 VDD90.n389 VSS 0.0186f
C23726 VDD90.n390 VSS 0.0261f
C23727 VDD90.n391 VSS 0.0737f
C23728 VDD90.n392 VSS 0.173f
C23729 VDD90.n393 VSS 0.0727f
C23730 VDD90.n394 VSS 0.0193f
C23731 VDD90.n395 VSS 0.0609f
C23732 VDD90.t219 VSS 0.053f
C23733 VDD90.n396 VSS 0.0358f
C23734 VDD90.t311 VSS 0.0504f
C23735 VDD90.n397 VSS 0.0923f
C23736 VDD90.n398 VSS 0.0399f
C23737 VDD90.n399 VSS 0.047f
C23738 VDD90.n400 VSS 0.029f
C23739 VDD90.n401 VSS 0.0446f
C23740 VDD90.n402 VSS 0.0852f
C23741 VDD90.t170 VSS 0.00592f
C23742 VDD90.t135 VSS 0.0716f
C23743 VDD90.n403 VSS 0.00593f
C23744 VDD90.t248 VSS 0.00244f
C23745 VDD90.n404 VSS 0.00244f
C23746 VDD90.n405 VSS 0.00532f
C23747 VDD90.n406 VSS 0.00593f
C23748 VDD90.n407 VSS 0.0346f
C23749 VDD90.t80 VSS 0.0714f
C23750 VDD90.n408 VSS 5.86e-19
C23751 VDD90.t471 VSS 0.00385f
C23752 VDD90.t59 VSS 0.00508f
C23753 VDD90.n409 VSS 0.00992f
C23754 VDD90.n410 VSS 0.066f
C23755 VDD90.n411 VSS 0.0652f
C23756 VDD90.t479 VSS 0.00385f
C23757 VDD90.t79 VSS 0.00498f
C23758 VDD90.n412 VSS 0.00474f
C23759 VDD90.n413 VSS 0.00529f
C23760 VDD90.n414 VSS 8.37e-19
C23761 VDD90.n415 VSS 0.00442f
C23762 VDD90.n416 VSS 0.00553f
C23763 VDD90.n417 VSS 0.0138f
C23764 VDD90.t451 VSS 0.00244f
C23765 VDD90.n418 VSS 0.00244f
C23766 VDD90.n419 VSS 0.00532f
C23767 VDD90.n420 VSS 0.0338f
C23768 VDD90.n421 VSS 0.0338f
C23769 VDD90.n422 VSS 0.0368f
C23770 VDD90.t450 VSS 0.0404f
C23771 VDD90.t176 VSS 0.0872f
C23772 VDD90.t198 VSS 0.0716f
C23773 VDD90.t337 VSS 0.0872f
C23774 VDD90.t247 VSS 0.0404f
C23775 VDD90.n423 VSS 0.0368f
C23776 VDD90.n424 VSS 0.0183f
C23777 VDD90.n425 VSS 0.0338f
C23778 VDD90.n426 VSS 0.0345f
C23779 VDD90.t3 VSS 0.00592f
C23780 VDD90.n427 VSS 0.00593f
C23781 VDD90.n428 VSS 0.0272f
C23782 VDD90.n429 VSS 0.0293f
C23783 VDD90.n430 VSS 0.0205f
C23784 VDD90.n431 VSS 0.0368f
C23785 VDD90.t2 VSS 0.0781f
C23786 VDD90.t279 VSS 0.0716f
C23787 VDD90.t169 VSS 0.077f
C23788 VDD90.n432 VSS 0.0368f
C23789 VDD90.n433 VSS 0.0205f
C23790 VDD90.n434 VSS 0.0511f
C23791 VDD90.t372 VSS 0.00592f
C23792 VDD90.n435 VSS 0.00593f
C23793 VDD90.n436 VSS 0.0221f
C23794 VDD90.t164 VSS 0.0407f
C23795 VDD90.n437 VSS 0.00593f
C23796 VDD90.n438 VSS 0.00618f
C23797 VDD90.t457 VSS 0.0524f
C23798 VDD90.n439 VSS 0.055f
C23799 VDD90.n440 VSS 0.028f
C23800 VDD90.n441 VSS 0.0183f
C23801 VDD90.n442 VSS 0.0368f
C23802 VDD90.t452 VSS 0.0404f
C23803 VDD90.t368 VSS 0.0872f
C23804 VDD90.t100 VSS 0.0716f
C23805 VDD90.n443 VSS 0.00593f
C23806 VDD90.n444 VSS 0.0258f
C23807 VDD90.n445 VSS 0.0164f
C23808 VDD90.n446 VSS 0.0368f
C23809 VDD90.t138 VSS 0.0781f
C23810 VDD90.t334 VSS 0.0716f
C23811 VDD90.n447 VSS 0.00593f
C23812 VDD90.n448 VSS 0.0196f
C23813 VDD90.t1 VSS 0.00592f
C23814 VDD90.n449 VSS 0.0235f
C23815 VDD90.n450 VSS 0.0205f
C23816 VDD90.n451 VSS 0.0368f
C23817 VDD90.t0 VSS 0.0781f
C23818 VDD90.t189 VSS 0.0716f
C23819 VDD90.t371 VSS 0.077f
C23820 VDD90.n452 VSS 0.0368f
C23821 VDD90.n453 VSS 0.0205f
C23822 VDD90.n454 VSS 0.0286f
C23823 VDD90.n455 VSS 0.0416f
C23824 VDD90.n456 VSS 0.0059f
C23825 VDD90.n457 VSS 0.00593f
C23826 VDD90.n458 VSS 0.0261f
C23827 VDD90.t462 VSS 0.0524f
C23828 VDD90.n459 VSS 0.0137f
C23829 VDD90.t332 VSS 0.0781f
C23830 VDD90.n460 VSS 0.00593f
C23831 VDD90.t461 VSS 0.00244f
C23832 VDD90.n461 VSS 0.00244f
C23833 VDD90.n462 VSS 0.00532f
C23834 VDD90.n463 VSS 0.0462f
C23835 VDD90.n464 VSS 0.0191f
C23836 VDD90.n465 VSS 0.0258f
C23837 VDD90.t333 VSS 0.00592f
C23838 VDD90.n466 VSS 0.00593f
C23839 VDD90.t323 VSS 0.0716f
C23840 VDD90.n467 VSS 0.0368f
C23841 VDD90.t5 VSS 0.00592f
C23842 VDD90.n468 VSS 0.00593f
C23843 VDD90.t4 VSS 0.0781f
C23844 VDD90.t179 VSS 0.0716f
C23845 VDD90.t167 VSS 0.077f
C23846 VDD90.n469 VSS 0.0368f
C23847 VDD90.t168 VSS 0.00592f
C23848 VDD90.t224 VSS 0.00592f
C23849 VDD90.t329 VSS 0.0716f
C23850 VDD90.n470 VSS 0.00593f
C23851 VDD90.t246 VSS 0.00244f
C23852 VDD90.n471 VSS 0.00244f
C23853 VDD90.n472 VSS 0.00532f
C23854 VDD90.n473 VSS 0.00593f
C23855 VDD90.n474 VSS 0.0346f
C23856 VDD90.t60 VSS 0.0714f
C23857 VDD90.n475 VSS 0.00635f
C23858 VDD90.t466 VSS 0.00244f
C23859 VDD90.n476 VSS 0.00244f
C23860 VDD90.n477 VSS 0.00532f
C23861 VDD90.n478 VSS 0.0338f
C23862 VDD90.n479 VSS 0.0456f
C23863 VDD90.n480 VSS 0.0368f
C23864 VDD90.t465 VSS 0.0404f
C23865 VDD90.t220 VSS 0.0872f
C23866 VDD90.t143 VSS 0.0716f
C23867 VDD90.t326 VSS 0.0872f
C23868 VDD90.t245 VSS 0.0404f
C23869 VDD90.n481 VSS 0.0368f
C23870 VDD90.n482 VSS 0.0183f
C23871 VDD90.n483 VSS 0.0338f
C23872 VDD90.n484 VSS 0.0345f
C23873 VDD90.t7 VSS 0.00592f
C23874 VDD90.n485 VSS 0.00593f
C23875 VDD90.n486 VSS 0.0272f
C23876 VDD90.n487 VSS 0.0293f
C23877 VDD90.n488 VSS 0.0205f
C23878 VDD90.n489 VSS 0.0368f
C23879 VDD90.t6 VSS 0.0781f
C23880 VDD90.t140 VSS 0.0716f
C23881 VDD90.t223 VSS 0.077f
C23882 VDD90.n490 VSS 0.0368f
C23883 VDD90.n491 VSS 0.0205f
C23884 VDD90.n492 VSS 0.0558f
C23885 VDD90.n493 VSS 0.0634f
C23886 VDD90.n494 VSS 0.0205f
C23887 VDD90.n495 VSS 0.0272f
C23888 VDD90.n496 VSS 0.0293f
C23889 VDD90.n497 VSS 0.0205f
C23890 VDD90.n498 VSS 0.0272f
C23891 VDD90.n499 VSS 0.0293f
C23892 VDD90.n500 VSS 0.0205f
C23893 VDD90.n501 VSS 0.0368f
C23894 VDD90.t376 VSS 0.0716f
C23895 VDD90.t161 VSS 0.0872f
C23896 VDD90.t460 VSS 0.0404f
C23897 VDD90.n502 VSS 0.0368f
C23898 VDD90.t171 VSS 0.0407f
C23899 VDD90.n503 VSS 0.055f
C23900 VDD90.n504 VSS 0.0188f
C23901 VDD90.n505 VSS 0.0847f
C23902 VDD90.n506 VSS 0.185f
C23903 VDD90.n507 VSS 0.184f
C23904 VDD90.n508 VSS 0.15f
C23905 VDD90.n509 VSS 0.04f
C23906 VDD90.n510 VSS 0.0487f
C23907 VDD90.n511 VSS 0.014f
C23908 VDD90.n512 VSS 0.326f
C23909 VDD90.n513 VSS 0.00163f
C23910 VDD90.n514 VSS 0.00592f
C23911 VDD90.n515 VSS 0.0153f
C23912 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n0 VSS 2.07f
C23913 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t0 VSS 0.0344f
C23914 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n1 VSS 0.0344f
C23915 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n2 VSS 0.0734f
C23916 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t3 VSS 0.0774f
C23917 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t2 VSS 0.0493f
C23918 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n3 VSS 0.137f
C23919 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t7 VSS 0.0552f
C23920 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t5 VSS 0.0708f
C23921 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n4 VSS 0.141f
C23922 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t4 VSS 0.055f
C23923 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.t6 VSS 0.044f
C23924 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n5 VSS 0.131f
C23925 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n6 VSS 1.18f
C23926 CLK_div_90_mag_0.CLK_div_3_mag_0.JK_FF_mag_1.K.n7 VSS 0.215f
.ends

