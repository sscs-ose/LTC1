magic
tech gf180mcuC
magscale 1 10
timestamp 1693883759
<< error_p >>
rect -1303 -48 -1257 48
rect -1143 -48 -1097 48
rect -983 -48 -937 48
rect -823 -48 -777 48
rect -663 -48 -617 48
rect -503 -48 -457 48
rect -343 -48 -297 48
rect -183 -48 -137 48
rect -23 -48 23 48
rect 137 -48 183 48
rect 297 -48 343 48
rect 457 -48 503 48
rect 617 -48 663 48
rect 777 -48 823 48
rect 937 -48 983 48
rect 1097 -48 1143 48
rect 1257 -48 1303 48
<< nwell >>
rect -1402 -180 1402 180
<< pmos >>
rect -1228 -50 -1172 50
rect -1068 -50 -1012 50
rect -908 -50 -852 50
rect -748 -50 -692 50
rect -588 -50 -532 50
rect -428 -50 -372 50
rect -268 -50 -212 50
rect -108 -50 -52 50
rect 52 -50 108 50
rect 212 -50 268 50
rect 372 -50 428 50
rect 532 -50 588 50
rect 692 -50 748 50
rect 852 -50 908 50
rect 1012 -50 1068 50
rect 1172 -50 1228 50
<< pdiff >>
rect -1316 37 -1228 50
rect -1316 -37 -1303 37
rect -1257 -37 -1228 37
rect -1316 -50 -1228 -37
rect -1172 37 -1068 50
rect -1172 -37 -1143 37
rect -1097 -37 -1068 37
rect -1172 -50 -1068 -37
rect -1012 37 -908 50
rect -1012 -37 -983 37
rect -937 -37 -908 37
rect -1012 -50 -908 -37
rect -852 37 -748 50
rect -852 -37 -823 37
rect -777 -37 -748 37
rect -852 -50 -748 -37
rect -692 37 -588 50
rect -692 -37 -663 37
rect -617 -37 -588 37
rect -692 -50 -588 -37
rect -532 37 -428 50
rect -532 -37 -503 37
rect -457 -37 -428 37
rect -532 -50 -428 -37
rect -372 37 -268 50
rect -372 -37 -343 37
rect -297 -37 -268 37
rect -372 -50 -268 -37
rect -212 37 -108 50
rect -212 -37 -183 37
rect -137 -37 -108 37
rect -212 -50 -108 -37
rect -52 37 52 50
rect -52 -37 -23 37
rect 23 -37 52 37
rect -52 -50 52 -37
rect 108 37 212 50
rect 108 -37 137 37
rect 183 -37 212 37
rect 108 -50 212 -37
rect 268 37 372 50
rect 268 -37 297 37
rect 343 -37 372 37
rect 268 -50 372 -37
rect 428 37 532 50
rect 428 -37 457 37
rect 503 -37 532 37
rect 428 -50 532 -37
rect 588 37 692 50
rect 588 -37 617 37
rect 663 -37 692 37
rect 588 -50 692 -37
rect 748 37 852 50
rect 748 -37 777 37
rect 823 -37 852 37
rect 748 -50 852 -37
rect 908 37 1012 50
rect 908 -37 937 37
rect 983 -37 1012 37
rect 908 -50 1012 -37
rect 1068 37 1172 50
rect 1068 -37 1097 37
rect 1143 -37 1172 37
rect 1068 -50 1172 -37
rect 1228 37 1316 50
rect 1228 -37 1257 37
rect 1303 -37 1316 37
rect 1228 -50 1316 -37
<< pdiffc >>
rect -1303 -37 -1257 37
rect -1143 -37 -1097 37
rect -983 -37 -937 37
rect -823 -37 -777 37
rect -663 -37 -617 37
rect -503 -37 -457 37
rect -343 -37 -297 37
rect -183 -37 -137 37
rect -23 -37 23 37
rect 137 -37 183 37
rect 297 -37 343 37
rect 457 -37 503 37
rect 617 -37 663 37
rect 777 -37 823 37
rect 937 -37 983 37
rect 1097 -37 1143 37
rect 1257 -37 1303 37
<< polysilicon >>
rect -1228 50 -1172 94
rect -1068 50 -1012 94
rect -908 50 -852 94
rect -748 50 -692 94
rect -588 50 -532 94
rect -428 50 -372 94
rect -268 50 -212 94
rect -108 50 -52 94
rect 52 50 108 94
rect 212 50 268 94
rect 372 50 428 94
rect 532 50 588 94
rect 692 50 748 94
rect 852 50 908 94
rect 1012 50 1068 94
rect 1172 50 1228 94
rect -1228 -94 -1172 -50
rect -1068 -94 -1012 -50
rect -908 -94 -852 -50
rect -748 -94 -692 -50
rect -588 -94 -532 -50
rect -428 -94 -372 -50
rect -268 -94 -212 -50
rect -108 -94 -52 -50
rect 52 -94 108 -50
rect 212 -94 268 -50
rect 372 -94 428 -50
rect 532 -94 588 -50
rect 692 -94 748 -50
rect 852 -94 908 -50
rect 1012 -94 1068 -50
rect 1172 -94 1228 -50
<< metal1 >>
rect -1303 37 -1257 48
rect -1303 -48 -1257 -37
rect -1143 37 -1097 48
rect -1143 -48 -1097 -37
rect -983 37 -937 48
rect -983 -48 -937 -37
rect -823 37 -777 48
rect -823 -48 -777 -37
rect -663 37 -617 48
rect -663 -48 -617 -37
rect -503 37 -457 48
rect -503 -48 -457 -37
rect -343 37 -297 48
rect -343 -48 -297 -37
rect -183 37 -137 48
rect -183 -48 -137 -37
rect -23 37 23 48
rect -23 -48 23 -37
rect 137 37 183 48
rect 137 -48 183 -37
rect 297 37 343 48
rect 297 -48 343 -37
rect 457 37 503 48
rect 457 -48 503 -37
rect 617 37 663 48
rect 617 -48 663 -37
rect 777 37 823 48
rect 777 -48 823 -37
rect 937 37 983 48
rect 937 -48 983 -37
rect 1097 37 1143 48
rect 1097 -48 1143 -37
rect 1257 37 1303 48
rect 1257 -48 1303 -37
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 0.500 l 0.280 m 1 nf 16 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
