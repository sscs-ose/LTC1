magic
tech gf180mcuC
magscale 1 10
timestamp 1699351161
<< nwell >>
rect 34658 11207 34858 11407
rect 35028 11207 35228 11407
rect 35398 11207 35598 11407
rect 35768 11207 35968 11407
rect 36138 11207 36338 11407
rect 36508 11207 36708 11407
rect 36878 11207 37078 11407
rect 37248 11207 37448 11407
rect 37618 11207 37818 11407
rect 37988 11207 38188 11407
rect 38358 11207 38558 11407
rect 38728 11207 38928 11407
rect 39098 11207 39298 11407
rect 39468 11207 39668 11407
rect 39838 11207 40038 11407
rect 40208 11207 40408 11407
rect 40578 11207 40778 11407
rect 40948 11207 41148 11407
rect 41318 11207 41518 11407
rect 41688 11207 41888 11407
rect 42058 11207 42258 11407
rect 42428 11207 42628 11407
rect 42798 11207 42998 11407
rect 34658 10826 34858 11026
rect 35028 10826 35228 11026
rect 35398 10826 35598 11026
rect 35768 10826 35968 11026
rect 36138 10826 36338 11026
rect 36508 10826 36708 11026
rect 36878 10826 37078 11026
rect 37248 10826 37448 11026
rect 37618 10826 37818 11026
rect 37988 10826 38188 11026
rect 38358 10826 38558 11026
rect 38728 10826 38928 11026
rect 39098 10826 39298 11026
rect 39468 10826 39668 11026
rect 39838 10826 40038 11026
rect 40208 10826 40408 11026
rect 40578 10826 40778 11026
rect 40948 10826 41148 11026
rect 41318 10826 41518 11026
rect 41688 10826 41888 11026
rect 42058 10826 42258 11026
rect 42428 10826 42628 11026
rect 42798 10826 42998 11026
rect 34658 10445 34858 10645
rect 35028 10445 35228 10645
rect 35398 10445 35598 10645
rect 35768 10445 35968 10645
rect 36138 10445 36338 10645
rect 36508 10445 36708 10645
rect 36878 10445 37078 10645
rect 37248 10445 37448 10645
rect 37618 10445 37818 10645
rect 37988 10445 38188 10645
rect 38358 10445 38558 10645
rect 38728 10445 38928 10645
rect 39098 10445 39298 10645
rect 39468 10445 39668 10645
rect 39838 10445 40038 10645
rect 40208 10445 40408 10645
rect 40578 10445 40778 10645
rect 40948 10445 41148 10645
rect 41318 10445 41518 10645
rect 41688 10445 41888 10645
rect 42058 10445 42258 10645
rect 42428 10445 42628 10645
rect 42798 10445 42998 10645
rect 43378 2071 43473 2203
<< psubdiff >>
rect 21556 -22872 21756 -22844
rect 21556 -23024 21576 -22872
rect 21729 -23024 21756 -22872
rect 21556 -23044 21756 -23024
rect 21841 -22872 22041 -22844
rect 21841 -23024 21861 -22872
rect 22014 -23024 22041 -22872
rect 21841 -23044 22041 -23024
rect 22126 -22872 22326 -22844
rect 22126 -23024 22146 -22872
rect 22299 -23024 22326 -22872
rect 22126 -23044 22326 -23024
rect 22411 -22872 22611 -22844
rect 22411 -23024 22431 -22872
rect 22584 -23024 22611 -22872
rect 22411 -23044 22611 -23024
rect 22696 -22872 22896 -22844
rect 22696 -23024 22716 -22872
rect 22869 -23024 22896 -22872
rect 22696 -23044 22896 -23024
rect 22981 -22872 23181 -22844
rect 22981 -23024 23001 -22872
rect 23154 -23024 23181 -22872
rect 22981 -23044 23181 -23024
rect 23266 -22872 23466 -22844
rect 23266 -23024 23286 -22872
rect 23439 -23024 23466 -22872
rect 23266 -23044 23466 -23024
rect 23551 -22872 23751 -22844
rect 23551 -23024 23571 -22872
rect 23724 -23024 23751 -22872
rect 23551 -23044 23751 -23024
rect 23836 -22872 24036 -22844
rect 23836 -23024 23856 -22872
rect 24009 -23024 24036 -22872
rect 23836 -23044 24036 -23024
rect 24121 -22872 24321 -22844
rect 24121 -23024 24141 -22872
rect 24294 -23024 24321 -22872
rect 24121 -23044 24321 -23024
rect 24406 -22872 24606 -22844
rect 24406 -23024 24426 -22872
rect 24579 -23024 24606 -22872
rect 24406 -23044 24606 -23024
rect 24691 -22872 24891 -22844
rect 24691 -23024 24711 -22872
rect 24864 -23024 24891 -22872
rect 24691 -23044 24891 -23024
rect 24976 -22872 25176 -22844
rect 24976 -23024 24996 -22872
rect 25149 -23024 25176 -22872
rect 24976 -23044 25176 -23024
rect 25261 -22872 25461 -22844
rect 25261 -23024 25281 -22872
rect 25434 -23024 25461 -22872
rect 25261 -23044 25461 -23024
rect 25546 -22872 25746 -22844
rect 25546 -23024 25566 -22872
rect 25719 -23024 25746 -22872
rect 25546 -23044 25746 -23024
rect 25831 -22872 26031 -22844
rect 25831 -23024 25851 -22872
rect 26004 -23024 26031 -22872
rect 25831 -23044 26031 -23024
rect 26116 -22872 26316 -22844
rect 26116 -23024 26136 -22872
rect 26289 -23024 26316 -22872
rect 26116 -23044 26316 -23024
rect 26401 -22872 26601 -22844
rect 26401 -23024 26421 -22872
rect 26574 -23024 26601 -22872
rect 26401 -23044 26601 -23024
rect 26686 -22872 26886 -22844
rect 26686 -23024 26706 -22872
rect 26859 -23024 26886 -22872
rect 26686 -23044 26886 -23024
rect 26971 -22872 27171 -22844
rect 26971 -23024 26991 -22872
rect 27144 -23024 27171 -22872
rect 26971 -23044 27171 -23024
rect 27256 -22872 27456 -22844
rect 27256 -23024 27276 -22872
rect 27429 -23024 27456 -22872
rect 27256 -23044 27456 -23024
rect 27541 -22872 27741 -22844
rect 27541 -23024 27561 -22872
rect 27714 -23024 27741 -22872
rect 27541 -23044 27741 -23024
rect 27826 -22872 28026 -22844
rect 27826 -23024 27846 -22872
rect 27999 -23024 28026 -22872
rect 27826 -23044 28026 -23024
rect 28111 -22872 28311 -22844
rect 28111 -23024 28131 -22872
rect 28284 -23024 28311 -22872
rect 28111 -23044 28311 -23024
rect 28396 -22872 28596 -22844
rect 28396 -23024 28416 -22872
rect 28569 -23024 28596 -22872
rect 28396 -23044 28596 -23024
rect 28681 -22872 28881 -22844
rect 28681 -23024 28701 -22872
rect 28854 -23024 28881 -22872
rect 28681 -23044 28881 -23024
rect 28966 -22872 29166 -22844
rect 28966 -23024 28986 -22872
rect 29139 -23024 29166 -22872
rect 28966 -23044 29166 -23024
rect 29251 -22872 29451 -22844
rect 29251 -23024 29271 -22872
rect 29424 -23024 29451 -22872
rect 29251 -23044 29451 -23024
rect 29536 -22872 29736 -22844
rect 29536 -23024 29556 -22872
rect 29709 -23024 29736 -22872
rect 29536 -23044 29736 -23024
rect 29821 -22872 30021 -22844
rect 29821 -23024 29841 -22872
rect 29994 -23024 30021 -22872
rect 29821 -23044 30021 -23024
rect 30106 -22872 30306 -22844
rect 30106 -23024 30126 -22872
rect 30279 -23024 30306 -22872
rect 30106 -23044 30306 -23024
rect 30391 -22872 30591 -22844
rect 30391 -23024 30411 -22872
rect 30564 -23024 30591 -22872
rect 30391 -23044 30591 -23024
rect 30676 -22872 30876 -22844
rect 30676 -23024 30696 -22872
rect 30849 -23024 30876 -22872
rect 30676 -23044 30876 -23024
rect 30961 -22872 31161 -22844
rect 30961 -23024 30981 -22872
rect 31134 -23024 31161 -22872
rect 30961 -23044 31161 -23024
rect 31246 -22872 31446 -22844
rect 31246 -23024 31266 -22872
rect 31419 -23024 31446 -22872
rect 31246 -23044 31446 -23024
rect 31531 -22872 31731 -22844
rect 31531 -23024 31551 -22872
rect 31704 -23024 31731 -22872
rect 31531 -23044 31731 -23024
rect 31816 -22872 32016 -22844
rect 31816 -23024 31836 -22872
rect 31989 -23024 32016 -22872
rect 31816 -23044 32016 -23024
rect 32101 -22872 32301 -22844
rect 32101 -23024 32121 -22872
rect 32274 -23024 32301 -22872
rect 32101 -23044 32301 -23024
rect 32386 -22872 32586 -22844
rect 32386 -23024 32406 -22872
rect 32559 -23024 32586 -22872
rect 32386 -23044 32586 -23024
rect 32671 -22872 32871 -22844
rect 32671 -23024 32691 -22872
rect 32844 -23024 32871 -22872
rect 32671 -23044 32871 -23024
rect 32956 -22872 33156 -22844
rect 32956 -23024 32976 -22872
rect 33129 -23024 33156 -22872
rect 32956 -23044 33156 -23024
rect 33241 -22872 33441 -22844
rect 33241 -23024 33261 -22872
rect 33414 -23024 33441 -22872
rect 33241 -23044 33441 -23024
rect 33526 -22872 33726 -22844
rect 33526 -23024 33546 -22872
rect 33699 -23024 33726 -22872
rect 33526 -23044 33726 -23024
rect 33811 -22872 34011 -22844
rect 33811 -23024 33831 -22872
rect 33984 -23024 34011 -22872
rect 33811 -23044 34011 -23024
rect 34096 -22872 34296 -22844
rect 34096 -23024 34116 -22872
rect 34269 -23024 34296 -22872
rect 34096 -23044 34296 -23024
rect 34381 -22872 34581 -22844
rect 34381 -23024 34401 -22872
rect 34554 -23024 34581 -22872
rect 34381 -23044 34581 -23024
rect 34666 -22872 34866 -22844
rect 34666 -23024 34686 -22872
rect 34839 -23024 34866 -22872
rect 34666 -23044 34866 -23024
rect 34951 -22872 35151 -22844
rect 34951 -23024 34971 -22872
rect 35124 -23024 35151 -22872
rect 34951 -23044 35151 -23024
rect 35236 -22872 35436 -22844
rect 35236 -23024 35256 -22872
rect 35409 -23024 35436 -22872
rect 35236 -23044 35436 -23024
rect 35521 -22872 35721 -22844
rect 35521 -23024 35541 -22872
rect 35694 -23024 35721 -22872
rect 35521 -23044 35721 -23024
rect 35806 -22872 36006 -22844
rect 35806 -23024 35826 -22872
rect 35979 -23024 36006 -22872
rect 35806 -23044 36006 -23024
rect 36091 -22872 36291 -22844
rect 36091 -23024 36111 -22872
rect 36264 -23024 36291 -22872
rect 36091 -23044 36291 -23024
rect 36376 -22872 36576 -22844
rect 36376 -23024 36396 -22872
rect 36549 -23024 36576 -22872
rect 36376 -23044 36576 -23024
rect 36661 -22872 36861 -22844
rect 36661 -23024 36681 -22872
rect 36834 -23024 36861 -22872
rect 36661 -23044 36861 -23024
rect 36946 -22872 37146 -22844
rect 36946 -23024 36966 -22872
rect 37119 -23024 37146 -22872
rect 36946 -23044 37146 -23024
rect 37231 -22872 37431 -22844
rect 37231 -23024 37251 -22872
rect 37404 -23024 37431 -22872
rect 37231 -23044 37431 -23024
rect 37516 -22872 37716 -22844
rect 37516 -23024 37536 -22872
rect 37689 -23024 37716 -22872
rect 37516 -23044 37716 -23024
rect 37801 -22872 38001 -22844
rect 37801 -23024 37821 -22872
rect 37974 -23024 38001 -22872
rect 37801 -23044 38001 -23024
rect 38086 -22872 38286 -22844
rect 38086 -23024 38106 -22872
rect 38259 -23024 38286 -22872
rect 38086 -23044 38286 -23024
rect 38371 -22872 38571 -22844
rect 38371 -23024 38391 -22872
rect 38544 -23024 38571 -22872
rect 38371 -23044 38571 -23024
rect 38656 -22872 38856 -22844
rect 38656 -23024 38676 -22872
rect 38829 -23024 38856 -22872
rect 38656 -23044 38856 -23024
rect 38941 -22872 39141 -22844
rect 38941 -23024 38961 -22872
rect 39114 -23024 39141 -22872
rect 38941 -23044 39141 -23024
rect 39226 -22872 39426 -22844
rect 39226 -23024 39246 -22872
rect 39399 -23024 39426 -22872
rect 39226 -23044 39426 -23024
rect 39511 -22872 39711 -22844
rect 39511 -23024 39531 -22872
rect 39684 -23024 39711 -22872
rect 39511 -23044 39711 -23024
rect 39796 -22872 39996 -22844
rect 39796 -23024 39816 -22872
rect 39969 -23024 39996 -22872
rect 39796 -23044 39996 -23024
rect 40081 -22872 40281 -22844
rect 40081 -23024 40101 -22872
rect 40254 -23024 40281 -22872
rect 40081 -23044 40281 -23024
rect 40366 -22872 40566 -22844
rect 40366 -23024 40386 -22872
rect 40539 -23024 40566 -22872
rect 40366 -23044 40566 -23024
rect 40651 -22872 40851 -22844
rect 40651 -23024 40671 -22872
rect 40824 -23024 40851 -22872
rect 40651 -23044 40851 -23024
rect 40936 -22872 41136 -22844
rect 40936 -23024 40956 -22872
rect 41109 -23024 41136 -22872
rect 40936 -23044 41136 -23024
rect 41221 -22872 41421 -22844
rect 41221 -23024 41241 -22872
rect 41394 -23024 41421 -22872
rect 41221 -23044 41421 -23024
rect 41506 -22872 41706 -22844
rect 41506 -23024 41526 -22872
rect 41679 -23024 41706 -22872
rect 41506 -23044 41706 -23024
rect 41791 -22872 41991 -22844
rect 41791 -23024 41811 -22872
rect 41964 -23024 41991 -22872
rect 41791 -23044 41991 -23024
rect 42076 -22872 42276 -22844
rect 42076 -23024 42096 -22872
rect 42249 -23024 42276 -22872
rect 42076 -23044 42276 -23024
rect 42361 -22872 42561 -22844
rect 42361 -23024 42381 -22872
rect 42534 -23024 42561 -22872
rect 42361 -23044 42561 -23024
rect 42646 -22872 42846 -22844
rect 42646 -23024 42666 -22872
rect 42819 -23024 42846 -22872
rect 42646 -23044 42846 -23024
rect 42931 -22872 43131 -22844
rect 42931 -23024 42951 -22872
rect 43104 -23024 43131 -22872
rect 42931 -23044 43131 -23024
rect 43216 -22872 43416 -22844
rect 43216 -23024 43236 -22872
rect 43389 -23024 43416 -22872
rect 43216 -23044 43416 -23024
rect 43501 -22872 43701 -22844
rect 43501 -23024 43521 -22872
rect 43674 -23024 43701 -22872
rect 43501 -23044 43701 -23024
rect 43786 -22872 43986 -22844
rect 43786 -23024 43806 -22872
rect 43959 -23024 43986 -22872
rect 43786 -23044 43986 -23024
rect 44071 -22872 44271 -22844
rect 44071 -23024 44091 -22872
rect 44244 -23024 44271 -22872
rect 44071 -23044 44271 -23024
rect 44356 -22872 44556 -22844
rect 44356 -23024 44376 -22872
rect 44529 -23024 44556 -22872
rect 44356 -23044 44556 -23024
rect 44641 -22872 44841 -22844
rect 44641 -23024 44661 -22872
rect 44814 -23024 44841 -22872
rect 44641 -23044 44841 -23024
rect 44926 -22872 45126 -22844
rect 44926 -23024 44946 -22872
rect 45099 -23024 45126 -22872
rect 44926 -23044 45126 -23024
rect 45211 -22872 45411 -22844
rect 45211 -23024 45231 -22872
rect 45384 -23024 45411 -22872
rect 45211 -23044 45411 -23024
rect 45496 -22872 45696 -22844
rect 45496 -23024 45516 -22872
rect 45669 -23024 45696 -22872
rect 45496 -23044 45696 -23024
rect 45781 -22872 45981 -22844
rect 45781 -23024 45801 -22872
rect 45954 -23024 45981 -22872
rect 45781 -23044 45981 -23024
rect 46066 -22872 46266 -22844
rect 46066 -23024 46086 -22872
rect 46239 -23024 46266 -22872
rect 46066 -23044 46266 -23024
rect 46351 -22872 46551 -22844
rect 46351 -23024 46371 -22872
rect 46524 -23024 46551 -22872
rect 46351 -23044 46551 -23024
rect 46636 -22872 46836 -22844
rect 46636 -23024 46656 -22872
rect 46809 -23024 46836 -22872
rect 46636 -23044 46836 -23024
rect 46921 -22872 47121 -22844
rect 46921 -23024 46941 -22872
rect 47094 -23024 47121 -22872
rect 46921 -23044 47121 -23024
rect 47206 -22872 47406 -22844
rect 47206 -23024 47226 -22872
rect 47379 -23024 47406 -22872
rect 47206 -23044 47406 -23024
rect 47491 -22872 47691 -22844
rect 47491 -23024 47511 -22872
rect 47664 -23024 47691 -22872
rect 47491 -23044 47691 -23024
rect 47776 -22872 47976 -22844
rect 47776 -23024 47796 -22872
rect 47949 -23024 47976 -22872
rect 47776 -23044 47976 -23024
rect 48061 -22872 48261 -22844
rect 48061 -23024 48081 -22872
rect 48234 -23024 48261 -22872
rect 48061 -23044 48261 -23024
rect 48346 -22872 48546 -22844
rect 48346 -23024 48366 -22872
rect 48519 -23024 48546 -22872
rect 48346 -23044 48546 -23024
rect 48631 -22872 48831 -22844
rect 48631 -23024 48651 -22872
rect 48804 -23024 48831 -22872
rect 48631 -23044 48831 -23024
rect 48916 -22872 49116 -22844
rect 48916 -23024 48936 -22872
rect 49089 -23024 49116 -22872
rect 48916 -23044 49116 -23024
rect 49201 -22872 49401 -22844
rect 49201 -23024 49221 -22872
rect 49374 -23024 49401 -22872
rect 49201 -23044 49401 -23024
rect 49486 -22872 49686 -22844
rect 49486 -23024 49506 -22872
rect 49659 -23024 49686 -22872
rect 49486 -23044 49686 -23024
rect 49771 -22872 49971 -22844
rect 49771 -23024 49791 -22872
rect 49944 -23024 49971 -22872
rect 49771 -23044 49971 -23024
rect 50056 -22872 50256 -22844
rect 50056 -23024 50076 -22872
rect 50229 -23024 50256 -22872
rect 50056 -23044 50256 -23024
rect 50341 -22872 50541 -22844
rect 50341 -23024 50361 -22872
rect 50514 -23024 50541 -22872
rect 50341 -23044 50541 -23024
rect 50626 -22872 50826 -22844
rect 50626 -23024 50646 -22872
rect 50799 -23024 50826 -22872
rect 50626 -23044 50826 -23024
rect 50911 -22872 51111 -22844
rect 50911 -23024 50931 -22872
rect 51084 -23024 51111 -22872
rect 50911 -23044 51111 -23024
rect 51196 -22872 51396 -22844
rect 51196 -23024 51216 -22872
rect 51369 -23024 51396 -22872
rect 51196 -23044 51396 -23024
rect 51481 -22872 51681 -22844
rect 51481 -23024 51501 -22872
rect 51654 -23024 51681 -22872
rect 51481 -23044 51681 -23024
rect 51766 -22872 51966 -22844
rect 51766 -23024 51786 -22872
rect 51939 -23024 51966 -22872
rect 51766 -23044 51966 -23024
rect 52051 -22872 52251 -22844
rect 52051 -23024 52071 -22872
rect 52224 -23024 52251 -22872
rect 52051 -23044 52251 -23024
rect 52336 -22872 52536 -22844
rect 52336 -23024 52356 -22872
rect 52509 -23024 52536 -22872
rect 52336 -23044 52536 -23024
rect 52621 -22872 52821 -22844
rect 52621 -23024 52641 -22872
rect 52794 -23024 52821 -22872
rect 52621 -23044 52821 -23024
rect 52906 -22872 53106 -22844
rect 52906 -23024 52926 -22872
rect 53079 -23024 53106 -22872
rect 52906 -23044 53106 -23024
rect 53191 -22872 53391 -22844
rect 53191 -23024 53211 -22872
rect 53364 -23024 53391 -22872
rect 53191 -23044 53391 -23024
rect 53476 -22872 53676 -22844
rect 53476 -23024 53496 -22872
rect 53649 -23024 53676 -22872
rect 53476 -23044 53676 -23024
rect 53761 -22872 53961 -22844
rect 53761 -23024 53781 -22872
rect 53934 -23024 53961 -22872
rect 53761 -23044 53961 -23024
rect 54046 -22872 54246 -22844
rect 54046 -23024 54066 -22872
rect 54219 -23024 54246 -22872
rect 54046 -23044 54246 -23024
rect 54331 -22872 54531 -22844
rect 54331 -23024 54351 -22872
rect 54504 -23024 54531 -22872
rect 54331 -23044 54531 -23024
rect 54616 -22872 54816 -22844
rect 54616 -23024 54636 -22872
rect 54789 -23024 54816 -22872
rect 54616 -23044 54816 -23024
rect 54901 -22872 55101 -22844
rect 54901 -23024 54921 -22872
rect 55074 -23024 55101 -22872
rect 54901 -23044 55101 -23024
rect 55186 -22872 55386 -22844
rect 55186 -23024 55206 -22872
rect 55359 -23024 55386 -22872
rect 55186 -23044 55386 -23024
rect 55471 -22872 55671 -22844
rect 55471 -23024 55491 -22872
rect 55644 -23024 55671 -22872
rect 55471 -23044 55671 -23024
rect 55756 -22872 55956 -22844
rect 55756 -23024 55776 -22872
rect 55929 -23024 55956 -22872
rect 55756 -23044 55956 -23024
rect 21556 -23145 21756 -23117
rect 21556 -23297 21576 -23145
rect 21729 -23297 21756 -23145
rect 21556 -23317 21756 -23297
rect 21841 -23145 22041 -23117
rect 21841 -23297 21861 -23145
rect 22014 -23297 22041 -23145
rect 21841 -23317 22041 -23297
rect 22126 -23145 22326 -23117
rect 22126 -23297 22146 -23145
rect 22299 -23297 22326 -23145
rect 22126 -23317 22326 -23297
rect 22411 -23145 22611 -23117
rect 22411 -23297 22431 -23145
rect 22584 -23297 22611 -23145
rect 22411 -23317 22611 -23297
rect 22696 -23145 22896 -23117
rect 22696 -23297 22716 -23145
rect 22869 -23297 22896 -23145
rect 22696 -23317 22896 -23297
rect 22981 -23145 23181 -23117
rect 22981 -23297 23001 -23145
rect 23154 -23297 23181 -23145
rect 22981 -23317 23181 -23297
rect 23266 -23145 23466 -23117
rect 23266 -23297 23286 -23145
rect 23439 -23297 23466 -23145
rect 23266 -23317 23466 -23297
rect 23551 -23145 23751 -23117
rect 23551 -23297 23571 -23145
rect 23724 -23297 23751 -23145
rect 23551 -23317 23751 -23297
rect 23836 -23145 24036 -23117
rect 23836 -23297 23856 -23145
rect 24009 -23297 24036 -23145
rect 23836 -23317 24036 -23297
rect 24121 -23145 24321 -23117
rect 24121 -23297 24141 -23145
rect 24294 -23297 24321 -23145
rect 24121 -23317 24321 -23297
rect 24406 -23145 24606 -23117
rect 24406 -23297 24426 -23145
rect 24579 -23297 24606 -23145
rect 24406 -23317 24606 -23297
rect 24691 -23145 24891 -23117
rect 24691 -23297 24711 -23145
rect 24864 -23297 24891 -23145
rect 24691 -23317 24891 -23297
rect 24976 -23145 25176 -23117
rect 24976 -23297 24996 -23145
rect 25149 -23297 25176 -23145
rect 24976 -23317 25176 -23297
rect 25261 -23145 25461 -23117
rect 25261 -23297 25281 -23145
rect 25434 -23297 25461 -23145
rect 25261 -23317 25461 -23297
rect 25546 -23145 25746 -23117
rect 25546 -23297 25566 -23145
rect 25719 -23297 25746 -23145
rect 25546 -23317 25746 -23297
rect 25831 -23145 26031 -23117
rect 25831 -23297 25851 -23145
rect 26004 -23297 26031 -23145
rect 25831 -23317 26031 -23297
rect 26116 -23145 26316 -23117
rect 26116 -23297 26136 -23145
rect 26289 -23297 26316 -23145
rect 26116 -23317 26316 -23297
rect 26401 -23145 26601 -23117
rect 26401 -23297 26421 -23145
rect 26574 -23297 26601 -23145
rect 26401 -23317 26601 -23297
rect 26686 -23145 26886 -23117
rect 26686 -23297 26706 -23145
rect 26859 -23297 26886 -23145
rect 26686 -23317 26886 -23297
rect 26971 -23145 27171 -23117
rect 26971 -23297 26991 -23145
rect 27144 -23297 27171 -23145
rect 26971 -23317 27171 -23297
rect 27256 -23145 27456 -23117
rect 27256 -23297 27276 -23145
rect 27429 -23297 27456 -23145
rect 27256 -23317 27456 -23297
rect 27541 -23145 27741 -23117
rect 27541 -23297 27561 -23145
rect 27714 -23297 27741 -23145
rect 27541 -23317 27741 -23297
rect 27826 -23145 28026 -23117
rect 27826 -23297 27846 -23145
rect 27999 -23297 28026 -23145
rect 27826 -23317 28026 -23297
rect 28111 -23145 28311 -23117
rect 28111 -23297 28131 -23145
rect 28284 -23297 28311 -23145
rect 28111 -23317 28311 -23297
rect 28396 -23145 28596 -23117
rect 28396 -23297 28416 -23145
rect 28569 -23297 28596 -23145
rect 28396 -23317 28596 -23297
rect 28681 -23145 28881 -23117
rect 28681 -23297 28701 -23145
rect 28854 -23297 28881 -23145
rect 28681 -23317 28881 -23297
rect 28966 -23145 29166 -23117
rect 28966 -23297 28986 -23145
rect 29139 -23297 29166 -23145
rect 28966 -23317 29166 -23297
rect 29251 -23145 29451 -23117
rect 29251 -23297 29271 -23145
rect 29424 -23297 29451 -23145
rect 29251 -23317 29451 -23297
rect 29536 -23145 29736 -23117
rect 29536 -23297 29556 -23145
rect 29709 -23297 29736 -23145
rect 29536 -23317 29736 -23297
rect 29821 -23145 30021 -23117
rect 29821 -23297 29841 -23145
rect 29994 -23297 30021 -23145
rect 29821 -23317 30021 -23297
rect 30106 -23145 30306 -23117
rect 30106 -23297 30126 -23145
rect 30279 -23297 30306 -23145
rect 30106 -23317 30306 -23297
rect 30391 -23145 30591 -23117
rect 30391 -23297 30411 -23145
rect 30564 -23297 30591 -23145
rect 30391 -23317 30591 -23297
rect 30676 -23145 30876 -23117
rect 30676 -23297 30696 -23145
rect 30849 -23297 30876 -23145
rect 30676 -23317 30876 -23297
rect 30961 -23145 31161 -23117
rect 30961 -23297 30981 -23145
rect 31134 -23297 31161 -23145
rect 30961 -23317 31161 -23297
rect 31246 -23145 31446 -23117
rect 31246 -23297 31266 -23145
rect 31419 -23297 31446 -23145
rect 31246 -23317 31446 -23297
rect 31531 -23145 31731 -23117
rect 31531 -23297 31551 -23145
rect 31704 -23297 31731 -23145
rect 31531 -23317 31731 -23297
rect 31816 -23145 32016 -23117
rect 31816 -23297 31836 -23145
rect 31989 -23297 32016 -23145
rect 31816 -23317 32016 -23297
rect 32101 -23145 32301 -23117
rect 32101 -23297 32121 -23145
rect 32274 -23297 32301 -23145
rect 32101 -23317 32301 -23297
rect 32386 -23145 32586 -23117
rect 32386 -23297 32406 -23145
rect 32559 -23297 32586 -23145
rect 32386 -23317 32586 -23297
rect 32671 -23145 32871 -23117
rect 32671 -23297 32691 -23145
rect 32844 -23297 32871 -23145
rect 32671 -23317 32871 -23297
rect 32956 -23145 33156 -23117
rect 32956 -23297 32976 -23145
rect 33129 -23297 33156 -23145
rect 32956 -23317 33156 -23297
rect 33241 -23145 33441 -23117
rect 33241 -23297 33261 -23145
rect 33414 -23297 33441 -23145
rect 33241 -23317 33441 -23297
rect 33526 -23145 33726 -23117
rect 33526 -23297 33546 -23145
rect 33699 -23297 33726 -23145
rect 33526 -23317 33726 -23297
rect 33811 -23145 34011 -23117
rect 33811 -23297 33831 -23145
rect 33984 -23297 34011 -23145
rect 33811 -23317 34011 -23297
rect 34096 -23145 34296 -23117
rect 34096 -23297 34116 -23145
rect 34269 -23297 34296 -23145
rect 34096 -23317 34296 -23297
rect 34381 -23145 34581 -23117
rect 34381 -23297 34401 -23145
rect 34554 -23297 34581 -23145
rect 34381 -23317 34581 -23297
rect 34666 -23145 34866 -23117
rect 34666 -23297 34686 -23145
rect 34839 -23297 34866 -23145
rect 34666 -23317 34866 -23297
rect 34951 -23145 35151 -23117
rect 34951 -23297 34971 -23145
rect 35124 -23297 35151 -23145
rect 34951 -23317 35151 -23297
rect 35236 -23145 35436 -23117
rect 35236 -23297 35256 -23145
rect 35409 -23297 35436 -23145
rect 35236 -23317 35436 -23297
rect 35521 -23145 35721 -23117
rect 35521 -23297 35541 -23145
rect 35694 -23297 35721 -23145
rect 35521 -23317 35721 -23297
rect 35806 -23145 36006 -23117
rect 35806 -23297 35826 -23145
rect 35979 -23297 36006 -23145
rect 35806 -23317 36006 -23297
rect 36091 -23145 36291 -23117
rect 36091 -23297 36111 -23145
rect 36264 -23297 36291 -23145
rect 36091 -23317 36291 -23297
rect 36376 -23145 36576 -23117
rect 36376 -23297 36396 -23145
rect 36549 -23297 36576 -23145
rect 36376 -23317 36576 -23297
rect 36661 -23145 36861 -23117
rect 36661 -23297 36681 -23145
rect 36834 -23297 36861 -23145
rect 36661 -23317 36861 -23297
rect 36946 -23145 37146 -23117
rect 36946 -23297 36966 -23145
rect 37119 -23297 37146 -23145
rect 36946 -23317 37146 -23297
rect 37231 -23145 37431 -23117
rect 37231 -23297 37251 -23145
rect 37404 -23297 37431 -23145
rect 37231 -23317 37431 -23297
rect 37516 -23145 37716 -23117
rect 37516 -23297 37536 -23145
rect 37689 -23297 37716 -23145
rect 37516 -23317 37716 -23297
rect 37801 -23145 38001 -23117
rect 37801 -23297 37821 -23145
rect 37974 -23297 38001 -23145
rect 37801 -23317 38001 -23297
rect 38086 -23145 38286 -23117
rect 38086 -23297 38106 -23145
rect 38259 -23297 38286 -23145
rect 38086 -23317 38286 -23297
rect 38371 -23145 38571 -23117
rect 38371 -23297 38391 -23145
rect 38544 -23297 38571 -23145
rect 38371 -23317 38571 -23297
rect 38656 -23145 38856 -23117
rect 38656 -23297 38676 -23145
rect 38829 -23297 38856 -23145
rect 38656 -23317 38856 -23297
rect 38941 -23145 39141 -23117
rect 38941 -23297 38961 -23145
rect 39114 -23297 39141 -23145
rect 38941 -23317 39141 -23297
rect 39226 -23145 39426 -23117
rect 39226 -23297 39246 -23145
rect 39399 -23297 39426 -23145
rect 39226 -23317 39426 -23297
rect 39511 -23145 39711 -23117
rect 39511 -23297 39531 -23145
rect 39684 -23297 39711 -23145
rect 39511 -23317 39711 -23297
rect 39796 -23145 39996 -23117
rect 39796 -23297 39816 -23145
rect 39969 -23297 39996 -23145
rect 39796 -23317 39996 -23297
rect 40081 -23145 40281 -23117
rect 40081 -23297 40101 -23145
rect 40254 -23297 40281 -23145
rect 40081 -23317 40281 -23297
rect 40366 -23145 40566 -23117
rect 40366 -23297 40386 -23145
rect 40539 -23297 40566 -23145
rect 40366 -23317 40566 -23297
rect 40651 -23145 40851 -23117
rect 40651 -23297 40671 -23145
rect 40824 -23297 40851 -23145
rect 40651 -23317 40851 -23297
rect 40936 -23145 41136 -23117
rect 40936 -23297 40956 -23145
rect 41109 -23297 41136 -23145
rect 40936 -23317 41136 -23297
rect 41221 -23145 41421 -23117
rect 41221 -23297 41241 -23145
rect 41394 -23297 41421 -23145
rect 41221 -23317 41421 -23297
rect 41506 -23145 41706 -23117
rect 41506 -23297 41526 -23145
rect 41679 -23297 41706 -23145
rect 41506 -23317 41706 -23297
rect 41791 -23145 41991 -23117
rect 41791 -23297 41811 -23145
rect 41964 -23297 41991 -23145
rect 41791 -23317 41991 -23297
rect 42076 -23145 42276 -23117
rect 42076 -23297 42096 -23145
rect 42249 -23297 42276 -23145
rect 42076 -23317 42276 -23297
rect 42361 -23145 42561 -23117
rect 42361 -23297 42381 -23145
rect 42534 -23297 42561 -23145
rect 42361 -23317 42561 -23297
rect 42646 -23145 42846 -23117
rect 42646 -23297 42666 -23145
rect 42819 -23297 42846 -23145
rect 42646 -23317 42846 -23297
rect 42931 -23145 43131 -23117
rect 42931 -23297 42951 -23145
rect 43104 -23297 43131 -23145
rect 42931 -23317 43131 -23297
rect 43216 -23145 43416 -23117
rect 43216 -23297 43236 -23145
rect 43389 -23297 43416 -23145
rect 43216 -23317 43416 -23297
rect 43501 -23145 43701 -23117
rect 43501 -23297 43521 -23145
rect 43674 -23297 43701 -23145
rect 43501 -23317 43701 -23297
rect 43786 -23145 43986 -23117
rect 43786 -23297 43806 -23145
rect 43959 -23297 43986 -23145
rect 43786 -23317 43986 -23297
rect 44071 -23145 44271 -23117
rect 44071 -23297 44091 -23145
rect 44244 -23297 44271 -23145
rect 44071 -23317 44271 -23297
rect 44356 -23145 44556 -23117
rect 44356 -23297 44376 -23145
rect 44529 -23297 44556 -23145
rect 44356 -23317 44556 -23297
rect 44641 -23145 44841 -23117
rect 44641 -23297 44661 -23145
rect 44814 -23297 44841 -23145
rect 44641 -23317 44841 -23297
rect 44926 -23145 45126 -23117
rect 44926 -23297 44946 -23145
rect 45099 -23297 45126 -23145
rect 44926 -23317 45126 -23297
rect 45211 -23145 45411 -23117
rect 45211 -23297 45231 -23145
rect 45384 -23297 45411 -23145
rect 45211 -23317 45411 -23297
rect 45496 -23145 45696 -23117
rect 45496 -23297 45516 -23145
rect 45669 -23297 45696 -23145
rect 45496 -23317 45696 -23297
rect 45781 -23145 45981 -23117
rect 45781 -23297 45801 -23145
rect 45954 -23297 45981 -23145
rect 45781 -23317 45981 -23297
rect 46066 -23145 46266 -23117
rect 46066 -23297 46086 -23145
rect 46239 -23297 46266 -23145
rect 46066 -23317 46266 -23297
rect 46351 -23145 46551 -23117
rect 46351 -23297 46371 -23145
rect 46524 -23297 46551 -23145
rect 46351 -23317 46551 -23297
rect 46636 -23145 46836 -23117
rect 46636 -23297 46656 -23145
rect 46809 -23297 46836 -23145
rect 46636 -23317 46836 -23297
rect 46921 -23145 47121 -23117
rect 46921 -23297 46941 -23145
rect 47094 -23297 47121 -23145
rect 46921 -23317 47121 -23297
rect 47206 -23145 47406 -23117
rect 47206 -23297 47226 -23145
rect 47379 -23297 47406 -23145
rect 47206 -23317 47406 -23297
rect 47491 -23145 47691 -23117
rect 47491 -23297 47511 -23145
rect 47664 -23297 47691 -23145
rect 47491 -23317 47691 -23297
rect 47776 -23145 47976 -23117
rect 47776 -23297 47796 -23145
rect 47949 -23297 47976 -23145
rect 47776 -23317 47976 -23297
rect 48061 -23145 48261 -23117
rect 48061 -23297 48081 -23145
rect 48234 -23297 48261 -23145
rect 48061 -23317 48261 -23297
rect 48346 -23145 48546 -23117
rect 48346 -23297 48366 -23145
rect 48519 -23297 48546 -23145
rect 48346 -23317 48546 -23297
rect 48631 -23145 48831 -23117
rect 48631 -23297 48651 -23145
rect 48804 -23297 48831 -23145
rect 48631 -23317 48831 -23297
rect 48916 -23145 49116 -23117
rect 48916 -23297 48936 -23145
rect 49089 -23297 49116 -23145
rect 48916 -23317 49116 -23297
rect 49201 -23145 49401 -23117
rect 49201 -23297 49221 -23145
rect 49374 -23297 49401 -23145
rect 49201 -23317 49401 -23297
rect 49486 -23145 49686 -23117
rect 49486 -23297 49506 -23145
rect 49659 -23297 49686 -23145
rect 49486 -23317 49686 -23297
rect 49771 -23145 49971 -23117
rect 49771 -23297 49791 -23145
rect 49944 -23297 49971 -23145
rect 49771 -23317 49971 -23297
rect 50056 -23145 50256 -23117
rect 50056 -23297 50076 -23145
rect 50229 -23297 50256 -23145
rect 50056 -23317 50256 -23297
rect 50341 -23145 50541 -23117
rect 50341 -23297 50361 -23145
rect 50514 -23297 50541 -23145
rect 50341 -23317 50541 -23297
rect 50626 -23145 50826 -23117
rect 50626 -23297 50646 -23145
rect 50799 -23297 50826 -23145
rect 50626 -23317 50826 -23297
rect 50911 -23145 51111 -23117
rect 50911 -23297 50931 -23145
rect 51084 -23297 51111 -23145
rect 50911 -23317 51111 -23297
rect 51196 -23145 51396 -23117
rect 51196 -23297 51216 -23145
rect 51369 -23297 51396 -23145
rect 51196 -23317 51396 -23297
rect 51481 -23145 51681 -23117
rect 51481 -23297 51501 -23145
rect 51654 -23297 51681 -23145
rect 51481 -23317 51681 -23297
rect 51766 -23145 51966 -23117
rect 51766 -23297 51786 -23145
rect 51939 -23297 51966 -23145
rect 51766 -23317 51966 -23297
rect 52051 -23145 52251 -23117
rect 52051 -23297 52071 -23145
rect 52224 -23297 52251 -23145
rect 52051 -23317 52251 -23297
rect 52336 -23145 52536 -23117
rect 52336 -23297 52356 -23145
rect 52509 -23297 52536 -23145
rect 52336 -23317 52536 -23297
rect 52621 -23145 52821 -23117
rect 52621 -23297 52641 -23145
rect 52794 -23297 52821 -23145
rect 52621 -23317 52821 -23297
rect 52906 -23145 53106 -23117
rect 52906 -23297 52926 -23145
rect 53079 -23297 53106 -23145
rect 52906 -23317 53106 -23297
rect 53191 -23145 53391 -23117
rect 53191 -23297 53211 -23145
rect 53364 -23297 53391 -23145
rect 53191 -23317 53391 -23297
rect 53476 -23145 53676 -23117
rect 53476 -23297 53496 -23145
rect 53649 -23297 53676 -23145
rect 53476 -23317 53676 -23297
rect 53761 -23145 53961 -23117
rect 53761 -23297 53781 -23145
rect 53934 -23297 53961 -23145
rect 53761 -23317 53961 -23297
rect 54046 -23145 54246 -23117
rect 54046 -23297 54066 -23145
rect 54219 -23297 54246 -23145
rect 54046 -23317 54246 -23297
rect 54331 -23145 54531 -23117
rect 54331 -23297 54351 -23145
rect 54504 -23297 54531 -23145
rect 54331 -23317 54531 -23297
rect 54616 -23145 54816 -23117
rect 54616 -23297 54636 -23145
rect 54789 -23297 54816 -23145
rect 54616 -23317 54816 -23297
rect 54901 -23145 55101 -23117
rect 54901 -23297 54921 -23145
rect 55074 -23297 55101 -23145
rect 54901 -23317 55101 -23297
rect 55186 -23145 55386 -23117
rect 55186 -23297 55206 -23145
rect 55359 -23297 55386 -23145
rect 55186 -23317 55386 -23297
rect 55471 -23145 55671 -23117
rect 55471 -23297 55491 -23145
rect 55644 -23297 55671 -23145
rect 55471 -23317 55671 -23297
rect 55756 -23145 55956 -23117
rect 55756 -23297 55776 -23145
rect 55929 -23297 55956 -23145
rect 55756 -23317 55956 -23297
rect 21556 -23418 21756 -23390
rect 21556 -23570 21576 -23418
rect 21729 -23570 21756 -23418
rect 21556 -23590 21756 -23570
rect 21841 -23418 22041 -23390
rect 21841 -23570 21861 -23418
rect 22014 -23570 22041 -23418
rect 21841 -23590 22041 -23570
rect 22126 -23418 22326 -23390
rect 22126 -23570 22146 -23418
rect 22299 -23570 22326 -23418
rect 22126 -23590 22326 -23570
rect 22411 -23418 22611 -23390
rect 22411 -23570 22431 -23418
rect 22584 -23570 22611 -23418
rect 22411 -23590 22611 -23570
rect 22696 -23418 22896 -23390
rect 22696 -23570 22716 -23418
rect 22869 -23570 22896 -23418
rect 22696 -23590 22896 -23570
rect 22981 -23418 23181 -23390
rect 22981 -23570 23001 -23418
rect 23154 -23570 23181 -23418
rect 22981 -23590 23181 -23570
rect 23266 -23418 23466 -23390
rect 23266 -23570 23286 -23418
rect 23439 -23570 23466 -23418
rect 23266 -23590 23466 -23570
rect 23551 -23418 23751 -23390
rect 23551 -23570 23571 -23418
rect 23724 -23570 23751 -23418
rect 23551 -23590 23751 -23570
rect 23836 -23418 24036 -23390
rect 23836 -23570 23856 -23418
rect 24009 -23570 24036 -23418
rect 23836 -23590 24036 -23570
rect 24121 -23418 24321 -23390
rect 24121 -23570 24141 -23418
rect 24294 -23570 24321 -23418
rect 24121 -23590 24321 -23570
rect 24406 -23418 24606 -23390
rect 24406 -23570 24426 -23418
rect 24579 -23570 24606 -23418
rect 24406 -23590 24606 -23570
rect 24691 -23418 24891 -23390
rect 24691 -23570 24711 -23418
rect 24864 -23570 24891 -23418
rect 24691 -23590 24891 -23570
rect 24976 -23418 25176 -23390
rect 24976 -23570 24996 -23418
rect 25149 -23570 25176 -23418
rect 24976 -23590 25176 -23570
rect 25261 -23418 25461 -23390
rect 25261 -23570 25281 -23418
rect 25434 -23570 25461 -23418
rect 25261 -23590 25461 -23570
rect 25546 -23418 25746 -23390
rect 25546 -23570 25566 -23418
rect 25719 -23570 25746 -23418
rect 25546 -23590 25746 -23570
rect 25831 -23418 26031 -23390
rect 25831 -23570 25851 -23418
rect 26004 -23570 26031 -23418
rect 25831 -23590 26031 -23570
rect 26116 -23418 26316 -23390
rect 26116 -23570 26136 -23418
rect 26289 -23570 26316 -23418
rect 26116 -23590 26316 -23570
rect 26401 -23418 26601 -23390
rect 26401 -23570 26421 -23418
rect 26574 -23570 26601 -23418
rect 26401 -23590 26601 -23570
rect 26686 -23418 26886 -23390
rect 26686 -23570 26706 -23418
rect 26859 -23570 26886 -23418
rect 26686 -23590 26886 -23570
rect 26971 -23418 27171 -23390
rect 26971 -23570 26991 -23418
rect 27144 -23570 27171 -23418
rect 26971 -23590 27171 -23570
rect 27256 -23418 27456 -23390
rect 27256 -23570 27276 -23418
rect 27429 -23570 27456 -23418
rect 27256 -23590 27456 -23570
rect 27541 -23418 27741 -23390
rect 27541 -23570 27561 -23418
rect 27714 -23570 27741 -23418
rect 27541 -23590 27741 -23570
rect 27826 -23418 28026 -23390
rect 27826 -23570 27846 -23418
rect 27999 -23570 28026 -23418
rect 27826 -23590 28026 -23570
rect 28111 -23418 28311 -23390
rect 28111 -23570 28131 -23418
rect 28284 -23570 28311 -23418
rect 28111 -23590 28311 -23570
rect 28396 -23418 28596 -23390
rect 28396 -23570 28416 -23418
rect 28569 -23570 28596 -23418
rect 28396 -23590 28596 -23570
rect 28681 -23418 28881 -23390
rect 28681 -23570 28701 -23418
rect 28854 -23570 28881 -23418
rect 28681 -23590 28881 -23570
rect 28966 -23418 29166 -23390
rect 28966 -23570 28986 -23418
rect 29139 -23570 29166 -23418
rect 28966 -23590 29166 -23570
rect 29251 -23418 29451 -23390
rect 29251 -23570 29271 -23418
rect 29424 -23570 29451 -23418
rect 29251 -23590 29451 -23570
rect 29536 -23418 29736 -23390
rect 29536 -23570 29556 -23418
rect 29709 -23570 29736 -23418
rect 29536 -23590 29736 -23570
rect 29821 -23418 30021 -23390
rect 29821 -23570 29841 -23418
rect 29994 -23570 30021 -23418
rect 29821 -23590 30021 -23570
rect 30106 -23418 30306 -23390
rect 30106 -23570 30126 -23418
rect 30279 -23570 30306 -23418
rect 30106 -23590 30306 -23570
rect 30391 -23418 30591 -23390
rect 30391 -23570 30411 -23418
rect 30564 -23570 30591 -23418
rect 30391 -23590 30591 -23570
rect 30676 -23418 30876 -23390
rect 30676 -23570 30696 -23418
rect 30849 -23570 30876 -23418
rect 30676 -23590 30876 -23570
rect 30961 -23418 31161 -23390
rect 30961 -23570 30981 -23418
rect 31134 -23570 31161 -23418
rect 30961 -23590 31161 -23570
rect 31246 -23418 31446 -23390
rect 31246 -23570 31266 -23418
rect 31419 -23570 31446 -23418
rect 31246 -23590 31446 -23570
rect 31531 -23418 31731 -23390
rect 31531 -23570 31551 -23418
rect 31704 -23570 31731 -23418
rect 31531 -23590 31731 -23570
rect 31816 -23418 32016 -23390
rect 31816 -23570 31836 -23418
rect 31989 -23570 32016 -23418
rect 31816 -23590 32016 -23570
rect 32101 -23418 32301 -23390
rect 32101 -23570 32121 -23418
rect 32274 -23570 32301 -23418
rect 32101 -23590 32301 -23570
rect 32386 -23418 32586 -23390
rect 32386 -23570 32406 -23418
rect 32559 -23570 32586 -23418
rect 32386 -23590 32586 -23570
rect 32671 -23418 32871 -23390
rect 32671 -23570 32691 -23418
rect 32844 -23570 32871 -23418
rect 32671 -23590 32871 -23570
rect 32956 -23418 33156 -23390
rect 32956 -23570 32976 -23418
rect 33129 -23570 33156 -23418
rect 32956 -23590 33156 -23570
rect 33241 -23418 33441 -23390
rect 33241 -23570 33261 -23418
rect 33414 -23570 33441 -23418
rect 33241 -23590 33441 -23570
rect 33526 -23418 33726 -23390
rect 33526 -23570 33546 -23418
rect 33699 -23570 33726 -23418
rect 33526 -23590 33726 -23570
rect 33811 -23418 34011 -23390
rect 33811 -23570 33831 -23418
rect 33984 -23570 34011 -23418
rect 33811 -23590 34011 -23570
rect 34096 -23418 34296 -23390
rect 34096 -23570 34116 -23418
rect 34269 -23570 34296 -23418
rect 34096 -23590 34296 -23570
rect 34381 -23418 34581 -23390
rect 34381 -23570 34401 -23418
rect 34554 -23570 34581 -23418
rect 34381 -23590 34581 -23570
rect 34666 -23418 34866 -23390
rect 34666 -23570 34686 -23418
rect 34839 -23570 34866 -23418
rect 34666 -23590 34866 -23570
rect 34951 -23418 35151 -23390
rect 34951 -23570 34971 -23418
rect 35124 -23570 35151 -23418
rect 34951 -23590 35151 -23570
rect 35236 -23418 35436 -23390
rect 35236 -23570 35256 -23418
rect 35409 -23570 35436 -23418
rect 35236 -23590 35436 -23570
rect 35521 -23418 35721 -23390
rect 35521 -23570 35541 -23418
rect 35694 -23570 35721 -23418
rect 35521 -23590 35721 -23570
rect 35806 -23418 36006 -23390
rect 35806 -23570 35826 -23418
rect 35979 -23570 36006 -23418
rect 35806 -23590 36006 -23570
rect 36091 -23418 36291 -23390
rect 36091 -23570 36111 -23418
rect 36264 -23570 36291 -23418
rect 36091 -23590 36291 -23570
rect 36376 -23418 36576 -23390
rect 36376 -23570 36396 -23418
rect 36549 -23570 36576 -23418
rect 36376 -23590 36576 -23570
rect 36661 -23418 36861 -23390
rect 36661 -23570 36681 -23418
rect 36834 -23570 36861 -23418
rect 36661 -23590 36861 -23570
rect 36946 -23418 37146 -23390
rect 36946 -23570 36966 -23418
rect 37119 -23570 37146 -23418
rect 36946 -23590 37146 -23570
rect 37231 -23418 37431 -23390
rect 37231 -23570 37251 -23418
rect 37404 -23570 37431 -23418
rect 37231 -23590 37431 -23570
rect 37516 -23418 37716 -23390
rect 37516 -23570 37536 -23418
rect 37689 -23570 37716 -23418
rect 37516 -23590 37716 -23570
rect 37801 -23418 38001 -23390
rect 37801 -23570 37821 -23418
rect 37974 -23570 38001 -23418
rect 37801 -23590 38001 -23570
rect 38086 -23418 38286 -23390
rect 38086 -23570 38106 -23418
rect 38259 -23570 38286 -23418
rect 38086 -23590 38286 -23570
rect 38371 -23418 38571 -23390
rect 38371 -23570 38391 -23418
rect 38544 -23570 38571 -23418
rect 38371 -23590 38571 -23570
rect 38656 -23418 38856 -23390
rect 38656 -23570 38676 -23418
rect 38829 -23570 38856 -23418
rect 38656 -23590 38856 -23570
rect 38941 -23418 39141 -23390
rect 38941 -23570 38961 -23418
rect 39114 -23570 39141 -23418
rect 38941 -23590 39141 -23570
rect 39226 -23418 39426 -23390
rect 39226 -23570 39246 -23418
rect 39399 -23570 39426 -23418
rect 39226 -23590 39426 -23570
rect 39511 -23418 39711 -23390
rect 39511 -23570 39531 -23418
rect 39684 -23570 39711 -23418
rect 39511 -23590 39711 -23570
rect 39796 -23418 39996 -23390
rect 39796 -23570 39816 -23418
rect 39969 -23570 39996 -23418
rect 39796 -23590 39996 -23570
rect 40081 -23418 40281 -23390
rect 40081 -23570 40101 -23418
rect 40254 -23570 40281 -23418
rect 40081 -23590 40281 -23570
rect 40366 -23418 40566 -23390
rect 40366 -23570 40386 -23418
rect 40539 -23570 40566 -23418
rect 40366 -23590 40566 -23570
rect 40651 -23418 40851 -23390
rect 40651 -23570 40671 -23418
rect 40824 -23570 40851 -23418
rect 40651 -23590 40851 -23570
rect 40936 -23418 41136 -23390
rect 40936 -23570 40956 -23418
rect 41109 -23570 41136 -23418
rect 40936 -23590 41136 -23570
rect 41221 -23418 41421 -23390
rect 41221 -23570 41241 -23418
rect 41394 -23570 41421 -23418
rect 41221 -23590 41421 -23570
rect 41506 -23418 41706 -23390
rect 41506 -23570 41526 -23418
rect 41679 -23570 41706 -23418
rect 41506 -23590 41706 -23570
rect 41791 -23418 41991 -23390
rect 41791 -23570 41811 -23418
rect 41964 -23570 41991 -23418
rect 41791 -23590 41991 -23570
rect 42076 -23418 42276 -23390
rect 42076 -23570 42096 -23418
rect 42249 -23570 42276 -23418
rect 42076 -23590 42276 -23570
rect 42361 -23418 42561 -23390
rect 42361 -23570 42381 -23418
rect 42534 -23570 42561 -23418
rect 42361 -23590 42561 -23570
rect 42646 -23418 42846 -23390
rect 42646 -23570 42666 -23418
rect 42819 -23570 42846 -23418
rect 42646 -23590 42846 -23570
rect 42931 -23418 43131 -23390
rect 42931 -23570 42951 -23418
rect 43104 -23570 43131 -23418
rect 42931 -23590 43131 -23570
rect 43216 -23418 43416 -23390
rect 43216 -23570 43236 -23418
rect 43389 -23570 43416 -23418
rect 43216 -23590 43416 -23570
rect 43501 -23418 43701 -23390
rect 43501 -23570 43521 -23418
rect 43674 -23570 43701 -23418
rect 43501 -23590 43701 -23570
rect 43786 -23418 43986 -23390
rect 43786 -23570 43806 -23418
rect 43959 -23570 43986 -23418
rect 43786 -23590 43986 -23570
rect 44071 -23418 44271 -23390
rect 44071 -23570 44091 -23418
rect 44244 -23570 44271 -23418
rect 44071 -23590 44271 -23570
rect 44356 -23418 44556 -23390
rect 44356 -23570 44376 -23418
rect 44529 -23570 44556 -23418
rect 44356 -23590 44556 -23570
rect 44641 -23418 44841 -23390
rect 44641 -23570 44661 -23418
rect 44814 -23570 44841 -23418
rect 44641 -23590 44841 -23570
rect 44926 -23418 45126 -23390
rect 44926 -23570 44946 -23418
rect 45099 -23570 45126 -23418
rect 44926 -23590 45126 -23570
rect 45211 -23418 45411 -23390
rect 45211 -23570 45231 -23418
rect 45384 -23570 45411 -23418
rect 45211 -23590 45411 -23570
rect 45496 -23418 45696 -23390
rect 45496 -23570 45516 -23418
rect 45669 -23570 45696 -23418
rect 45496 -23590 45696 -23570
rect 45781 -23418 45981 -23390
rect 45781 -23570 45801 -23418
rect 45954 -23570 45981 -23418
rect 45781 -23590 45981 -23570
rect 46066 -23418 46266 -23390
rect 46066 -23570 46086 -23418
rect 46239 -23570 46266 -23418
rect 46066 -23590 46266 -23570
rect 46351 -23418 46551 -23390
rect 46351 -23570 46371 -23418
rect 46524 -23570 46551 -23418
rect 46351 -23590 46551 -23570
rect 46636 -23418 46836 -23390
rect 46636 -23570 46656 -23418
rect 46809 -23570 46836 -23418
rect 46636 -23590 46836 -23570
rect 46921 -23418 47121 -23390
rect 46921 -23570 46941 -23418
rect 47094 -23570 47121 -23418
rect 46921 -23590 47121 -23570
rect 47206 -23418 47406 -23390
rect 47206 -23570 47226 -23418
rect 47379 -23570 47406 -23418
rect 47206 -23590 47406 -23570
rect 47491 -23418 47691 -23390
rect 47491 -23570 47511 -23418
rect 47664 -23570 47691 -23418
rect 47491 -23590 47691 -23570
rect 47776 -23418 47976 -23390
rect 47776 -23570 47796 -23418
rect 47949 -23570 47976 -23418
rect 47776 -23590 47976 -23570
rect 48061 -23418 48261 -23390
rect 48061 -23570 48081 -23418
rect 48234 -23570 48261 -23418
rect 48061 -23590 48261 -23570
rect 48346 -23418 48546 -23390
rect 48346 -23570 48366 -23418
rect 48519 -23570 48546 -23418
rect 48346 -23590 48546 -23570
rect 48631 -23418 48831 -23390
rect 48631 -23570 48651 -23418
rect 48804 -23570 48831 -23418
rect 48631 -23590 48831 -23570
rect 48916 -23418 49116 -23390
rect 48916 -23570 48936 -23418
rect 49089 -23570 49116 -23418
rect 48916 -23590 49116 -23570
rect 49201 -23418 49401 -23390
rect 49201 -23570 49221 -23418
rect 49374 -23570 49401 -23418
rect 49201 -23590 49401 -23570
rect 49486 -23418 49686 -23390
rect 49486 -23570 49506 -23418
rect 49659 -23570 49686 -23418
rect 49486 -23590 49686 -23570
rect 49771 -23418 49971 -23390
rect 49771 -23570 49791 -23418
rect 49944 -23570 49971 -23418
rect 49771 -23590 49971 -23570
rect 50056 -23418 50256 -23390
rect 50056 -23570 50076 -23418
rect 50229 -23570 50256 -23418
rect 50056 -23590 50256 -23570
rect 50341 -23418 50541 -23390
rect 50341 -23570 50361 -23418
rect 50514 -23570 50541 -23418
rect 50341 -23590 50541 -23570
rect 50626 -23418 50826 -23390
rect 50626 -23570 50646 -23418
rect 50799 -23570 50826 -23418
rect 50626 -23590 50826 -23570
rect 50911 -23418 51111 -23390
rect 50911 -23570 50931 -23418
rect 51084 -23570 51111 -23418
rect 50911 -23590 51111 -23570
rect 51196 -23418 51396 -23390
rect 51196 -23570 51216 -23418
rect 51369 -23570 51396 -23418
rect 51196 -23590 51396 -23570
rect 51481 -23418 51681 -23390
rect 51481 -23570 51501 -23418
rect 51654 -23570 51681 -23418
rect 51481 -23590 51681 -23570
rect 51766 -23418 51966 -23390
rect 51766 -23570 51786 -23418
rect 51939 -23570 51966 -23418
rect 51766 -23590 51966 -23570
rect 52051 -23418 52251 -23390
rect 52051 -23570 52071 -23418
rect 52224 -23570 52251 -23418
rect 52051 -23590 52251 -23570
rect 52336 -23418 52536 -23390
rect 52336 -23570 52356 -23418
rect 52509 -23570 52536 -23418
rect 52336 -23590 52536 -23570
rect 52621 -23418 52821 -23390
rect 52621 -23570 52641 -23418
rect 52794 -23570 52821 -23418
rect 52621 -23590 52821 -23570
rect 52906 -23418 53106 -23390
rect 52906 -23570 52926 -23418
rect 53079 -23570 53106 -23418
rect 52906 -23590 53106 -23570
rect 53191 -23418 53391 -23390
rect 53191 -23570 53211 -23418
rect 53364 -23570 53391 -23418
rect 53191 -23590 53391 -23570
rect 53476 -23418 53676 -23390
rect 53476 -23570 53496 -23418
rect 53649 -23570 53676 -23418
rect 53476 -23590 53676 -23570
rect 53761 -23418 53961 -23390
rect 53761 -23570 53781 -23418
rect 53934 -23570 53961 -23418
rect 53761 -23590 53961 -23570
rect 54046 -23418 54246 -23390
rect 54046 -23570 54066 -23418
rect 54219 -23570 54246 -23418
rect 54046 -23590 54246 -23570
rect 54331 -23418 54531 -23390
rect 54331 -23570 54351 -23418
rect 54504 -23570 54531 -23418
rect 54331 -23590 54531 -23570
rect 54616 -23418 54816 -23390
rect 54616 -23570 54636 -23418
rect 54789 -23570 54816 -23418
rect 54616 -23590 54816 -23570
rect 54901 -23418 55101 -23390
rect 54901 -23570 54921 -23418
rect 55074 -23570 55101 -23418
rect 54901 -23590 55101 -23570
rect 55186 -23418 55386 -23390
rect 55186 -23570 55206 -23418
rect 55359 -23570 55386 -23418
rect 55186 -23590 55386 -23570
rect 55471 -23418 55671 -23390
rect 55471 -23570 55491 -23418
rect 55644 -23570 55671 -23418
rect 55471 -23590 55671 -23570
rect 55756 -23418 55956 -23390
rect 55756 -23570 55776 -23418
rect 55929 -23570 55956 -23418
rect 55756 -23590 55956 -23570
rect 21556 -23691 21756 -23663
rect 21556 -23843 21576 -23691
rect 21729 -23843 21756 -23691
rect 21556 -23863 21756 -23843
rect 21841 -23691 22041 -23663
rect 21841 -23843 21861 -23691
rect 22014 -23843 22041 -23691
rect 21841 -23863 22041 -23843
rect 22126 -23691 22326 -23663
rect 22126 -23843 22146 -23691
rect 22299 -23843 22326 -23691
rect 22126 -23863 22326 -23843
rect 22411 -23691 22611 -23663
rect 22411 -23843 22431 -23691
rect 22584 -23843 22611 -23691
rect 22411 -23863 22611 -23843
rect 22696 -23691 22896 -23663
rect 22696 -23843 22716 -23691
rect 22869 -23843 22896 -23691
rect 22696 -23863 22896 -23843
rect 22981 -23691 23181 -23663
rect 22981 -23843 23001 -23691
rect 23154 -23843 23181 -23691
rect 22981 -23863 23181 -23843
rect 23266 -23691 23466 -23663
rect 23266 -23843 23286 -23691
rect 23439 -23843 23466 -23691
rect 23266 -23863 23466 -23843
rect 23551 -23691 23751 -23663
rect 23551 -23843 23571 -23691
rect 23724 -23843 23751 -23691
rect 23551 -23863 23751 -23843
rect 23836 -23691 24036 -23663
rect 23836 -23843 23856 -23691
rect 24009 -23843 24036 -23691
rect 23836 -23863 24036 -23843
rect 24121 -23691 24321 -23663
rect 24121 -23843 24141 -23691
rect 24294 -23843 24321 -23691
rect 24121 -23863 24321 -23843
rect 24406 -23691 24606 -23663
rect 24406 -23843 24426 -23691
rect 24579 -23843 24606 -23691
rect 24406 -23863 24606 -23843
rect 24691 -23691 24891 -23663
rect 24691 -23843 24711 -23691
rect 24864 -23843 24891 -23691
rect 24691 -23863 24891 -23843
rect 24976 -23691 25176 -23663
rect 24976 -23843 24996 -23691
rect 25149 -23843 25176 -23691
rect 24976 -23863 25176 -23843
rect 25261 -23691 25461 -23663
rect 25261 -23843 25281 -23691
rect 25434 -23843 25461 -23691
rect 25261 -23863 25461 -23843
rect 25546 -23691 25746 -23663
rect 25546 -23843 25566 -23691
rect 25719 -23843 25746 -23691
rect 25546 -23863 25746 -23843
rect 25831 -23691 26031 -23663
rect 25831 -23843 25851 -23691
rect 26004 -23843 26031 -23691
rect 25831 -23863 26031 -23843
rect 26116 -23691 26316 -23663
rect 26116 -23843 26136 -23691
rect 26289 -23843 26316 -23691
rect 26116 -23863 26316 -23843
rect 26401 -23691 26601 -23663
rect 26401 -23843 26421 -23691
rect 26574 -23843 26601 -23691
rect 26401 -23863 26601 -23843
rect 26686 -23691 26886 -23663
rect 26686 -23843 26706 -23691
rect 26859 -23843 26886 -23691
rect 26686 -23863 26886 -23843
rect 26971 -23691 27171 -23663
rect 26971 -23843 26991 -23691
rect 27144 -23843 27171 -23691
rect 26971 -23863 27171 -23843
rect 27256 -23691 27456 -23663
rect 27256 -23843 27276 -23691
rect 27429 -23843 27456 -23691
rect 27256 -23863 27456 -23843
rect 27541 -23691 27741 -23663
rect 27541 -23843 27561 -23691
rect 27714 -23843 27741 -23691
rect 27541 -23863 27741 -23843
rect 27826 -23691 28026 -23663
rect 27826 -23843 27846 -23691
rect 27999 -23843 28026 -23691
rect 27826 -23863 28026 -23843
rect 28111 -23691 28311 -23663
rect 28111 -23843 28131 -23691
rect 28284 -23843 28311 -23691
rect 28111 -23863 28311 -23843
rect 28396 -23691 28596 -23663
rect 28396 -23843 28416 -23691
rect 28569 -23843 28596 -23691
rect 28396 -23863 28596 -23843
rect 28681 -23691 28881 -23663
rect 28681 -23843 28701 -23691
rect 28854 -23843 28881 -23691
rect 28681 -23863 28881 -23843
rect 28966 -23691 29166 -23663
rect 28966 -23843 28986 -23691
rect 29139 -23843 29166 -23691
rect 28966 -23863 29166 -23843
rect 29251 -23691 29451 -23663
rect 29251 -23843 29271 -23691
rect 29424 -23843 29451 -23691
rect 29251 -23863 29451 -23843
rect 29536 -23691 29736 -23663
rect 29536 -23843 29556 -23691
rect 29709 -23843 29736 -23691
rect 29536 -23863 29736 -23843
rect 29821 -23691 30021 -23663
rect 29821 -23843 29841 -23691
rect 29994 -23843 30021 -23691
rect 29821 -23863 30021 -23843
rect 30106 -23691 30306 -23663
rect 30106 -23843 30126 -23691
rect 30279 -23843 30306 -23691
rect 30106 -23863 30306 -23843
rect 30391 -23691 30591 -23663
rect 30391 -23843 30411 -23691
rect 30564 -23843 30591 -23691
rect 30391 -23863 30591 -23843
rect 30676 -23691 30876 -23663
rect 30676 -23843 30696 -23691
rect 30849 -23843 30876 -23691
rect 30676 -23863 30876 -23843
rect 30961 -23691 31161 -23663
rect 30961 -23843 30981 -23691
rect 31134 -23843 31161 -23691
rect 30961 -23863 31161 -23843
rect 31246 -23691 31446 -23663
rect 31246 -23843 31266 -23691
rect 31419 -23843 31446 -23691
rect 31246 -23863 31446 -23843
rect 31531 -23691 31731 -23663
rect 31531 -23843 31551 -23691
rect 31704 -23843 31731 -23691
rect 31531 -23863 31731 -23843
rect 31816 -23691 32016 -23663
rect 31816 -23843 31836 -23691
rect 31989 -23843 32016 -23691
rect 31816 -23863 32016 -23843
rect 32101 -23691 32301 -23663
rect 32101 -23843 32121 -23691
rect 32274 -23843 32301 -23691
rect 32101 -23863 32301 -23843
rect 32386 -23691 32586 -23663
rect 32386 -23843 32406 -23691
rect 32559 -23843 32586 -23691
rect 32386 -23863 32586 -23843
rect 32671 -23691 32871 -23663
rect 32671 -23843 32691 -23691
rect 32844 -23843 32871 -23691
rect 32671 -23863 32871 -23843
rect 32956 -23691 33156 -23663
rect 32956 -23843 32976 -23691
rect 33129 -23843 33156 -23691
rect 32956 -23863 33156 -23843
rect 33241 -23691 33441 -23663
rect 33241 -23843 33261 -23691
rect 33414 -23843 33441 -23691
rect 33241 -23863 33441 -23843
rect 33526 -23691 33726 -23663
rect 33526 -23843 33546 -23691
rect 33699 -23843 33726 -23691
rect 33526 -23863 33726 -23843
rect 33811 -23691 34011 -23663
rect 33811 -23843 33831 -23691
rect 33984 -23843 34011 -23691
rect 33811 -23863 34011 -23843
rect 34096 -23691 34296 -23663
rect 34096 -23843 34116 -23691
rect 34269 -23843 34296 -23691
rect 34096 -23863 34296 -23843
rect 34381 -23691 34581 -23663
rect 34381 -23843 34401 -23691
rect 34554 -23843 34581 -23691
rect 34381 -23863 34581 -23843
rect 34666 -23691 34866 -23663
rect 34666 -23843 34686 -23691
rect 34839 -23843 34866 -23691
rect 34666 -23863 34866 -23843
rect 34951 -23691 35151 -23663
rect 34951 -23843 34971 -23691
rect 35124 -23843 35151 -23691
rect 34951 -23863 35151 -23843
rect 35236 -23691 35436 -23663
rect 35236 -23843 35256 -23691
rect 35409 -23843 35436 -23691
rect 35236 -23863 35436 -23843
rect 35521 -23691 35721 -23663
rect 35521 -23843 35541 -23691
rect 35694 -23843 35721 -23691
rect 35521 -23863 35721 -23843
rect 35806 -23691 36006 -23663
rect 35806 -23843 35826 -23691
rect 35979 -23843 36006 -23691
rect 35806 -23863 36006 -23843
rect 36091 -23691 36291 -23663
rect 36091 -23843 36111 -23691
rect 36264 -23843 36291 -23691
rect 36091 -23863 36291 -23843
rect 36376 -23691 36576 -23663
rect 36376 -23843 36396 -23691
rect 36549 -23843 36576 -23691
rect 36376 -23863 36576 -23843
rect 36661 -23691 36861 -23663
rect 36661 -23843 36681 -23691
rect 36834 -23843 36861 -23691
rect 36661 -23863 36861 -23843
rect 36946 -23691 37146 -23663
rect 36946 -23843 36966 -23691
rect 37119 -23843 37146 -23691
rect 36946 -23863 37146 -23843
rect 37231 -23691 37431 -23663
rect 37231 -23843 37251 -23691
rect 37404 -23843 37431 -23691
rect 37231 -23863 37431 -23843
rect 37516 -23691 37716 -23663
rect 37516 -23843 37536 -23691
rect 37689 -23843 37716 -23691
rect 37516 -23863 37716 -23843
rect 37801 -23691 38001 -23663
rect 37801 -23843 37821 -23691
rect 37974 -23843 38001 -23691
rect 37801 -23863 38001 -23843
rect 38086 -23691 38286 -23663
rect 38086 -23843 38106 -23691
rect 38259 -23843 38286 -23691
rect 38086 -23863 38286 -23843
rect 38371 -23691 38571 -23663
rect 38371 -23843 38391 -23691
rect 38544 -23843 38571 -23691
rect 38371 -23863 38571 -23843
rect 38656 -23691 38856 -23663
rect 38656 -23843 38676 -23691
rect 38829 -23843 38856 -23691
rect 38656 -23863 38856 -23843
rect 38941 -23691 39141 -23663
rect 38941 -23843 38961 -23691
rect 39114 -23843 39141 -23691
rect 38941 -23863 39141 -23843
rect 39226 -23691 39426 -23663
rect 39226 -23843 39246 -23691
rect 39399 -23843 39426 -23691
rect 39226 -23863 39426 -23843
rect 39511 -23691 39711 -23663
rect 39511 -23843 39531 -23691
rect 39684 -23843 39711 -23691
rect 39511 -23863 39711 -23843
rect 39796 -23691 39996 -23663
rect 39796 -23843 39816 -23691
rect 39969 -23843 39996 -23691
rect 39796 -23863 39996 -23843
rect 40081 -23691 40281 -23663
rect 40081 -23843 40101 -23691
rect 40254 -23843 40281 -23691
rect 40081 -23863 40281 -23843
rect 40366 -23691 40566 -23663
rect 40366 -23843 40386 -23691
rect 40539 -23843 40566 -23691
rect 40366 -23863 40566 -23843
rect 40651 -23691 40851 -23663
rect 40651 -23843 40671 -23691
rect 40824 -23843 40851 -23691
rect 40651 -23863 40851 -23843
rect 40936 -23691 41136 -23663
rect 40936 -23843 40956 -23691
rect 41109 -23843 41136 -23691
rect 40936 -23863 41136 -23843
rect 41221 -23691 41421 -23663
rect 41221 -23843 41241 -23691
rect 41394 -23843 41421 -23691
rect 41221 -23863 41421 -23843
rect 41506 -23691 41706 -23663
rect 41506 -23843 41526 -23691
rect 41679 -23843 41706 -23691
rect 41506 -23863 41706 -23843
rect 41791 -23691 41991 -23663
rect 41791 -23843 41811 -23691
rect 41964 -23843 41991 -23691
rect 41791 -23863 41991 -23843
rect 42076 -23691 42276 -23663
rect 42076 -23843 42096 -23691
rect 42249 -23843 42276 -23691
rect 42076 -23863 42276 -23843
rect 42361 -23691 42561 -23663
rect 42361 -23843 42381 -23691
rect 42534 -23843 42561 -23691
rect 42361 -23863 42561 -23843
rect 42646 -23691 42846 -23663
rect 42646 -23843 42666 -23691
rect 42819 -23843 42846 -23691
rect 42646 -23863 42846 -23843
rect 42931 -23691 43131 -23663
rect 42931 -23843 42951 -23691
rect 43104 -23843 43131 -23691
rect 42931 -23863 43131 -23843
rect 43216 -23691 43416 -23663
rect 43216 -23843 43236 -23691
rect 43389 -23843 43416 -23691
rect 43216 -23863 43416 -23843
rect 43501 -23691 43701 -23663
rect 43501 -23843 43521 -23691
rect 43674 -23843 43701 -23691
rect 43501 -23863 43701 -23843
rect 43786 -23691 43986 -23663
rect 43786 -23843 43806 -23691
rect 43959 -23843 43986 -23691
rect 43786 -23863 43986 -23843
rect 44071 -23691 44271 -23663
rect 44071 -23843 44091 -23691
rect 44244 -23843 44271 -23691
rect 44071 -23863 44271 -23843
rect 44356 -23691 44556 -23663
rect 44356 -23843 44376 -23691
rect 44529 -23843 44556 -23691
rect 44356 -23863 44556 -23843
rect 44641 -23691 44841 -23663
rect 44641 -23843 44661 -23691
rect 44814 -23843 44841 -23691
rect 44641 -23863 44841 -23843
rect 44926 -23691 45126 -23663
rect 44926 -23843 44946 -23691
rect 45099 -23843 45126 -23691
rect 44926 -23863 45126 -23843
rect 45211 -23691 45411 -23663
rect 45211 -23843 45231 -23691
rect 45384 -23843 45411 -23691
rect 45211 -23863 45411 -23843
rect 45496 -23691 45696 -23663
rect 45496 -23843 45516 -23691
rect 45669 -23843 45696 -23691
rect 45496 -23863 45696 -23843
rect 45781 -23691 45981 -23663
rect 45781 -23843 45801 -23691
rect 45954 -23843 45981 -23691
rect 45781 -23863 45981 -23843
rect 46066 -23691 46266 -23663
rect 46066 -23843 46086 -23691
rect 46239 -23843 46266 -23691
rect 46066 -23863 46266 -23843
rect 46351 -23691 46551 -23663
rect 46351 -23843 46371 -23691
rect 46524 -23843 46551 -23691
rect 46351 -23863 46551 -23843
rect 46636 -23691 46836 -23663
rect 46636 -23843 46656 -23691
rect 46809 -23843 46836 -23691
rect 46636 -23863 46836 -23843
rect 46921 -23691 47121 -23663
rect 46921 -23843 46941 -23691
rect 47094 -23843 47121 -23691
rect 46921 -23863 47121 -23843
rect 47206 -23691 47406 -23663
rect 47206 -23843 47226 -23691
rect 47379 -23843 47406 -23691
rect 47206 -23863 47406 -23843
rect 47491 -23691 47691 -23663
rect 47491 -23843 47511 -23691
rect 47664 -23843 47691 -23691
rect 47491 -23863 47691 -23843
rect 47776 -23691 47976 -23663
rect 47776 -23843 47796 -23691
rect 47949 -23843 47976 -23691
rect 47776 -23863 47976 -23843
rect 48061 -23691 48261 -23663
rect 48061 -23843 48081 -23691
rect 48234 -23843 48261 -23691
rect 48061 -23863 48261 -23843
rect 48346 -23691 48546 -23663
rect 48346 -23843 48366 -23691
rect 48519 -23843 48546 -23691
rect 48346 -23863 48546 -23843
rect 48631 -23691 48831 -23663
rect 48631 -23843 48651 -23691
rect 48804 -23843 48831 -23691
rect 48631 -23863 48831 -23843
rect 48916 -23691 49116 -23663
rect 48916 -23843 48936 -23691
rect 49089 -23843 49116 -23691
rect 48916 -23863 49116 -23843
rect 49201 -23691 49401 -23663
rect 49201 -23843 49221 -23691
rect 49374 -23843 49401 -23691
rect 49201 -23863 49401 -23843
rect 49486 -23691 49686 -23663
rect 49486 -23843 49506 -23691
rect 49659 -23843 49686 -23691
rect 49486 -23863 49686 -23843
rect 49771 -23691 49971 -23663
rect 49771 -23843 49791 -23691
rect 49944 -23843 49971 -23691
rect 49771 -23863 49971 -23843
rect 50056 -23691 50256 -23663
rect 50056 -23843 50076 -23691
rect 50229 -23843 50256 -23691
rect 50056 -23863 50256 -23843
rect 50341 -23691 50541 -23663
rect 50341 -23843 50361 -23691
rect 50514 -23843 50541 -23691
rect 50341 -23863 50541 -23843
rect 50626 -23691 50826 -23663
rect 50626 -23843 50646 -23691
rect 50799 -23843 50826 -23691
rect 50626 -23863 50826 -23843
rect 50911 -23691 51111 -23663
rect 50911 -23843 50931 -23691
rect 51084 -23843 51111 -23691
rect 50911 -23863 51111 -23843
rect 51196 -23691 51396 -23663
rect 51196 -23843 51216 -23691
rect 51369 -23843 51396 -23691
rect 51196 -23863 51396 -23843
rect 51481 -23691 51681 -23663
rect 51481 -23843 51501 -23691
rect 51654 -23843 51681 -23691
rect 51481 -23863 51681 -23843
rect 51766 -23691 51966 -23663
rect 51766 -23843 51786 -23691
rect 51939 -23843 51966 -23691
rect 51766 -23863 51966 -23843
rect 52051 -23691 52251 -23663
rect 52051 -23843 52071 -23691
rect 52224 -23843 52251 -23691
rect 52051 -23863 52251 -23843
rect 52336 -23691 52536 -23663
rect 52336 -23843 52356 -23691
rect 52509 -23843 52536 -23691
rect 52336 -23863 52536 -23843
rect 52621 -23691 52821 -23663
rect 52621 -23843 52641 -23691
rect 52794 -23843 52821 -23691
rect 52621 -23863 52821 -23843
rect 52906 -23691 53106 -23663
rect 52906 -23843 52926 -23691
rect 53079 -23843 53106 -23691
rect 52906 -23863 53106 -23843
rect 53191 -23691 53391 -23663
rect 53191 -23843 53211 -23691
rect 53364 -23843 53391 -23691
rect 53191 -23863 53391 -23843
rect 53476 -23691 53676 -23663
rect 53476 -23843 53496 -23691
rect 53649 -23843 53676 -23691
rect 53476 -23863 53676 -23843
rect 53761 -23691 53961 -23663
rect 53761 -23843 53781 -23691
rect 53934 -23843 53961 -23691
rect 53761 -23863 53961 -23843
rect 54046 -23691 54246 -23663
rect 54046 -23843 54066 -23691
rect 54219 -23843 54246 -23691
rect 54046 -23863 54246 -23843
rect 54331 -23691 54531 -23663
rect 54331 -23843 54351 -23691
rect 54504 -23843 54531 -23691
rect 54331 -23863 54531 -23843
rect 54616 -23691 54816 -23663
rect 54616 -23843 54636 -23691
rect 54789 -23843 54816 -23691
rect 54616 -23863 54816 -23843
rect 54901 -23691 55101 -23663
rect 54901 -23843 54921 -23691
rect 55074 -23843 55101 -23691
rect 54901 -23863 55101 -23843
rect 55186 -23691 55386 -23663
rect 55186 -23843 55206 -23691
rect 55359 -23843 55386 -23691
rect 55186 -23863 55386 -23843
rect 55471 -23691 55671 -23663
rect 55471 -23843 55491 -23691
rect 55644 -23843 55671 -23691
rect 55471 -23863 55671 -23843
rect 55756 -23691 55956 -23663
rect 55756 -23843 55776 -23691
rect 55929 -23843 55956 -23691
rect 55756 -23863 55956 -23843
<< nsubdiff >>
rect 34683 11358 34828 11380
rect 34683 11261 34707 11358
rect 34805 11261 34828 11358
rect 34683 11236 34828 11261
rect 35053 11358 35198 11380
rect 35053 11261 35077 11358
rect 35175 11261 35198 11358
rect 35053 11236 35198 11261
rect 35423 11358 35568 11380
rect 35423 11261 35447 11358
rect 35545 11261 35568 11358
rect 35423 11236 35568 11261
rect 35793 11358 35938 11380
rect 35793 11261 35817 11358
rect 35915 11261 35938 11358
rect 35793 11236 35938 11261
rect 36163 11358 36308 11380
rect 36163 11261 36187 11358
rect 36285 11261 36308 11358
rect 36163 11236 36308 11261
rect 36533 11358 36678 11380
rect 36533 11261 36557 11358
rect 36655 11261 36678 11358
rect 36533 11236 36678 11261
rect 36903 11358 37048 11380
rect 36903 11261 36927 11358
rect 37025 11261 37048 11358
rect 36903 11236 37048 11261
rect 37273 11358 37418 11380
rect 37273 11261 37297 11358
rect 37395 11261 37418 11358
rect 37273 11236 37418 11261
rect 37643 11358 37788 11380
rect 37643 11261 37667 11358
rect 37765 11261 37788 11358
rect 37643 11236 37788 11261
rect 38013 11358 38158 11380
rect 38013 11261 38037 11358
rect 38135 11261 38158 11358
rect 38013 11236 38158 11261
rect 38383 11358 38528 11380
rect 38383 11261 38407 11358
rect 38505 11261 38528 11358
rect 38383 11236 38528 11261
rect 38753 11358 38898 11380
rect 38753 11261 38777 11358
rect 38875 11261 38898 11358
rect 38753 11236 38898 11261
rect 39123 11358 39268 11380
rect 39123 11261 39147 11358
rect 39245 11261 39268 11358
rect 39123 11236 39268 11261
rect 39493 11358 39638 11380
rect 39493 11261 39517 11358
rect 39615 11261 39638 11358
rect 39493 11236 39638 11261
rect 39863 11358 40008 11380
rect 39863 11261 39887 11358
rect 39985 11261 40008 11358
rect 39863 11236 40008 11261
rect 40233 11358 40378 11380
rect 40233 11261 40257 11358
rect 40355 11261 40378 11358
rect 40233 11236 40378 11261
rect 40603 11358 40748 11380
rect 40603 11261 40627 11358
rect 40725 11261 40748 11358
rect 40603 11236 40748 11261
rect 40973 11358 41118 11380
rect 40973 11261 40997 11358
rect 41095 11261 41118 11358
rect 40973 11236 41118 11261
rect 41343 11358 41488 11380
rect 41343 11261 41367 11358
rect 41465 11261 41488 11358
rect 41343 11236 41488 11261
rect 41713 11358 41858 11380
rect 41713 11261 41737 11358
rect 41835 11261 41858 11358
rect 41713 11236 41858 11261
rect 42083 11358 42228 11380
rect 42083 11261 42107 11358
rect 42205 11261 42228 11358
rect 42083 11236 42228 11261
rect 42453 11358 42598 11380
rect 42453 11261 42477 11358
rect 42575 11261 42598 11358
rect 42453 11236 42598 11261
rect 42823 11358 42968 11380
rect 42823 11261 42847 11358
rect 42945 11261 42968 11358
rect 42823 11236 42968 11261
rect 34683 10977 34828 10999
rect 34683 10880 34707 10977
rect 34805 10880 34828 10977
rect 34683 10855 34828 10880
rect 35053 10977 35198 10999
rect 35053 10880 35077 10977
rect 35175 10880 35198 10977
rect 35053 10855 35198 10880
rect 35423 10977 35568 10999
rect 35423 10880 35447 10977
rect 35545 10880 35568 10977
rect 35423 10855 35568 10880
rect 35793 10977 35938 10999
rect 35793 10880 35817 10977
rect 35915 10880 35938 10977
rect 35793 10855 35938 10880
rect 36163 10977 36308 10999
rect 36163 10880 36187 10977
rect 36285 10880 36308 10977
rect 36163 10855 36308 10880
rect 36533 10977 36678 10999
rect 36533 10880 36557 10977
rect 36655 10880 36678 10977
rect 36533 10855 36678 10880
rect 36903 10977 37048 10999
rect 36903 10880 36927 10977
rect 37025 10880 37048 10977
rect 36903 10855 37048 10880
rect 37273 10977 37418 10999
rect 37273 10880 37297 10977
rect 37395 10880 37418 10977
rect 37273 10855 37418 10880
rect 37643 10977 37788 10999
rect 37643 10880 37667 10977
rect 37765 10880 37788 10977
rect 37643 10855 37788 10880
rect 38013 10977 38158 10999
rect 38013 10880 38037 10977
rect 38135 10880 38158 10977
rect 38013 10855 38158 10880
rect 38383 10977 38528 10999
rect 38383 10880 38407 10977
rect 38505 10880 38528 10977
rect 38383 10855 38528 10880
rect 38753 10977 38898 10999
rect 38753 10880 38777 10977
rect 38875 10880 38898 10977
rect 38753 10855 38898 10880
rect 39123 10977 39268 10999
rect 39123 10880 39147 10977
rect 39245 10880 39268 10977
rect 39123 10855 39268 10880
rect 39493 10977 39638 10999
rect 39493 10880 39517 10977
rect 39615 10880 39638 10977
rect 39493 10855 39638 10880
rect 39863 10977 40008 10999
rect 39863 10880 39887 10977
rect 39985 10880 40008 10977
rect 39863 10855 40008 10880
rect 40233 10977 40378 10999
rect 40233 10880 40257 10977
rect 40355 10880 40378 10977
rect 40233 10855 40378 10880
rect 40603 10977 40748 10999
rect 40603 10880 40627 10977
rect 40725 10880 40748 10977
rect 40603 10855 40748 10880
rect 40973 10977 41118 10999
rect 40973 10880 40997 10977
rect 41095 10880 41118 10977
rect 40973 10855 41118 10880
rect 41343 10977 41488 10999
rect 41343 10880 41367 10977
rect 41465 10880 41488 10977
rect 41343 10855 41488 10880
rect 41713 10977 41858 10999
rect 41713 10880 41737 10977
rect 41835 10880 41858 10977
rect 41713 10855 41858 10880
rect 42083 10977 42228 10999
rect 42083 10880 42107 10977
rect 42205 10880 42228 10977
rect 42083 10855 42228 10880
rect 42453 10977 42598 10999
rect 42453 10880 42477 10977
rect 42575 10880 42598 10977
rect 42453 10855 42598 10880
rect 42823 10977 42968 10999
rect 42823 10880 42847 10977
rect 42945 10880 42968 10977
rect 42823 10855 42968 10880
rect 34683 10596 34828 10618
rect 34683 10499 34707 10596
rect 34805 10499 34828 10596
rect 34683 10474 34828 10499
rect 35053 10596 35198 10618
rect 35053 10499 35077 10596
rect 35175 10499 35198 10596
rect 35053 10474 35198 10499
rect 35423 10596 35568 10618
rect 35423 10499 35447 10596
rect 35545 10499 35568 10596
rect 35423 10474 35568 10499
rect 35793 10596 35938 10618
rect 35793 10499 35817 10596
rect 35915 10499 35938 10596
rect 35793 10474 35938 10499
rect 36163 10596 36308 10618
rect 36163 10499 36187 10596
rect 36285 10499 36308 10596
rect 36163 10474 36308 10499
rect 36533 10596 36678 10618
rect 36533 10499 36557 10596
rect 36655 10499 36678 10596
rect 36533 10474 36678 10499
rect 36903 10596 37048 10618
rect 36903 10499 36927 10596
rect 37025 10499 37048 10596
rect 36903 10474 37048 10499
rect 37273 10596 37418 10618
rect 37273 10499 37297 10596
rect 37395 10499 37418 10596
rect 37273 10474 37418 10499
rect 37643 10596 37788 10618
rect 37643 10499 37667 10596
rect 37765 10499 37788 10596
rect 37643 10474 37788 10499
rect 38013 10596 38158 10618
rect 38013 10499 38037 10596
rect 38135 10499 38158 10596
rect 38013 10474 38158 10499
rect 38383 10596 38528 10618
rect 38383 10499 38407 10596
rect 38505 10499 38528 10596
rect 38383 10474 38528 10499
rect 38753 10596 38898 10618
rect 38753 10499 38777 10596
rect 38875 10499 38898 10596
rect 38753 10474 38898 10499
rect 39123 10596 39268 10618
rect 39123 10499 39147 10596
rect 39245 10499 39268 10596
rect 39123 10474 39268 10499
rect 39493 10596 39638 10618
rect 39493 10499 39517 10596
rect 39615 10499 39638 10596
rect 39493 10474 39638 10499
rect 39863 10596 40008 10618
rect 39863 10499 39887 10596
rect 39985 10499 40008 10596
rect 39863 10474 40008 10499
rect 40233 10596 40378 10618
rect 40233 10499 40257 10596
rect 40355 10499 40378 10596
rect 40233 10474 40378 10499
rect 40603 10596 40748 10618
rect 40603 10499 40627 10596
rect 40725 10499 40748 10596
rect 40603 10474 40748 10499
rect 40973 10596 41118 10618
rect 40973 10499 40997 10596
rect 41095 10499 41118 10596
rect 40973 10474 41118 10499
rect 41343 10596 41488 10618
rect 41343 10499 41367 10596
rect 41465 10499 41488 10596
rect 41343 10474 41488 10499
rect 41713 10596 41858 10618
rect 41713 10499 41737 10596
rect 41835 10499 41858 10596
rect 41713 10474 41858 10499
rect 42083 10596 42228 10618
rect 42083 10499 42107 10596
rect 42205 10499 42228 10596
rect 42083 10474 42228 10499
rect 42453 10596 42598 10618
rect 42453 10499 42477 10596
rect 42575 10499 42598 10596
rect 42453 10474 42598 10499
rect 42823 10596 42968 10618
rect 42823 10499 42847 10596
rect 42945 10499 42968 10596
rect 42823 10474 42968 10499
<< psubdiffcont >>
rect 21576 -23024 21729 -22872
rect 21861 -23024 22014 -22872
rect 22146 -23024 22299 -22872
rect 22431 -23024 22584 -22872
rect 22716 -23024 22869 -22872
rect 23001 -23024 23154 -22872
rect 23286 -23024 23439 -22872
rect 23571 -23024 23724 -22872
rect 23856 -23024 24009 -22872
rect 24141 -23024 24294 -22872
rect 24426 -23024 24579 -22872
rect 24711 -23024 24864 -22872
rect 24996 -23024 25149 -22872
rect 25281 -23024 25434 -22872
rect 25566 -23024 25719 -22872
rect 25851 -23024 26004 -22872
rect 26136 -23024 26289 -22872
rect 26421 -23024 26574 -22872
rect 26706 -23024 26859 -22872
rect 26991 -23024 27144 -22872
rect 27276 -23024 27429 -22872
rect 27561 -23024 27714 -22872
rect 27846 -23024 27999 -22872
rect 28131 -23024 28284 -22872
rect 28416 -23024 28569 -22872
rect 28701 -23024 28854 -22872
rect 28986 -23024 29139 -22872
rect 29271 -23024 29424 -22872
rect 29556 -23024 29709 -22872
rect 29841 -23024 29994 -22872
rect 30126 -23024 30279 -22872
rect 30411 -23024 30564 -22872
rect 30696 -23024 30849 -22872
rect 30981 -23024 31134 -22872
rect 31266 -23024 31419 -22872
rect 31551 -23024 31704 -22872
rect 31836 -23024 31989 -22872
rect 32121 -23024 32274 -22872
rect 32406 -23024 32559 -22872
rect 32691 -23024 32844 -22872
rect 32976 -23024 33129 -22872
rect 33261 -23024 33414 -22872
rect 33546 -23024 33699 -22872
rect 33831 -23024 33984 -22872
rect 34116 -23024 34269 -22872
rect 34401 -23024 34554 -22872
rect 34686 -23024 34839 -22872
rect 34971 -23024 35124 -22872
rect 35256 -23024 35409 -22872
rect 35541 -23024 35694 -22872
rect 35826 -23024 35979 -22872
rect 36111 -23024 36264 -22872
rect 36396 -23024 36549 -22872
rect 36681 -23024 36834 -22872
rect 36966 -23024 37119 -22872
rect 37251 -23024 37404 -22872
rect 37536 -23024 37689 -22872
rect 37821 -23024 37974 -22872
rect 38106 -23024 38259 -22872
rect 38391 -23024 38544 -22872
rect 38676 -23024 38829 -22872
rect 38961 -23024 39114 -22872
rect 39246 -23024 39399 -22872
rect 39531 -23024 39684 -22872
rect 39816 -23024 39969 -22872
rect 40101 -23024 40254 -22872
rect 40386 -23024 40539 -22872
rect 40671 -23024 40824 -22872
rect 40956 -23024 41109 -22872
rect 41241 -23024 41394 -22872
rect 41526 -23024 41679 -22872
rect 41811 -23024 41964 -22872
rect 42096 -23024 42249 -22872
rect 42381 -23024 42534 -22872
rect 42666 -23024 42819 -22872
rect 42951 -23024 43104 -22872
rect 43236 -23024 43389 -22872
rect 43521 -23024 43674 -22872
rect 43806 -23024 43959 -22872
rect 44091 -23024 44244 -22872
rect 44376 -23024 44529 -22872
rect 44661 -23024 44814 -22872
rect 44946 -23024 45099 -22872
rect 45231 -23024 45384 -22872
rect 45516 -23024 45669 -22872
rect 45801 -23024 45954 -22872
rect 46086 -23024 46239 -22872
rect 46371 -23024 46524 -22872
rect 46656 -23024 46809 -22872
rect 46941 -23024 47094 -22872
rect 47226 -23024 47379 -22872
rect 47511 -23024 47664 -22872
rect 47796 -23024 47949 -22872
rect 48081 -23024 48234 -22872
rect 48366 -23024 48519 -22872
rect 48651 -23024 48804 -22872
rect 48936 -23024 49089 -22872
rect 49221 -23024 49374 -22872
rect 49506 -23024 49659 -22872
rect 49791 -23024 49944 -22872
rect 50076 -23024 50229 -22872
rect 50361 -23024 50514 -22872
rect 50646 -23024 50799 -22872
rect 50931 -23024 51084 -22872
rect 51216 -23024 51369 -22872
rect 51501 -23024 51654 -22872
rect 51786 -23024 51939 -22872
rect 52071 -23024 52224 -22872
rect 52356 -23024 52509 -22872
rect 52641 -23024 52794 -22872
rect 52926 -23024 53079 -22872
rect 53211 -23024 53364 -22872
rect 53496 -23024 53649 -22872
rect 53781 -23024 53934 -22872
rect 54066 -23024 54219 -22872
rect 54351 -23024 54504 -22872
rect 54636 -23024 54789 -22872
rect 54921 -23024 55074 -22872
rect 55206 -23024 55359 -22872
rect 55491 -23024 55644 -22872
rect 55776 -23024 55929 -22872
rect 21576 -23297 21729 -23145
rect 21861 -23297 22014 -23145
rect 22146 -23297 22299 -23145
rect 22431 -23297 22584 -23145
rect 22716 -23297 22869 -23145
rect 23001 -23297 23154 -23145
rect 23286 -23297 23439 -23145
rect 23571 -23297 23724 -23145
rect 23856 -23297 24009 -23145
rect 24141 -23297 24294 -23145
rect 24426 -23297 24579 -23145
rect 24711 -23297 24864 -23145
rect 24996 -23297 25149 -23145
rect 25281 -23297 25434 -23145
rect 25566 -23297 25719 -23145
rect 25851 -23297 26004 -23145
rect 26136 -23297 26289 -23145
rect 26421 -23297 26574 -23145
rect 26706 -23297 26859 -23145
rect 26991 -23297 27144 -23145
rect 27276 -23297 27429 -23145
rect 27561 -23297 27714 -23145
rect 27846 -23297 27999 -23145
rect 28131 -23297 28284 -23145
rect 28416 -23297 28569 -23145
rect 28701 -23297 28854 -23145
rect 28986 -23297 29139 -23145
rect 29271 -23297 29424 -23145
rect 29556 -23297 29709 -23145
rect 29841 -23297 29994 -23145
rect 30126 -23297 30279 -23145
rect 30411 -23297 30564 -23145
rect 30696 -23297 30849 -23145
rect 30981 -23297 31134 -23145
rect 31266 -23297 31419 -23145
rect 31551 -23297 31704 -23145
rect 31836 -23297 31989 -23145
rect 32121 -23297 32274 -23145
rect 32406 -23297 32559 -23145
rect 32691 -23297 32844 -23145
rect 32976 -23297 33129 -23145
rect 33261 -23297 33414 -23145
rect 33546 -23297 33699 -23145
rect 33831 -23297 33984 -23145
rect 34116 -23297 34269 -23145
rect 34401 -23297 34554 -23145
rect 34686 -23297 34839 -23145
rect 34971 -23297 35124 -23145
rect 35256 -23297 35409 -23145
rect 35541 -23297 35694 -23145
rect 35826 -23297 35979 -23145
rect 36111 -23297 36264 -23145
rect 36396 -23297 36549 -23145
rect 36681 -23297 36834 -23145
rect 36966 -23297 37119 -23145
rect 37251 -23297 37404 -23145
rect 37536 -23297 37689 -23145
rect 37821 -23297 37974 -23145
rect 38106 -23297 38259 -23145
rect 38391 -23297 38544 -23145
rect 38676 -23297 38829 -23145
rect 38961 -23297 39114 -23145
rect 39246 -23297 39399 -23145
rect 39531 -23297 39684 -23145
rect 39816 -23297 39969 -23145
rect 40101 -23297 40254 -23145
rect 40386 -23297 40539 -23145
rect 40671 -23297 40824 -23145
rect 40956 -23297 41109 -23145
rect 41241 -23297 41394 -23145
rect 41526 -23297 41679 -23145
rect 41811 -23297 41964 -23145
rect 42096 -23297 42249 -23145
rect 42381 -23297 42534 -23145
rect 42666 -23297 42819 -23145
rect 42951 -23297 43104 -23145
rect 43236 -23297 43389 -23145
rect 43521 -23297 43674 -23145
rect 43806 -23297 43959 -23145
rect 44091 -23297 44244 -23145
rect 44376 -23297 44529 -23145
rect 44661 -23297 44814 -23145
rect 44946 -23297 45099 -23145
rect 45231 -23297 45384 -23145
rect 45516 -23297 45669 -23145
rect 45801 -23297 45954 -23145
rect 46086 -23297 46239 -23145
rect 46371 -23297 46524 -23145
rect 46656 -23297 46809 -23145
rect 46941 -23297 47094 -23145
rect 47226 -23297 47379 -23145
rect 47511 -23297 47664 -23145
rect 47796 -23297 47949 -23145
rect 48081 -23297 48234 -23145
rect 48366 -23297 48519 -23145
rect 48651 -23297 48804 -23145
rect 48936 -23297 49089 -23145
rect 49221 -23297 49374 -23145
rect 49506 -23297 49659 -23145
rect 49791 -23297 49944 -23145
rect 50076 -23297 50229 -23145
rect 50361 -23297 50514 -23145
rect 50646 -23297 50799 -23145
rect 50931 -23297 51084 -23145
rect 51216 -23297 51369 -23145
rect 51501 -23297 51654 -23145
rect 51786 -23297 51939 -23145
rect 52071 -23297 52224 -23145
rect 52356 -23297 52509 -23145
rect 52641 -23297 52794 -23145
rect 52926 -23297 53079 -23145
rect 53211 -23297 53364 -23145
rect 53496 -23297 53649 -23145
rect 53781 -23297 53934 -23145
rect 54066 -23297 54219 -23145
rect 54351 -23297 54504 -23145
rect 54636 -23297 54789 -23145
rect 54921 -23297 55074 -23145
rect 55206 -23297 55359 -23145
rect 55491 -23297 55644 -23145
rect 55776 -23297 55929 -23145
rect 21576 -23570 21729 -23418
rect 21861 -23570 22014 -23418
rect 22146 -23570 22299 -23418
rect 22431 -23570 22584 -23418
rect 22716 -23570 22869 -23418
rect 23001 -23570 23154 -23418
rect 23286 -23570 23439 -23418
rect 23571 -23570 23724 -23418
rect 23856 -23570 24009 -23418
rect 24141 -23570 24294 -23418
rect 24426 -23570 24579 -23418
rect 24711 -23570 24864 -23418
rect 24996 -23570 25149 -23418
rect 25281 -23570 25434 -23418
rect 25566 -23570 25719 -23418
rect 25851 -23570 26004 -23418
rect 26136 -23570 26289 -23418
rect 26421 -23570 26574 -23418
rect 26706 -23570 26859 -23418
rect 26991 -23570 27144 -23418
rect 27276 -23570 27429 -23418
rect 27561 -23570 27714 -23418
rect 27846 -23570 27999 -23418
rect 28131 -23570 28284 -23418
rect 28416 -23570 28569 -23418
rect 28701 -23570 28854 -23418
rect 28986 -23570 29139 -23418
rect 29271 -23570 29424 -23418
rect 29556 -23570 29709 -23418
rect 29841 -23570 29994 -23418
rect 30126 -23570 30279 -23418
rect 30411 -23570 30564 -23418
rect 30696 -23570 30849 -23418
rect 30981 -23570 31134 -23418
rect 31266 -23570 31419 -23418
rect 31551 -23570 31704 -23418
rect 31836 -23570 31989 -23418
rect 32121 -23570 32274 -23418
rect 32406 -23570 32559 -23418
rect 32691 -23570 32844 -23418
rect 32976 -23570 33129 -23418
rect 33261 -23570 33414 -23418
rect 33546 -23570 33699 -23418
rect 33831 -23570 33984 -23418
rect 34116 -23570 34269 -23418
rect 34401 -23570 34554 -23418
rect 34686 -23570 34839 -23418
rect 34971 -23570 35124 -23418
rect 35256 -23570 35409 -23418
rect 35541 -23570 35694 -23418
rect 35826 -23570 35979 -23418
rect 36111 -23570 36264 -23418
rect 36396 -23570 36549 -23418
rect 36681 -23570 36834 -23418
rect 36966 -23570 37119 -23418
rect 37251 -23570 37404 -23418
rect 37536 -23570 37689 -23418
rect 37821 -23570 37974 -23418
rect 38106 -23570 38259 -23418
rect 38391 -23570 38544 -23418
rect 38676 -23570 38829 -23418
rect 38961 -23570 39114 -23418
rect 39246 -23570 39399 -23418
rect 39531 -23570 39684 -23418
rect 39816 -23570 39969 -23418
rect 40101 -23570 40254 -23418
rect 40386 -23570 40539 -23418
rect 40671 -23570 40824 -23418
rect 40956 -23570 41109 -23418
rect 41241 -23570 41394 -23418
rect 41526 -23570 41679 -23418
rect 41811 -23570 41964 -23418
rect 42096 -23570 42249 -23418
rect 42381 -23570 42534 -23418
rect 42666 -23570 42819 -23418
rect 42951 -23570 43104 -23418
rect 43236 -23570 43389 -23418
rect 43521 -23570 43674 -23418
rect 43806 -23570 43959 -23418
rect 44091 -23570 44244 -23418
rect 44376 -23570 44529 -23418
rect 44661 -23570 44814 -23418
rect 44946 -23570 45099 -23418
rect 45231 -23570 45384 -23418
rect 45516 -23570 45669 -23418
rect 45801 -23570 45954 -23418
rect 46086 -23570 46239 -23418
rect 46371 -23570 46524 -23418
rect 46656 -23570 46809 -23418
rect 46941 -23570 47094 -23418
rect 47226 -23570 47379 -23418
rect 47511 -23570 47664 -23418
rect 47796 -23570 47949 -23418
rect 48081 -23570 48234 -23418
rect 48366 -23570 48519 -23418
rect 48651 -23570 48804 -23418
rect 48936 -23570 49089 -23418
rect 49221 -23570 49374 -23418
rect 49506 -23570 49659 -23418
rect 49791 -23570 49944 -23418
rect 50076 -23570 50229 -23418
rect 50361 -23570 50514 -23418
rect 50646 -23570 50799 -23418
rect 50931 -23570 51084 -23418
rect 51216 -23570 51369 -23418
rect 51501 -23570 51654 -23418
rect 51786 -23570 51939 -23418
rect 52071 -23570 52224 -23418
rect 52356 -23570 52509 -23418
rect 52641 -23570 52794 -23418
rect 52926 -23570 53079 -23418
rect 53211 -23570 53364 -23418
rect 53496 -23570 53649 -23418
rect 53781 -23570 53934 -23418
rect 54066 -23570 54219 -23418
rect 54351 -23570 54504 -23418
rect 54636 -23570 54789 -23418
rect 54921 -23570 55074 -23418
rect 55206 -23570 55359 -23418
rect 55491 -23570 55644 -23418
rect 55776 -23570 55929 -23418
rect 21576 -23843 21729 -23691
rect 21861 -23843 22014 -23691
rect 22146 -23843 22299 -23691
rect 22431 -23843 22584 -23691
rect 22716 -23843 22869 -23691
rect 23001 -23843 23154 -23691
rect 23286 -23843 23439 -23691
rect 23571 -23843 23724 -23691
rect 23856 -23843 24009 -23691
rect 24141 -23843 24294 -23691
rect 24426 -23843 24579 -23691
rect 24711 -23843 24864 -23691
rect 24996 -23843 25149 -23691
rect 25281 -23843 25434 -23691
rect 25566 -23843 25719 -23691
rect 25851 -23843 26004 -23691
rect 26136 -23843 26289 -23691
rect 26421 -23843 26574 -23691
rect 26706 -23843 26859 -23691
rect 26991 -23843 27144 -23691
rect 27276 -23843 27429 -23691
rect 27561 -23843 27714 -23691
rect 27846 -23843 27999 -23691
rect 28131 -23843 28284 -23691
rect 28416 -23843 28569 -23691
rect 28701 -23843 28854 -23691
rect 28986 -23843 29139 -23691
rect 29271 -23843 29424 -23691
rect 29556 -23843 29709 -23691
rect 29841 -23843 29994 -23691
rect 30126 -23843 30279 -23691
rect 30411 -23843 30564 -23691
rect 30696 -23843 30849 -23691
rect 30981 -23843 31134 -23691
rect 31266 -23843 31419 -23691
rect 31551 -23843 31704 -23691
rect 31836 -23843 31989 -23691
rect 32121 -23843 32274 -23691
rect 32406 -23843 32559 -23691
rect 32691 -23843 32844 -23691
rect 32976 -23843 33129 -23691
rect 33261 -23843 33414 -23691
rect 33546 -23843 33699 -23691
rect 33831 -23843 33984 -23691
rect 34116 -23843 34269 -23691
rect 34401 -23843 34554 -23691
rect 34686 -23843 34839 -23691
rect 34971 -23843 35124 -23691
rect 35256 -23843 35409 -23691
rect 35541 -23843 35694 -23691
rect 35826 -23843 35979 -23691
rect 36111 -23843 36264 -23691
rect 36396 -23843 36549 -23691
rect 36681 -23843 36834 -23691
rect 36966 -23843 37119 -23691
rect 37251 -23843 37404 -23691
rect 37536 -23843 37689 -23691
rect 37821 -23843 37974 -23691
rect 38106 -23843 38259 -23691
rect 38391 -23843 38544 -23691
rect 38676 -23843 38829 -23691
rect 38961 -23843 39114 -23691
rect 39246 -23843 39399 -23691
rect 39531 -23843 39684 -23691
rect 39816 -23843 39969 -23691
rect 40101 -23843 40254 -23691
rect 40386 -23843 40539 -23691
rect 40671 -23843 40824 -23691
rect 40956 -23843 41109 -23691
rect 41241 -23843 41394 -23691
rect 41526 -23843 41679 -23691
rect 41811 -23843 41964 -23691
rect 42096 -23843 42249 -23691
rect 42381 -23843 42534 -23691
rect 42666 -23843 42819 -23691
rect 42951 -23843 43104 -23691
rect 43236 -23843 43389 -23691
rect 43521 -23843 43674 -23691
rect 43806 -23843 43959 -23691
rect 44091 -23843 44244 -23691
rect 44376 -23843 44529 -23691
rect 44661 -23843 44814 -23691
rect 44946 -23843 45099 -23691
rect 45231 -23843 45384 -23691
rect 45516 -23843 45669 -23691
rect 45801 -23843 45954 -23691
rect 46086 -23843 46239 -23691
rect 46371 -23843 46524 -23691
rect 46656 -23843 46809 -23691
rect 46941 -23843 47094 -23691
rect 47226 -23843 47379 -23691
rect 47511 -23843 47664 -23691
rect 47796 -23843 47949 -23691
rect 48081 -23843 48234 -23691
rect 48366 -23843 48519 -23691
rect 48651 -23843 48804 -23691
rect 48936 -23843 49089 -23691
rect 49221 -23843 49374 -23691
rect 49506 -23843 49659 -23691
rect 49791 -23843 49944 -23691
rect 50076 -23843 50229 -23691
rect 50361 -23843 50514 -23691
rect 50646 -23843 50799 -23691
rect 50931 -23843 51084 -23691
rect 51216 -23843 51369 -23691
rect 51501 -23843 51654 -23691
rect 51786 -23843 51939 -23691
rect 52071 -23843 52224 -23691
rect 52356 -23843 52509 -23691
rect 52641 -23843 52794 -23691
rect 52926 -23843 53079 -23691
rect 53211 -23843 53364 -23691
rect 53496 -23843 53649 -23691
rect 53781 -23843 53934 -23691
rect 54066 -23843 54219 -23691
rect 54351 -23843 54504 -23691
rect 54636 -23843 54789 -23691
rect 54921 -23843 55074 -23691
rect 55206 -23843 55359 -23691
rect 55491 -23843 55644 -23691
rect 55776 -23843 55929 -23691
<< nsubdiffcont >>
rect 34707 11261 34805 11358
rect 35077 11261 35175 11358
rect 35447 11261 35545 11358
rect 35817 11261 35915 11358
rect 36187 11261 36285 11358
rect 36557 11261 36655 11358
rect 36927 11261 37025 11358
rect 37297 11261 37395 11358
rect 37667 11261 37765 11358
rect 38037 11261 38135 11358
rect 38407 11261 38505 11358
rect 38777 11261 38875 11358
rect 39147 11261 39245 11358
rect 39517 11261 39615 11358
rect 39887 11261 39985 11358
rect 40257 11261 40355 11358
rect 40627 11261 40725 11358
rect 40997 11261 41095 11358
rect 41367 11261 41465 11358
rect 41737 11261 41835 11358
rect 42107 11261 42205 11358
rect 42477 11261 42575 11358
rect 42847 11261 42945 11358
rect 34707 10880 34805 10977
rect 35077 10880 35175 10977
rect 35447 10880 35545 10977
rect 35817 10880 35915 10977
rect 36187 10880 36285 10977
rect 36557 10880 36655 10977
rect 36927 10880 37025 10977
rect 37297 10880 37395 10977
rect 37667 10880 37765 10977
rect 38037 10880 38135 10977
rect 38407 10880 38505 10977
rect 38777 10880 38875 10977
rect 39147 10880 39245 10977
rect 39517 10880 39615 10977
rect 39887 10880 39985 10977
rect 40257 10880 40355 10977
rect 40627 10880 40725 10977
rect 40997 10880 41095 10977
rect 41367 10880 41465 10977
rect 41737 10880 41835 10977
rect 42107 10880 42205 10977
rect 42477 10880 42575 10977
rect 42847 10880 42945 10977
rect 34707 10499 34805 10596
rect 35077 10499 35175 10596
rect 35447 10499 35545 10596
rect 35817 10499 35915 10596
rect 36187 10499 36285 10596
rect 36557 10499 36655 10596
rect 36927 10499 37025 10596
rect 37297 10499 37395 10596
rect 37667 10499 37765 10596
rect 38037 10499 38135 10596
rect 38407 10499 38505 10596
rect 38777 10499 38875 10596
rect 39147 10499 39245 10596
rect 39517 10499 39615 10596
rect 39887 10499 39985 10596
rect 40257 10499 40355 10596
rect 40627 10499 40725 10596
rect 40997 10499 41095 10596
rect 41367 10499 41465 10596
rect 41737 10499 41835 10596
rect 42107 10499 42205 10596
rect 42477 10499 42575 10596
rect 42847 10499 42945 10596
<< metal1 >>
rect 41644 12213 42163 12279
rect 34910 12114 35109 12141
rect 34910 11960 34943 12114
rect 35080 11960 35109 12114
rect 34910 11930 35109 11960
rect 35173 12121 35372 12144
rect 35173 11965 35195 12121
rect 35347 11965 35372 12121
rect 35173 11931 35372 11965
rect 35500 12114 35699 12142
rect 35500 11961 35531 12114
rect 35675 11961 35699 12114
rect 35500 11929 35699 11961
rect 41644 11933 41698 12213
rect 42092 11933 42163 12213
rect 41644 11850 42163 11933
rect 34570 11358 43150 11600
rect 17816 11251 18569 11314
rect 17816 10801 17869 11251
rect 18491 10801 18569 11251
rect 17816 10741 18569 10801
rect 18869 11248 19620 11309
rect 18869 10845 18958 11248
rect 19533 10845 19620 11248
rect 18869 10739 19620 10845
rect 34570 11261 34707 11358
rect 34805 11261 35077 11358
rect 35175 11261 35447 11358
rect 35545 11261 35817 11358
rect 35915 11261 36187 11358
rect 36285 11261 36557 11358
rect 36655 11261 36927 11358
rect 37025 11261 37297 11358
rect 37395 11261 37667 11358
rect 37765 11261 38037 11358
rect 38135 11261 38407 11358
rect 38505 11261 38777 11358
rect 38875 11261 39147 11358
rect 39245 11261 39517 11358
rect 39615 11261 39887 11358
rect 39985 11261 40257 11358
rect 40355 11261 40627 11358
rect 40725 11261 40997 11358
rect 41095 11261 41367 11358
rect 41465 11261 41737 11358
rect 41835 11261 42107 11358
rect 42205 11261 42477 11358
rect 42575 11261 42847 11358
rect 42945 11261 43150 11358
rect 34570 10977 43150 11261
rect 34570 10880 34707 10977
rect 34805 10880 35077 10977
rect 35175 10880 35447 10977
rect 35545 10880 35817 10977
rect 35915 10880 36187 10977
rect 36285 10880 36557 10977
rect 36655 10880 36927 10977
rect 37025 10880 37297 10977
rect 37395 10880 37667 10977
rect 37765 10880 38037 10977
rect 38135 10880 38407 10977
rect 38505 10880 38777 10977
rect 38875 10880 39147 10977
rect 39245 10880 39517 10977
rect 39615 10880 39887 10977
rect 39985 10880 40257 10977
rect 40355 10880 40627 10977
rect 40725 10880 40997 10977
rect 41095 10880 41367 10977
rect 41465 10880 41737 10977
rect 41835 10880 42107 10977
rect 42205 10880 42477 10977
rect 42575 10880 42847 10977
rect 42945 10880 43150 10977
rect 34570 10596 43150 10880
rect 34570 10499 34707 10596
rect 34805 10499 35077 10596
rect 35175 10499 35447 10596
rect 35545 10499 35817 10596
rect 35915 10499 36187 10596
rect 36285 10499 36557 10596
rect 36655 10499 36927 10596
rect 37025 10499 37297 10596
rect 37395 10499 37667 10596
rect 37765 10499 38037 10596
rect 38135 10499 38407 10596
rect 38505 10499 38777 10596
rect 38875 10499 39147 10596
rect 39245 10499 39517 10596
rect 39615 10499 39887 10596
rect 39985 10499 40257 10596
rect 40355 10499 40627 10596
rect 40725 10499 40997 10596
rect 41095 10499 41367 10596
rect 41465 10499 41737 10596
rect 41835 10499 42107 10596
rect 42205 10499 42477 10596
rect 42575 10499 42847 10596
rect 42945 10499 43150 10596
rect 34570 10370 43150 10499
rect 34320 9992 34529 10022
rect 34320 9825 34351 9992
rect 34507 9825 34529 9992
rect 34320 9810 34529 9825
rect 33844 8358 34045 8418
rect 33844 8183 33891 8358
rect 34002 8183 34045 8358
rect 33844 8137 34045 8183
rect 36903 7505 37080 10370
rect 37400 7520 37577 10370
rect 37870 7540 38047 10370
rect 38380 7570 38557 10370
rect 38810 7580 38987 10370
rect 39230 7580 39407 10370
rect 39670 7570 39847 10370
rect 40120 7580 40297 10370
rect 38638 7368 38782 7432
rect 34933 7155 35087 7167
rect 34933 7068 34948 7155
rect 35070 7149 35087 7155
rect 35070 7068 35528 7149
rect 34933 7058 35087 7068
rect 36457 7055 36508 7176
rect 37583 7062 37648 7302
rect 38718 7062 38782 7368
rect 39835 7062 39899 7242
rect 33840 6681 35792 6705
rect 33840 6557 35864 6681
rect 33840 6547 35792 6557
rect 43492 6498 43650 6606
rect 35202 6148 35347 6164
rect 35202 6147 35524 6148
rect 35202 6036 35217 6147
rect 35329 6067 35524 6147
rect 35329 6036 35347 6067
rect 35202 6019 35347 6036
rect 36458 5988 36522 6156
rect 37583 5995 37634 6116
rect 38709 5788 38773 6156
rect 39838 5978 39902 6156
rect 57209 5698 57574 5773
rect 41704 5484 42114 5519
rect 39707 5464 39887 5470
rect 41704 5464 41778 5484
rect 39707 5451 41778 5464
rect 39707 5348 39733 5451
rect 39863 5348 41778 5451
rect 39707 5338 41778 5348
rect 42037 5338 42114 5484
rect 39707 5316 42114 5338
rect 39707 5309 39887 5316
rect 41704 5307 42114 5316
rect 57209 5367 57270 5698
rect 57533 5367 57574 5698
rect 34940 5268 38740 5280
rect 57209 5279 57574 5367
rect 34940 5158 34958 5268
rect 35071 5260 38740 5268
rect 35071 5170 38620 5260
rect 38730 5170 38740 5260
rect 35071 5158 38740 5170
rect 34940 5150 38740 5158
rect 41708 5090 42113 5094
rect 41702 5053 42113 5090
rect 41702 5009 41757 5053
rect 33758 4795 41757 5009
rect 42024 5009 42113 5053
rect 42024 4795 45064 5009
rect 33758 4728 45064 4795
rect 41702 4717 42113 4728
rect 41708 4689 42113 4717
rect 42708 4265 43121 4516
rect 32588 3449 33088 3505
rect 37815 3449 38032 3471
rect 32588 3415 38032 3449
rect 32588 3397 37856 3415
rect 32588 3159 32655 3397
rect 32948 3247 37856 3397
rect 38001 3247 38032 3415
rect 32948 3202 38032 3247
rect 32948 3159 33088 3202
rect 37815 3171 38032 3202
rect 32588 3048 33088 3159
rect 19154 2873 19426 2933
rect 19154 2716 19196 2873
rect 19360 2716 19426 2873
rect 42201 2792 42374 2793
rect 42199 2782 42377 2792
rect 42199 2780 42213 2782
rect 19154 2679 19426 2716
rect 34551 2763 42213 2780
rect 34551 2622 34562 2763
rect 34665 2622 42213 2763
rect 34551 2603 42213 2622
rect 42369 2603 42377 2782
rect 34551 2601 42377 2603
rect 42199 2591 42377 2601
rect 34731 2456 34935 2492
rect 41460 2456 41640 2470
rect 34731 2455 41640 2456
rect 33824 2330 34082 2367
rect 30436 2124 33880 2330
rect 34068 2124 34082 2330
rect 34731 2297 34759 2455
rect 34905 2450 41640 2455
rect 34905 2297 41480 2450
rect 34731 2280 41480 2297
rect 41630 2280 41640 2450
rect 34731 2272 41640 2280
rect 34731 2262 34935 2272
rect 41460 2250 41640 2272
rect 30436 2093 34082 2124
rect 33824 2062 34082 2093
rect 43378 2178 43473 2203
rect 43378 2098 43396 2178
rect 43457 2098 43473 2178
rect 43378 2071 43473 2098
rect 35185 2027 35372 2044
rect 37477 2027 37606 2030
rect 35185 2024 37606 2027
rect 35185 1899 35214 2024
rect 35346 2008 37606 2024
rect 35346 1902 37502 2008
rect 37585 1902 37606 2008
rect 35346 1899 37606 1902
rect 35185 1895 37606 1899
rect 35185 1872 35372 1895
rect 37477 1881 37606 1895
rect 28028 1821 28258 1856
rect 28028 1665 28065 1821
rect 28228 1665 28258 1821
rect 28028 1630 28258 1665
rect 33883 1660 34022 1666
rect 30611 1647 34022 1660
rect 30611 1630 33894 1647
rect 30605 1572 33894 1630
rect 30611 1541 33894 1572
rect 34008 1541 34022 1647
rect 30611 1532 34022 1541
rect 33883 1531 34022 1532
rect 34550 1175 34672 1193
rect 34550 1088 34564 1175
rect 34662 1137 34672 1175
rect 39734 1167 39882 1185
rect 39734 1157 39754 1167
rect 34662 1090 35116 1137
rect 36204 1134 36286 1146
rect 34662 1088 34672 1090
rect 34550 1068 34672 1088
rect 36204 1075 36213 1134
rect 36273 1075 36286 1134
rect 39485 1123 39754 1157
rect 36204 1066 36286 1075
rect 39307 1068 39754 1123
rect 39485 1051 39754 1068
rect 39734 1037 39754 1051
rect 39872 1037 39882 1167
rect 39734 1018 39882 1037
rect 41742 797 42116 892
rect 41742 758 41837 797
rect 39320 675 41837 758
rect 39289 515 41837 675
rect 41742 480 41837 515
rect 42106 480 42116 797
rect 43366 544 43458 551
rect 43366 488 43380 544
rect 43440 488 43458 544
rect 43366 482 43458 488
rect 41742 417 42116 480
rect 37238 271 37329 284
rect 37238 213 37251 271
rect 37308 213 37329 271
rect 37238 197 37329 213
rect 37252 75 37309 197
rect 37113 18 37309 75
rect 34767 -1892 34909 -1880
rect 34767 -2000 34780 -1892
rect 34897 -1912 34909 -1892
rect 34897 -1996 35159 -1912
rect 36196 -1929 36287 -1916
rect 36196 -1992 36210 -1929
rect 36276 -1992 36287 -1929
rect 34897 -2000 34909 -1996
rect 34767 -2017 34909 -2000
rect 36196 -2004 36287 -1992
rect 41701 -2990 42314 -2932
rect 41701 -3053 41771 -2990
rect 30721 -3242 41771 -3053
rect 42236 -3053 42314 -2990
rect 45023 -3053 45212 -2394
rect 42236 -3242 45212 -3053
rect 41701 -3316 42314 -3242
rect 18971 -4176 19435 -3950
rect 18971 -4572 19061 -4176
rect 19310 -4572 19435 -4176
rect 57240 -4138 57627 -3991
rect 18971 -4719 19435 -4572
rect 42454 -4299 42680 -4298
rect 42454 -4352 43394 -4299
rect 42454 -4605 42485 -4352
rect 42645 -4605 43394 -4352
rect 42454 -4632 43394 -4605
rect 57240 -4593 57314 -4138
rect 57541 -4593 57627 -4138
rect 42454 -4656 42680 -4632
rect 57240 -4718 57627 -4593
rect 34226 -4954 34596 -4895
rect 34226 -5168 34281 -4954
rect 34547 -5168 34596 -4954
rect 34226 -5220 34596 -5168
rect 34768 -5556 34931 -5539
rect 42328 -5549 42544 -5529
rect 42328 -5556 42348 -5549
rect 34768 -5560 42348 -5556
rect 34768 -5708 34788 -5560
rect 34910 -5708 42348 -5560
rect 34768 -5722 42348 -5708
rect 42526 -5722 42544 -5549
rect 34768 -5732 42544 -5722
rect 42328 -5756 42544 -5732
rect 42326 -7564 42560 -7540
rect 42326 -7604 42354 -7564
rect 19088 -7739 19417 -7703
rect 41311 -7728 42354 -7604
rect 42530 -7728 42560 -7564
rect 41311 -7734 42560 -7728
rect 19088 -8019 19119 -7739
rect 19368 -8019 19417 -7739
rect 42326 -7750 42560 -7734
rect 19088 -8079 19417 -8019
rect 55478 -8641 55756 -8589
rect 55478 -8825 55513 -8641
rect 55696 -8825 55756 -8641
rect 55478 -8880 55756 -8825
rect 57244 -9679 57490 -9673
rect 57211 -9746 57563 -9679
rect 57211 -10038 57251 -9746
rect 57457 -10038 57563 -9746
rect 57211 -10104 57563 -10038
rect 41438 -10171 42929 -10127
rect 41438 -10421 41745 -10171
rect 42266 -10421 42929 -10171
rect 41438 -10472 42929 -10421
rect 19826 -12000 21571 -11979
rect 19804 -12058 21571 -12000
rect 19804 -12310 19869 -12058
rect 20071 -12310 21571 -12058
rect 19804 -12397 21571 -12310
rect 19826 -12404 21571 -12397
rect 41273 -12235 41674 -12161
rect 41273 -12413 41335 -12235
rect 41604 -12413 41674 -12235
rect 41273 -12454 41674 -12413
rect 35138 -12875 35375 -12834
rect 35138 -12881 35169 -12875
rect 34924 -13041 35169 -12881
rect 35138 -13044 35169 -13041
rect 35348 -13044 35375 -12875
rect 35138 -13077 35375 -13044
rect 37211 -14965 40395 -14903
rect 37211 -15247 38672 -14965
rect 39016 -15247 40395 -14965
rect 37211 -15309 40395 -15247
rect 57220 -16173 57646 -16072
rect 57220 -16547 57289 -16173
rect 57564 -16547 57646 -16173
rect 57220 -16623 57646 -16547
rect 19108 -17013 19454 -16917
rect 19108 -17206 19180 -17013
rect 19363 -17206 19454 -17013
rect 19108 -17290 19454 -17206
rect 36001 -18806 36246 -18777
rect 36001 -19007 36043 -18806
rect 36207 -19007 36246 -18806
rect 36001 -19062 36246 -19007
rect 56390 -19738 56703 -19713
rect 56390 -19819 56421 -19738
rect 55676 -19888 56421 -19819
rect 56390 -19908 56421 -19888
rect 56676 -19908 56703 -19738
rect 56390 -19946 56703 -19908
rect 21421 -22872 56289 -22738
rect 21421 -23024 21576 -22872
rect 21729 -23024 21861 -22872
rect 22014 -23024 22146 -22872
rect 22299 -23024 22431 -22872
rect 22584 -23024 22716 -22872
rect 22869 -23024 23001 -22872
rect 23154 -23024 23286 -22872
rect 23439 -23024 23571 -22872
rect 23724 -23024 23856 -22872
rect 24009 -23024 24141 -22872
rect 24294 -23024 24426 -22872
rect 24579 -23024 24711 -22872
rect 24864 -23024 24996 -22872
rect 25149 -23024 25281 -22872
rect 25434 -23024 25566 -22872
rect 25719 -23024 25851 -22872
rect 26004 -23024 26136 -22872
rect 26289 -23024 26421 -22872
rect 26574 -23024 26706 -22872
rect 26859 -23024 26991 -22872
rect 27144 -23024 27276 -22872
rect 27429 -23024 27561 -22872
rect 27714 -23024 27846 -22872
rect 27999 -23024 28131 -22872
rect 28284 -23024 28416 -22872
rect 28569 -23024 28701 -22872
rect 28854 -23024 28986 -22872
rect 29139 -23024 29271 -22872
rect 29424 -23024 29556 -22872
rect 29709 -23024 29841 -22872
rect 29994 -23024 30126 -22872
rect 30279 -23024 30411 -22872
rect 30564 -23024 30696 -22872
rect 30849 -23024 30981 -22872
rect 31134 -23024 31266 -22872
rect 31419 -23024 31551 -22872
rect 31704 -23024 31836 -22872
rect 31989 -23024 32121 -22872
rect 32274 -23024 32406 -22872
rect 32559 -23024 32691 -22872
rect 32844 -23024 32976 -22872
rect 33129 -23024 33261 -22872
rect 33414 -23024 33546 -22872
rect 33699 -23024 33831 -22872
rect 33984 -23024 34116 -22872
rect 34269 -23024 34401 -22872
rect 34554 -23024 34686 -22872
rect 34839 -23024 34971 -22872
rect 35124 -23024 35256 -22872
rect 35409 -23024 35541 -22872
rect 35694 -23024 35826 -22872
rect 35979 -23024 36111 -22872
rect 36264 -23024 36396 -22872
rect 36549 -23024 36681 -22872
rect 36834 -23024 36966 -22872
rect 37119 -23024 37251 -22872
rect 37404 -23024 37536 -22872
rect 37689 -23024 37821 -22872
rect 37974 -23024 38106 -22872
rect 38259 -23024 38391 -22872
rect 38544 -23024 38676 -22872
rect 38829 -23024 38961 -22872
rect 39114 -23024 39246 -22872
rect 39399 -23024 39531 -22872
rect 39684 -23024 39816 -22872
rect 39969 -23024 40101 -22872
rect 40254 -23024 40386 -22872
rect 40539 -23024 40671 -22872
rect 40824 -23024 40956 -22872
rect 41109 -23024 41241 -22872
rect 41394 -23024 41526 -22872
rect 41679 -23024 41811 -22872
rect 41964 -23024 42096 -22872
rect 42249 -23024 42381 -22872
rect 42534 -23024 42666 -22872
rect 42819 -23024 42951 -22872
rect 43104 -23024 43236 -22872
rect 43389 -23024 43521 -22872
rect 43674 -23024 43806 -22872
rect 43959 -23024 44091 -22872
rect 44244 -23024 44376 -22872
rect 44529 -23024 44661 -22872
rect 44814 -23024 44946 -22872
rect 45099 -23024 45231 -22872
rect 45384 -23024 45516 -22872
rect 45669 -23024 45801 -22872
rect 45954 -23024 46086 -22872
rect 46239 -23024 46371 -22872
rect 46524 -23024 46656 -22872
rect 46809 -23024 46941 -22872
rect 47094 -23024 47226 -22872
rect 47379 -23024 47511 -22872
rect 47664 -23024 47796 -22872
rect 47949 -23024 48081 -22872
rect 48234 -23024 48366 -22872
rect 48519 -23024 48651 -22872
rect 48804 -23024 48936 -22872
rect 49089 -23024 49221 -22872
rect 49374 -23024 49506 -22872
rect 49659 -23024 49791 -22872
rect 49944 -23024 50076 -22872
rect 50229 -23024 50361 -22872
rect 50514 -23024 50646 -22872
rect 50799 -23024 50931 -22872
rect 51084 -23024 51216 -22872
rect 51369 -23024 51501 -22872
rect 51654 -23024 51786 -22872
rect 51939 -23024 52071 -22872
rect 52224 -23024 52356 -22872
rect 52509 -23024 52641 -22872
rect 52794 -23024 52926 -22872
rect 53079 -23024 53211 -22872
rect 53364 -23024 53496 -22872
rect 53649 -23024 53781 -22872
rect 53934 -23024 54066 -22872
rect 54219 -23024 54351 -22872
rect 54504 -23024 54636 -22872
rect 54789 -23024 54921 -22872
rect 55074 -23024 55206 -22872
rect 55359 -23024 55491 -22872
rect 55644 -23024 55776 -22872
rect 55929 -23024 56289 -22872
rect 21421 -23059 56289 -23024
rect 21421 -23145 38572 -23059
rect 39145 -23145 56289 -23059
rect 21421 -23297 21576 -23145
rect 21729 -23297 21861 -23145
rect 22014 -23297 22146 -23145
rect 22299 -23297 22431 -23145
rect 22584 -23297 22716 -23145
rect 22869 -23297 23001 -23145
rect 23154 -23297 23286 -23145
rect 23439 -23297 23571 -23145
rect 23724 -23297 23856 -23145
rect 24009 -23297 24141 -23145
rect 24294 -23297 24426 -23145
rect 24579 -23297 24711 -23145
rect 24864 -23297 24996 -23145
rect 25149 -23297 25281 -23145
rect 25434 -23297 25566 -23145
rect 25719 -23297 25851 -23145
rect 26004 -23297 26136 -23145
rect 26289 -23297 26421 -23145
rect 26574 -23297 26706 -23145
rect 26859 -23297 26991 -23145
rect 27144 -23297 27276 -23145
rect 27429 -23297 27561 -23145
rect 27714 -23297 27846 -23145
rect 27999 -23297 28131 -23145
rect 28284 -23297 28416 -23145
rect 28569 -23297 28701 -23145
rect 28854 -23297 28986 -23145
rect 29139 -23297 29271 -23145
rect 29424 -23297 29556 -23145
rect 29709 -23297 29841 -23145
rect 29994 -23297 30126 -23145
rect 30279 -23297 30411 -23145
rect 30564 -23297 30696 -23145
rect 30849 -23297 30981 -23145
rect 31134 -23297 31266 -23145
rect 31419 -23297 31551 -23145
rect 31704 -23297 31836 -23145
rect 31989 -23297 32121 -23145
rect 32274 -23297 32406 -23145
rect 32559 -23297 32691 -23145
rect 32844 -23297 32976 -23145
rect 33129 -23297 33261 -23145
rect 33414 -23297 33546 -23145
rect 33699 -23297 33831 -23145
rect 33984 -23297 34116 -23145
rect 34269 -23297 34401 -23145
rect 34554 -23297 34686 -23145
rect 34839 -23297 34971 -23145
rect 35124 -23297 35256 -23145
rect 35409 -23297 35541 -23145
rect 35694 -23297 35826 -23145
rect 35979 -23297 36111 -23145
rect 36264 -23297 36396 -23145
rect 36549 -23297 36681 -23145
rect 36834 -23297 36966 -23145
rect 37119 -23297 37251 -23145
rect 37404 -23297 37536 -23145
rect 37689 -23297 37821 -23145
rect 37974 -23297 38106 -23145
rect 38259 -23297 38391 -23145
rect 38544 -23297 38572 -23145
rect 39145 -23297 39246 -23145
rect 39399 -23297 39531 -23145
rect 39684 -23297 39816 -23145
rect 39969 -23297 40101 -23145
rect 40254 -23297 40386 -23145
rect 40539 -23297 40671 -23145
rect 40824 -23297 40956 -23145
rect 41109 -23297 41241 -23145
rect 41394 -23297 41526 -23145
rect 41679 -23297 41811 -23145
rect 41964 -23297 42096 -23145
rect 42249 -23297 42381 -23145
rect 42534 -23297 42666 -23145
rect 42819 -23297 42951 -23145
rect 43104 -23297 43236 -23145
rect 43389 -23297 43521 -23145
rect 43674 -23297 43806 -23145
rect 43959 -23297 44091 -23145
rect 44244 -23297 44376 -23145
rect 44529 -23297 44661 -23145
rect 44814 -23297 44946 -23145
rect 45099 -23297 45231 -23145
rect 45384 -23297 45516 -23145
rect 45669 -23297 45801 -23145
rect 45954 -23297 46086 -23145
rect 46239 -23297 46371 -23145
rect 46524 -23297 46656 -23145
rect 46809 -23297 46941 -23145
rect 47094 -23297 47226 -23145
rect 47379 -23297 47511 -23145
rect 47664 -23297 47796 -23145
rect 47949 -23297 48081 -23145
rect 48234 -23297 48366 -23145
rect 48519 -23297 48651 -23145
rect 48804 -23297 48936 -23145
rect 49089 -23297 49221 -23145
rect 49374 -23297 49506 -23145
rect 49659 -23297 49791 -23145
rect 49944 -23297 50076 -23145
rect 50229 -23297 50361 -23145
rect 50514 -23297 50646 -23145
rect 50799 -23297 50931 -23145
rect 51084 -23297 51216 -23145
rect 51369 -23297 51501 -23145
rect 51654 -23297 51786 -23145
rect 51939 -23297 52071 -23145
rect 52224 -23297 52356 -23145
rect 52509 -23297 52641 -23145
rect 52794 -23297 52926 -23145
rect 53079 -23297 53211 -23145
rect 53364 -23297 53496 -23145
rect 53649 -23297 53781 -23145
rect 53934 -23297 54066 -23145
rect 54219 -23297 54351 -23145
rect 54504 -23297 54636 -23145
rect 54789 -23297 54921 -23145
rect 55074 -23297 55206 -23145
rect 55359 -23297 55491 -23145
rect 55644 -23297 55776 -23145
rect 55929 -23297 56289 -23145
rect 21421 -23418 38572 -23297
rect 39145 -23418 56289 -23297
rect 21421 -23570 21576 -23418
rect 21729 -23570 21861 -23418
rect 22014 -23570 22146 -23418
rect 22299 -23570 22431 -23418
rect 22584 -23570 22716 -23418
rect 22869 -23570 23001 -23418
rect 23154 -23570 23286 -23418
rect 23439 -23570 23571 -23418
rect 23724 -23570 23856 -23418
rect 24009 -23570 24141 -23418
rect 24294 -23570 24426 -23418
rect 24579 -23570 24711 -23418
rect 24864 -23570 24996 -23418
rect 25149 -23570 25281 -23418
rect 25434 -23570 25566 -23418
rect 25719 -23570 25851 -23418
rect 26004 -23570 26136 -23418
rect 26289 -23570 26421 -23418
rect 26574 -23570 26706 -23418
rect 26859 -23570 26991 -23418
rect 27144 -23570 27276 -23418
rect 27429 -23570 27561 -23418
rect 27714 -23570 27846 -23418
rect 27999 -23570 28131 -23418
rect 28284 -23570 28416 -23418
rect 28569 -23570 28701 -23418
rect 28854 -23570 28986 -23418
rect 29139 -23570 29271 -23418
rect 29424 -23570 29556 -23418
rect 29709 -23570 29841 -23418
rect 29994 -23570 30126 -23418
rect 30279 -23570 30411 -23418
rect 30564 -23570 30696 -23418
rect 30849 -23570 30981 -23418
rect 31134 -23570 31266 -23418
rect 31419 -23570 31551 -23418
rect 31704 -23570 31836 -23418
rect 31989 -23570 32121 -23418
rect 32274 -23570 32406 -23418
rect 32559 -23570 32691 -23418
rect 32844 -23570 32976 -23418
rect 33129 -23570 33261 -23418
rect 33414 -23570 33546 -23418
rect 33699 -23570 33831 -23418
rect 33984 -23570 34116 -23418
rect 34269 -23570 34401 -23418
rect 34554 -23570 34686 -23418
rect 34839 -23570 34971 -23418
rect 35124 -23570 35256 -23418
rect 35409 -23570 35541 -23418
rect 35694 -23570 35826 -23418
rect 35979 -23570 36111 -23418
rect 36264 -23570 36396 -23418
rect 36549 -23570 36681 -23418
rect 36834 -23570 36966 -23418
rect 37119 -23570 37251 -23418
rect 37404 -23570 37536 -23418
rect 37689 -23570 37821 -23418
rect 37974 -23570 38106 -23418
rect 38259 -23570 38391 -23418
rect 38544 -23526 38572 -23418
rect 39145 -23526 39246 -23418
rect 38544 -23570 38676 -23526
rect 38829 -23570 38961 -23526
rect 39114 -23570 39246 -23526
rect 39399 -23570 39531 -23418
rect 39684 -23570 39816 -23418
rect 39969 -23570 40101 -23418
rect 40254 -23570 40386 -23418
rect 40539 -23570 40671 -23418
rect 40824 -23570 40956 -23418
rect 41109 -23570 41241 -23418
rect 41394 -23570 41526 -23418
rect 41679 -23570 41811 -23418
rect 41964 -23570 42096 -23418
rect 42249 -23570 42381 -23418
rect 42534 -23570 42666 -23418
rect 42819 -23570 42951 -23418
rect 43104 -23570 43236 -23418
rect 43389 -23570 43521 -23418
rect 43674 -23570 43806 -23418
rect 43959 -23570 44091 -23418
rect 44244 -23570 44376 -23418
rect 44529 -23570 44661 -23418
rect 44814 -23570 44946 -23418
rect 45099 -23570 45231 -23418
rect 45384 -23570 45516 -23418
rect 45669 -23570 45801 -23418
rect 45954 -23570 46086 -23418
rect 46239 -23570 46371 -23418
rect 46524 -23570 46656 -23418
rect 46809 -23570 46941 -23418
rect 47094 -23570 47226 -23418
rect 47379 -23570 47511 -23418
rect 47664 -23570 47796 -23418
rect 47949 -23570 48081 -23418
rect 48234 -23570 48366 -23418
rect 48519 -23570 48651 -23418
rect 48804 -23570 48936 -23418
rect 49089 -23570 49221 -23418
rect 49374 -23570 49506 -23418
rect 49659 -23570 49791 -23418
rect 49944 -23570 50076 -23418
rect 50229 -23570 50361 -23418
rect 50514 -23570 50646 -23418
rect 50799 -23570 50931 -23418
rect 51084 -23570 51216 -23418
rect 51369 -23570 51501 -23418
rect 51654 -23570 51786 -23418
rect 51939 -23570 52071 -23418
rect 52224 -23570 52356 -23418
rect 52509 -23570 52641 -23418
rect 52794 -23570 52926 -23418
rect 53079 -23570 53211 -23418
rect 53364 -23570 53496 -23418
rect 53649 -23570 53781 -23418
rect 53934 -23570 54066 -23418
rect 54219 -23570 54351 -23418
rect 54504 -23570 54636 -23418
rect 54789 -23570 54921 -23418
rect 55074 -23570 55206 -23418
rect 55359 -23570 55491 -23418
rect 55644 -23570 55776 -23418
rect 55929 -23570 56289 -23418
rect 21421 -23691 56289 -23570
rect 21421 -23843 21576 -23691
rect 21729 -23843 21861 -23691
rect 22014 -23843 22146 -23691
rect 22299 -23843 22431 -23691
rect 22584 -23843 22716 -23691
rect 22869 -23843 23001 -23691
rect 23154 -23843 23286 -23691
rect 23439 -23843 23571 -23691
rect 23724 -23843 23856 -23691
rect 24009 -23843 24141 -23691
rect 24294 -23843 24426 -23691
rect 24579 -23843 24711 -23691
rect 24864 -23843 24996 -23691
rect 25149 -23843 25281 -23691
rect 25434 -23843 25566 -23691
rect 25719 -23843 25851 -23691
rect 26004 -23843 26136 -23691
rect 26289 -23843 26421 -23691
rect 26574 -23843 26706 -23691
rect 26859 -23843 26991 -23691
rect 27144 -23843 27276 -23691
rect 27429 -23843 27561 -23691
rect 27714 -23843 27846 -23691
rect 27999 -23843 28131 -23691
rect 28284 -23843 28416 -23691
rect 28569 -23843 28701 -23691
rect 28854 -23843 28986 -23691
rect 29139 -23843 29271 -23691
rect 29424 -23843 29556 -23691
rect 29709 -23843 29841 -23691
rect 29994 -23843 30126 -23691
rect 30279 -23843 30411 -23691
rect 30564 -23843 30696 -23691
rect 30849 -23843 30981 -23691
rect 31134 -23843 31266 -23691
rect 31419 -23843 31551 -23691
rect 31704 -23843 31836 -23691
rect 31989 -23843 32121 -23691
rect 32274 -23843 32406 -23691
rect 32559 -23843 32691 -23691
rect 32844 -23843 32976 -23691
rect 33129 -23843 33261 -23691
rect 33414 -23843 33546 -23691
rect 33699 -23843 33831 -23691
rect 33984 -23843 34116 -23691
rect 34269 -23843 34401 -23691
rect 34554 -23843 34686 -23691
rect 34839 -23843 34971 -23691
rect 35124 -23843 35256 -23691
rect 35409 -23843 35541 -23691
rect 35694 -23843 35826 -23691
rect 35979 -23843 36111 -23691
rect 36264 -23843 36396 -23691
rect 36549 -23843 36681 -23691
rect 36834 -23843 36966 -23691
rect 37119 -23843 37251 -23691
rect 37404 -23843 37536 -23691
rect 37689 -23843 37821 -23691
rect 37974 -23843 38106 -23691
rect 38259 -23843 38391 -23691
rect 38544 -23843 38676 -23691
rect 38829 -23843 38961 -23691
rect 39114 -23843 39246 -23691
rect 39399 -23843 39531 -23691
rect 39684 -23843 39816 -23691
rect 39969 -23843 40101 -23691
rect 40254 -23843 40386 -23691
rect 40539 -23843 40671 -23691
rect 40824 -23843 40956 -23691
rect 41109 -23843 41241 -23691
rect 41394 -23843 41526 -23691
rect 41679 -23843 41811 -23691
rect 41964 -23843 42096 -23691
rect 42249 -23843 42381 -23691
rect 42534 -23843 42666 -23691
rect 42819 -23843 42951 -23691
rect 43104 -23843 43236 -23691
rect 43389 -23843 43521 -23691
rect 43674 -23843 43806 -23691
rect 43959 -23843 44091 -23691
rect 44244 -23843 44376 -23691
rect 44529 -23843 44661 -23691
rect 44814 -23843 44946 -23691
rect 45099 -23843 45231 -23691
rect 45384 -23843 45516 -23691
rect 45669 -23843 45801 -23691
rect 45954 -23843 46086 -23691
rect 46239 -23843 46371 -23691
rect 46524 -23843 46656 -23691
rect 46809 -23843 46941 -23691
rect 47094 -23843 47226 -23691
rect 47379 -23843 47511 -23691
rect 47664 -23843 47796 -23691
rect 47949 -23843 48081 -23691
rect 48234 -23843 48366 -23691
rect 48519 -23843 48651 -23691
rect 48804 -23843 48936 -23691
rect 49089 -23843 49221 -23691
rect 49374 -23843 49506 -23691
rect 49659 -23843 49791 -23691
rect 49944 -23843 50076 -23691
rect 50229 -23843 50361 -23691
rect 50514 -23843 50646 -23691
rect 50799 -23843 50931 -23691
rect 51084 -23843 51216 -23691
rect 51369 -23843 51501 -23691
rect 51654 -23843 51786 -23691
rect 51939 -23843 52071 -23691
rect 52224 -23843 52356 -23691
rect 52509 -23843 52641 -23691
rect 52794 -23843 52926 -23691
rect 53079 -23843 53211 -23691
rect 53364 -23843 53496 -23691
rect 53649 -23843 53781 -23691
rect 53934 -23843 54066 -23691
rect 54219 -23843 54351 -23691
rect 54504 -23843 54636 -23691
rect 54789 -23843 54921 -23691
rect 55074 -23843 55206 -23691
rect 55359 -23843 55491 -23691
rect 55644 -23843 55776 -23691
rect 55929 -23843 56289 -23691
rect 21421 -23960 56289 -23843
<< via1 >>
rect 34943 11960 35080 12114
rect 35195 11965 35347 12121
rect 35531 11961 35675 12114
rect 41698 11933 42092 12213
rect 17869 10801 18491 11251
rect 18958 10845 19533 11248
rect 34351 9825 34507 9992
rect 33891 8183 34002 8358
rect 43502 8412 43573 8494
rect 43521 7768 43575 7831
rect 33707 7359 33780 7419
rect 34948 7068 35070 7155
rect 35217 6036 35329 6147
rect 38878 5565 39010 5623
rect 39259 5563 39393 5623
rect 39733 5348 39863 5451
rect 41778 5338 42037 5484
rect 57270 5367 57533 5698
rect 34958 5158 35071 5268
rect 38620 5170 38730 5260
rect 41757 4795 42024 5053
rect 32655 3159 32948 3397
rect 37856 3247 38001 3415
rect 19196 2716 19360 2873
rect 34562 2622 34665 2763
rect 42213 2603 42369 2782
rect 33880 2124 34068 2330
rect 34759 2297 34905 2455
rect 41480 2280 41630 2450
rect 43396 2098 43457 2178
rect 35214 1899 35346 2024
rect 37502 1902 37585 2008
rect 28065 1665 28228 1821
rect 33894 1541 34008 1647
rect 38890 1560 39000 1650
rect 39270 1590 39390 1660
rect 34564 1088 34662 1175
rect 36213 1075 36273 1134
rect 39754 1037 39872 1167
rect 41837 480 42106 797
rect 43380 488 43440 544
rect 37251 213 37308 271
rect 35903 19 35972 73
rect 35902 -926 35975 -873
rect 37032 -927 37108 -874
rect 34780 -2000 34897 -1892
rect 36210 -1992 36276 -1929
rect 41771 -3242 42236 -2990
rect 19061 -4572 19310 -4176
rect 42485 -4605 42645 -4352
rect 57314 -4593 57541 -4138
rect 34281 -5168 34547 -4954
rect 34788 -5708 34910 -5560
rect 42348 -5722 42526 -5549
rect 42354 -7728 42530 -7564
rect 19119 -8019 19368 -7739
rect 55513 -8825 55696 -8641
rect 57251 -10038 57457 -9746
rect 38709 -10438 38970 -10288
rect 41745 -10421 42266 -10171
rect 19869 -12310 20071 -12058
rect 41335 -12413 41604 -12235
rect 35169 -13044 35348 -12875
rect 38672 -15247 39016 -14965
rect 57289 -16547 57564 -16173
rect 19180 -17206 19363 -17013
rect 36043 -19007 36207 -18806
rect 56421 -19908 56676 -19738
rect 38572 -23145 39145 -23059
rect 38572 -23297 38676 -23145
rect 38676 -23297 38829 -23145
rect 38829 -23297 38961 -23145
rect 38961 -23297 39114 -23145
rect 39114 -23297 39145 -23145
rect 38572 -23418 39145 -23297
rect 38572 -23526 38676 -23418
rect 38676 -23526 38829 -23418
rect 38829 -23526 38961 -23418
rect 38961 -23526 39114 -23418
rect 39114 -23526 39145 -23418
<< metal2 >>
rect 41644 12213 42163 12279
rect 34910 12114 35109 12141
rect 34910 11960 34943 12114
rect 35080 11960 35109 12114
rect 34910 11930 35109 11960
rect 35173 12121 35372 12144
rect 35173 11965 35195 12121
rect 35347 11965 35372 12121
rect 35173 11931 35372 11965
rect 35500 12114 35699 12142
rect 35500 11961 35531 12114
rect 35675 11961 35699 12114
rect 17817 11314 18567 11315
rect 17816 11251 18569 11314
rect 17816 10801 17869 11251
rect 18491 10801 18569 11251
rect 17816 10741 18569 10801
rect 18869 11273 19620 11309
rect 18869 11248 19621 11273
rect 18869 10845 18958 11248
rect 19533 10845 19621 11248
rect 17817 4646 18567 10741
rect 18869 10739 19621 10845
rect 17817 4174 18015 4646
rect 18361 4174 18567 4646
rect 17817 -5667 18567 4174
rect 17817 -6036 18068 -5667
rect 18326 -6036 18567 -5667
rect 17817 -21293 18567 -6036
rect 18871 2897 19621 10739
rect 34320 10022 34527 10023
rect 34320 9992 34529 10022
rect 34320 9825 34351 9992
rect 34507 9825 34529 9992
rect 34320 9810 34529 9825
rect 33844 8387 34045 8418
rect 33844 8160 33865 8387
rect 34022 8160 34045 8387
rect 33844 8137 34045 8160
rect 33855 8000 34077 8002
rect 33855 7980 34083 8000
rect 33855 7836 33877 7980
rect 34060 7836 34083 7980
rect 33855 7820 34083 7836
rect 33699 7436 33786 7447
rect 33699 7347 33707 7436
rect 33778 7419 33786 7436
rect 33780 7359 33786 7419
rect 33778 7347 33786 7359
rect 33699 7333 33786 7347
rect 27990 4485 28310 4525
rect 27990 4259 28023 4485
rect 28259 4259 28310 4485
rect 27990 4223 28310 4259
rect 20027 3416 20444 3462
rect 20027 3193 20069 3416
rect 20374 3193 20444 3416
rect 20027 3126 20444 3193
rect 18871 2703 19172 2897
rect 19390 2703 19621 2897
rect 18871 -4097 19621 2703
rect 18871 -4640 19016 -4097
rect 19333 -4640 19621 -4097
rect 18871 -7733 19621 -4640
rect 20070 -4934 20353 3126
rect 28027 1821 28261 4223
rect 32588 3464 33088 3505
rect 32588 3090 32613 3464
rect 33033 3090 33088 3464
rect 32588 3048 33088 3090
rect 33863 2387 34083 7820
rect 34140 7446 34252 7465
rect 34140 7338 34151 7446
rect 34237 7338 34252 7446
rect 34140 7321 34252 7338
rect 33863 2367 34082 2387
rect 33824 2330 34082 2367
rect 33824 2124 33880 2330
rect 34068 2124 34082 2330
rect 33824 2062 34082 2124
rect 28027 1665 28065 1821
rect 28228 1665 28261 1821
rect 28027 1626 28261 1665
rect 33883 1647 34022 1666
rect 33883 1541 33894 1647
rect 34008 1541 34022 1647
rect 33883 1531 34022 1541
rect 33883 -1051 34020 1531
rect 34149 -820 34229 7321
rect 34320 4580 34527 9810
rect 34703 7749 34882 7784
rect 34703 7639 34728 7749
rect 34864 7639 34882 7749
rect 34703 7594 34882 7639
rect 34289 4511 34610 4580
rect 34289 4239 34321 4511
rect 34580 4239 34610 4511
rect 34289 4173 34610 4239
rect 34704 3019 34846 7594
rect 34940 7167 35085 11930
rect 34933 7155 35087 7167
rect 34933 7068 34948 7155
rect 35070 7068 35087 7155
rect 34933 7058 35087 7068
rect 34940 5268 35085 7058
rect 34940 5158 34958 5268
rect 35071 5158 35085 5268
rect 34940 5150 35085 5158
rect 35201 6164 35346 11931
rect 35500 11929 35699 11961
rect 41644 11933 41698 12213
rect 42092 11933 42163 12213
rect 35540 8960 35681 11929
rect 41644 11850 42163 11933
rect 35500 8920 35710 8960
rect 35500 8790 35530 8920
rect 35670 8790 35710 8920
rect 35500 8760 35710 8790
rect 41030 8920 41190 8940
rect 41030 8790 41050 8920
rect 41170 8790 41190 8920
rect 41030 8770 41190 8790
rect 36673 8308 36811 8325
rect 36673 8211 36696 8308
rect 36795 8211 36811 8308
rect 36673 8187 36811 8211
rect 36723 7772 36810 8187
rect 36723 7756 36831 7772
rect 36723 7691 36743 7756
rect 36814 7691 36831 7756
rect 36723 7679 36831 7691
rect 36723 7676 36810 7679
rect 35201 6147 35347 6164
rect 35201 6036 35217 6147
rect 35329 6036 35347 6147
rect 35201 6019 35347 6036
rect 40463 6100 40523 6150
rect 41040 6130 41180 8770
rect 41040 6100 41610 6130
rect 34318 2877 34846 3019
rect 34108 -839 34251 -820
rect 34108 -969 34119 -839
rect 34237 -969 34251 -839
rect 34108 -982 34251 -969
rect 33879 -1061 34025 -1051
rect 33879 -1160 33893 -1061
rect 34011 -1160 34025 -1061
rect 33879 -1165 34025 -1160
rect 34318 -4895 34460 2877
rect 34551 2763 34680 2780
rect 34551 2622 34562 2763
rect 34665 2622 34680 2763
rect 34551 2601 34680 2622
rect 34558 1193 34663 2601
rect 34731 2455 34935 2492
rect 34731 2297 34759 2455
rect 34905 2297 34935 2455
rect 34731 2262 34935 2297
rect 34755 1225 34902 2262
rect 35201 2044 35346 6019
rect 40463 6000 41610 6100
rect 41040 5990 41610 6000
rect 38862 5623 39024 5630
rect 38862 5565 38878 5623
rect 39010 5565 39024 5623
rect 38862 5558 39024 5565
rect 39242 5623 39408 5635
rect 39242 5563 39259 5623
rect 39393 5563 39408 5623
rect 39242 5558 39408 5563
rect 37887 5487 38018 5511
rect 37887 5388 37904 5487
rect 37999 5388 38018 5487
rect 37887 5372 38018 5388
rect 37894 3471 38016 5372
rect 38610 5260 38740 5280
rect 38610 5170 38620 5260
rect 38730 5170 38740 5260
rect 38610 5150 38740 5170
rect 37815 3415 38032 3471
rect 37815 3247 37856 3415
rect 38001 3247 38032 3415
rect 37815 3171 38032 3247
rect 35185 2024 35372 2044
rect 35185 1899 35214 2024
rect 35346 1899 35372 2024
rect 35185 1872 35372 1899
rect 37477 2008 37606 2030
rect 37477 1902 37502 2008
rect 37585 1902 37606 2008
rect 37477 1881 37606 1902
rect 34550 1175 34672 1193
rect 34550 1088 34564 1175
rect 34662 1088 34672 1175
rect 34755 1162 35323 1225
rect 34550 1068 34672 1088
rect 36204 1139 36286 1146
rect 36204 1075 36211 1139
rect 36279 1075 36286 1139
rect 37512 1126 37575 1881
rect 38637 1170 38700 5150
rect 38870 1650 39020 5558
rect 38870 1560 38890 1650
rect 39000 1560 39020 1650
rect 39250 1660 39400 5558
rect 39707 5451 39887 5470
rect 39707 5348 39733 5451
rect 39863 5348 39887 5451
rect 39707 5309 39887 5348
rect 41140 5395 41368 5415
rect 39250 1590 39270 1660
rect 39390 1590 39400 1660
rect 39250 1580 39400 1590
rect 38870 1550 39020 1560
rect 39736 1185 39881 5309
rect 41140 5288 41168 5395
rect 41335 5288 41368 5395
rect 41140 5244 41368 5288
rect 40772 3478 40932 3492
rect 40772 3333 40784 3478
rect 40913 3333 40932 3478
rect 40772 3318 40932 3333
rect 40783 1850 40929 3318
rect 40758 1825 40961 1850
rect 40758 1710 40793 1825
rect 40930 1710 40961 1825
rect 40758 1684 40961 1710
rect 39734 1167 39882 1185
rect 36204 1066 36286 1075
rect 39734 1037 39754 1167
rect 39872 1037 39882 1167
rect 39734 1018 39882 1037
rect 39736 1016 39881 1018
rect 37238 272 37329 284
rect 40844 283 40979 302
rect 40844 277 40858 283
rect 37238 204 37249 272
rect 37317 204 37329 272
rect 37238 197 37329 204
rect 40843 200 40858 277
rect 40964 200 40979 283
rect 40843 182 40979 200
rect 35883 84 35985 94
rect 35883 7 35893 84
rect 35976 7 35985 84
rect 35883 -5 35985 7
rect 35889 -859 35982 -848
rect 35889 -938 35895 -859
rect 35978 -938 35982 -859
rect 35889 -949 35982 -938
rect 37013 -855 37113 -846
rect 37013 -933 37022 -855
rect 37101 -874 37113 -855
rect 37108 -927 37113 -874
rect 37101 -933 37113 -927
rect 37013 -940 37113 -933
rect 34767 -1892 34909 -1880
rect 34767 -2000 34780 -1892
rect 34897 -2000 34909 -1892
rect 34767 -2017 34909 -2000
rect 36196 -1924 36287 -1916
rect 36196 -1996 36205 -1924
rect 36279 -1996 36287 -1924
rect 36196 -2004 36287 -1996
rect 18871 -8031 19101 -7733
rect 19398 -8031 19621 -7733
rect 18871 -16979 19621 -8031
rect 19806 -5217 20353 -4934
rect 34226 -4954 34596 -4895
rect 34226 -5168 34281 -4954
rect 34547 -5168 34596 -4954
rect 19806 -10256 20089 -5217
rect 34226 -5220 34596 -5168
rect 34790 -5539 34904 -2017
rect 35155 -2569 35392 -2546
rect 40843 -2569 40971 182
rect 35155 -2707 35175 -2569
rect 35355 -2707 35392 -2569
rect 35155 -2732 35392 -2707
rect 40834 -2590 41014 -2569
rect 34768 -5560 34931 -5539
rect 34768 -5708 34788 -5560
rect 34910 -5708 34931 -5560
rect 34768 -5732 34931 -5708
rect 35189 -8000 35353 -2732
rect 40834 -2791 40849 -2590
rect 40987 -2791 41014 -2590
rect 40834 -2804 41014 -2791
rect 41169 -5943 41328 5244
rect 41470 2470 41610 5990
rect 41708 5519 42114 11850
rect 43491 8498 43585 8505
rect 43491 8407 43499 8498
rect 43577 8407 43585 8498
rect 43491 8394 43585 8407
rect 43136 8029 43257 8056
rect 43136 7945 43149 8029
rect 43238 7945 43257 8029
rect 43136 7932 43257 7945
rect 42436 7793 42610 7811
rect 42436 7690 42458 7793
rect 42589 7690 42610 7793
rect 42436 7676 42610 7690
rect 42204 7564 42373 7576
rect 42204 7438 42218 7564
rect 42355 7438 42373 7564
rect 42204 7419 42373 7438
rect 41704 5484 42114 5519
rect 41704 5338 41778 5484
rect 42037 5338 42114 5484
rect 41704 5307 42114 5338
rect 41708 5090 42114 5094
rect 41702 5053 42114 5090
rect 41702 4795 41757 5053
rect 42024 4795 42114 5053
rect 41702 4717 42114 4795
rect 41460 2450 41640 2470
rect 41460 2280 41480 2450
rect 41630 2280 41640 2450
rect 41460 2250 41640 2280
rect 41708 915 42114 4717
rect 42208 2793 42365 7419
rect 42201 2792 42374 2793
rect 42199 2782 42377 2792
rect 42199 2603 42213 2782
rect 42369 2603 42377 2782
rect 42199 2591 42377 2603
rect 41708 797 42116 915
rect 41708 480 41837 797
rect 42106 480 42116 797
rect 41708 317 42116 480
rect 41708 81 42118 317
rect 41708 -2854 42116 81
rect 41708 -2932 42316 -2854
rect 41701 -2990 42316 -2932
rect 41701 -3242 41771 -2990
rect 42236 -3242 42316 -2990
rect 41701 -3316 42316 -3242
rect 41708 -4991 42316 -3316
rect 42455 -4298 42603 7676
rect 42819 6613 42993 6614
rect 42818 6600 42993 6613
rect 42818 6474 42834 6600
rect 42970 6474 42993 6600
rect 42818 4516 42993 6474
rect 43151 6161 43255 7932
rect 43500 7836 43586 7846
rect 43500 7759 43510 7836
rect 43575 7759 43586 7836
rect 43500 7749 43586 7759
rect 43489 6590 43651 6606
rect 43489 6512 43530 6590
rect 43610 6512 43651 6590
rect 43489 6494 43651 6512
rect 43151 6057 43329 6161
rect 42708 4471 43121 4516
rect 42708 4310 42782 4471
rect 43061 4310 43121 4471
rect 42708 4265 43121 4310
rect 42890 -734 42947 4265
rect 43225 3483 43329 6057
rect 57001 5739 57751 8305
rect 57001 5320 57242 5739
rect 57547 5320 57751 5739
rect 43060 3379 43329 3483
rect 56354 3492 56692 3519
rect 43060 2187 43164 3379
rect 56354 3260 56384 3492
rect 56662 3260 56692 3492
rect 56354 3217 56692 3260
rect 43378 2187 43473 2203
rect 43060 2178 43473 2187
rect 43060 2098 43396 2178
rect 43457 2098 43473 2178
rect 43060 2083 43473 2098
rect 43378 2071 43473 2083
rect 43034 549 43146 560
rect 43034 473 43051 549
rect 43135 473 43146 549
rect 43366 547 43458 551
rect 43366 485 43376 547
rect 43448 485 43458 547
rect 43366 482 43458 485
rect 43034 458 43146 473
rect 43046 103 43140 458
rect 43040 87 43152 103
rect 43040 11 43056 87
rect 43140 11 43152 87
rect 43040 -1 43152 11
rect 42890 -791 43679 -734
rect 55980 -2585 56278 -2546
rect 55980 -2807 56003 -2585
rect 56241 -2807 56278 -2585
rect 55980 -2852 56278 -2807
rect 42454 -4352 42680 -4298
rect 42454 -4605 42485 -4352
rect 42645 -4605 42680 -4352
rect 42454 -4656 42680 -4605
rect 41169 -6102 41567 -5943
rect 35189 -8971 35271 -8000
rect 35189 -8972 35336 -8971
rect 19807 -12000 20087 -10256
rect 19804 -12058 20143 -12000
rect 19804 -12310 19869 -12058
rect 20071 -12310 20143 -12058
rect 19804 -12397 20143 -12310
rect 35186 -12834 35336 -8972
rect 38608 -10288 39073 -10254
rect 38608 -10438 38709 -10288
rect 38970 -10438 39073 -10288
rect 35138 -12875 35375 -12834
rect 35138 -13044 35169 -12875
rect 35348 -13044 35375 -12875
rect 35138 -13077 35375 -13044
rect 18871 -17246 19155 -16979
rect 19388 -17246 19621 -16979
rect 18871 -21147 19621 -17246
rect 38608 -14965 39073 -10438
rect 41408 -12161 41567 -6102
rect 41708 -9877 42116 -4991
rect 42328 -5549 42544 -5529
rect 56008 -5530 56265 -2852
rect 42328 -5722 42348 -5549
rect 42526 -5722 42544 -5549
rect 55770 -5666 56265 -5530
rect 42328 -5756 42544 -5722
rect 42350 -7540 42529 -5756
rect 42326 -7564 42560 -7540
rect 42326 -7728 42354 -7564
rect 42530 -7728 42560 -7564
rect 42326 -7750 42560 -7728
rect 55478 -8618 55756 -8589
rect 55478 -8866 55495 -8618
rect 55721 -8866 55756 -8618
rect 55478 -8880 55756 -8866
rect 41708 -10171 42316 -9877
rect 41708 -10421 41745 -10171
rect 42266 -10421 42316 -10171
rect 41708 -10469 42316 -10421
rect 41273 -12235 41674 -12161
rect 41273 -12413 41335 -12235
rect 41604 -12413 41674 -12235
rect 41273 -12454 41674 -12413
rect 38608 -15247 38672 -14965
rect 39016 -15247 39073 -14965
rect 35977 -18806 36310 -18773
rect 35977 -19007 36043 -18806
rect 36207 -19007 36310 -18806
rect 17794 -21374 18567 -21293
rect 17794 -21836 17929 -21374
rect 18465 -21836 18567 -21374
rect 35977 -21412 36310 -19007
rect 17794 -21924 18567 -21836
rect 35823 -21527 36450 -21412
rect 35823 -21809 35912 -21527
rect 36348 -21809 36450 -21527
rect 35823 -21873 36450 -21809
rect 17794 -21951 18560 -21924
rect 38608 -22941 39073 -15247
rect 41992 -16829 42276 -16807
rect 41992 -17003 42022 -16829
rect 42239 -17003 42276 -16829
rect 41992 -17041 42276 -17003
rect 42891 -16856 43179 -16830
rect 42891 -16990 42947 -16856
rect 43146 -16990 43179 -16856
rect 42891 -17026 43179 -16990
rect 42019 -21404 42241 -17041
rect 56404 -19713 56685 3217
rect 57001 -1680 57751 5320
rect 57001 -2071 57206 -1680
rect 57480 -2071 57751 -1680
rect 57001 -4082 57751 -2071
rect 57001 -4667 57286 -4082
rect 57576 -4667 57751 -4082
rect 57001 -9726 57751 -4667
rect 57001 -10051 57237 -9726
rect 57490 -10051 57751 -9726
rect 57001 -16141 57751 -10051
rect 57001 -16560 57269 -16141
rect 57584 -16560 57751 -16141
rect 56390 -19738 56703 -19713
rect 56390 -19908 56421 -19738
rect 56676 -19908 56703 -19738
rect 56390 -19946 56703 -19908
rect 57001 -21282 57751 -16560
rect 58223 4673 58973 8277
rect 58223 4114 58446 4673
rect 58860 4114 58973 4673
rect 58223 -8539 58973 4114
rect 58223 -8967 58398 -8539
rect 58813 -8967 58973 -8539
rect 58223 -21286 58973 -8967
rect 58202 -21340 58979 -21286
rect 41930 -21483 42382 -21404
rect 41930 -21764 41995 -21483
rect 42303 -21764 42382 -21483
rect 41930 -21823 42382 -21764
rect 58202 -21871 58283 -21340
rect 58922 -21871 58979 -21340
rect 58202 -21942 58979 -21871
rect 38465 -23059 39241 -22941
rect 38465 -23526 38572 -23059
rect 39145 -23526 39241 -23059
rect 38465 -23610 39241 -23526
<< via2 >>
rect 19179 10964 19388 11180
rect 18015 4174 18361 4646
rect 18068 -6036 18326 -5667
rect 33865 8358 34022 8387
rect 33865 8183 33891 8358
rect 33891 8183 34002 8358
rect 34002 8183 34022 8358
rect 33865 8160 34022 8183
rect 33877 7836 34060 7980
rect 33707 7419 33778 7436
rect 33707 7359 33778 7419
rect 33707 7347 33778 7359
rect 28023 4259 28259 4485
rect 20069 3193 20374 3416
rect 19172 2873 19390 2897
rect 19172 2716 19196 2873
rect 19196 2716 19360 2873
rect 19360 2716 19390 2873
rect 19172 2703 19390 2716
rect 19016 -4176 19333 -4097
rect 19016 -4572 19061 -4176
rect 19061 -4572 19310 -4176
rect 19310 -4572 19333 -4176
rect 19016 -4640 19333 -4572
rect 32613 3397 33033 3464
rect 32613 3159 32655 3397
rect 32655 3159 32948 3397
rect 32948 3159 33033 3397
rect 32613 3090 33033 3159
rect 34151 7338 34237 7446
rect 34728 7639 34864 7749
rect 34321 4239 34580 4511
rect 35530 8790 35670 8920
rect 41050 8790 41170 8920
rect 36696 8211 36795 8308
rect 36743 7691 36814 7756
rect 34119 -969 34237 -839
rect 33893 -1160 34011 -1061
rect 37904 5388 37999 5487
rect 36211 1134 36279 1139
rect 36211 1075 36213 1134
rect 36213 1075 36273 1134
rect 36273 1075 36279 1134
rect 41168 5288 41335 5395
rect 40784 3333 40913 3478
rect 40793 1710 40930 1825
rect 37249 271 37317 272
rect 37249 213 37251 271
rect 37251 213 37308 271
rect 37308 213 37317 271
rect 37249 204 37317 213
rect 40858 200 40964 283
rect 35893 73 35976 84
rect 35893 19 35903 73
rect 35903 19 35972 73
rect 35972 19 35976 73
rect 35893 7 35976 19
rect 35895 -873 35978 -859
rect 35895 -926 35902 -873
rect 35902 -926 35975 -873
rect 35975 -926 35978 -873
rect 35895 -938 35978 -926
rect 37022 -874 37101 -855
rect 37022 -927 37032 -874
rect 37032 -927 37101 -874
rect 37022 -933 37101 -927
rect 36205 -1929 36279 -1924
rect 36205 -1992 36210 -1929
rect 36210 -1992 36276 -1929
rect 36276 -1992 36279 -1929
rect 36205 -1996 36279 -1992
rect 19101 -7739 19398 -7733
rect 19101 -8019 19119 -7739
rect 19119 -8019 19368 -7739
rect 19368 -8019 19398 -7739
rect 19101 -8031 19398 -8019
rect 35175 -2707 35355 -2569
rect 40849 -2791 40987 -2590
rect 43499 8494 43577 8498
rect 43499 8412 43502 8494
rect 43502 8412 43573 8494
rect 43573 8412 43577 8494
rect 43499 8407 43577 8412
rect 43149 7945 43238 8029
rect 42458 7690 42589 7793
rect 42218 7438 42355 7564
rect 42834 6474 42970 6600
rect 43510 7831 43575 7836
rect 43510 7768 43521 7831
rect 43521 7768 43575 7831
rect 43510 7759 43575 7768
rect 43530 6512 43610 6590
rect 42782 4310 43061 4471
rect 57242 5698 57547 5739
rect 57242 5367 57270 5698
rect 57270 5367 57533 5698
rect 57533 5367 57547 5698
rect 57242 5320 57547 5367
rect 56384 3260 56662 3492
rect 43051 473 43135 549
rect 43376 544 43448 547
rect 43376 488 43380 544
rect 43380 488 43440 544
rect 43440 488 43448 544
rect 43376 485 43448 488
rect 43056 11 43140 87
rect 56003 -2807 56241 -2585
rect 19155 -17013 19388 -16979
rect 19155 -17206 19180 -17013
rect 19180 -17206 19363 -17013
rect 19363 -17206 19388 -17013
rect 19155 -17246 19388 -17206
rect 55495 -8641 55721 -8618
rect 55495 -8825 55513 -8641
rect 55513 -8825 55696 -8641
rect 55696 -8825 55721 -8641
rect 55495 -8866 55721 -8825
rect 17929 -21836 18465 -21374
rect 35912 -21809 36348 -21527
rect 42022 -17003 42239 -16829
rect 42947 -16990 43146 -16856
rect 57206 -2071 57480 -1680
rect 57286 -4138 57576 -4082
rect 57286 -4593 57314 -4138
rect 57314 -4593 57541 -4138
rect 57541 -4593 57576 -4138
rect 57286 -4667 57576 -4593
rect 57237 -9746 57490 -9726
rect 57237 -10038 57251 -9746
rect 57251 -10038 57457 -9746
rect 57457 -10038 57490 -9746
rect 57237 -10051 57490 -10038
rect 57269 -16173 57584 -16141
rect 57269 -16547 57289 -16173
rect 57289 -16547 57564 -16173
rect 57564 -16547 57584 -16173
rect 57269 -16560 57584 -16547
rect 58446 4114 58860 4673
rect 58398 -8967 58813 -8539
rect 41995 -21764 42303 -21483
rect 58283 -21871 58922 -21340
<< metal3 >>
rect 19158 11180 19415 11195
rect 19158 10964 19179 11180
rect 19388 11103 19415 11180
rect 19388 11026 21798 11103
rect 19388 10964 19415 11026
rect 19158 10929 19415 10964
rect 35500 8930 35710 8960
rect 41030 8930 41190 8940
rect 35500 8920 41190 8930
rect 35500 8790 35530 8920
rect 35670 8790 41050 8920
rect 41170 8790 41190 8920
rect 35500 8760 35710 8790
rect 41030 8770 41190 8790
rect 43491 8498 43585 8505
rect 43491 8493 43499 8498
rect 33844 8387 34045 8418
rect 33844 8160 33865 8387
rect 34022 8322 34045 8387
rect 38828 8407 43499 8493
rect 43577 8407 43585 8498
rect 36673 8322 36811 8325
rect 34022 8308 36811 8322
rect 34022 8211 36696 8308
rect 36795 8211 36811 8308
rect 34022 8187 36811 8211
rect 34022 8184 36808 8187
rect 34022 8160 34045 8184
rect 33844 8137 34045 8160
rect 33855 7998 34077 8002
rect 33855 7980 38123 7998
rect 33855 7836 33877 7980
rect 34060 7911 38123 7980
rect 34060 7910 37811 7911
rect 34060 7836 34077 7910
rect 33855 7820 34077 7836
rect 34703 7766 34882 7784
rect 34703 7749 36674 7766
rect 34703 7639 34728 7749
rect 34864 7700 36674 7749
rect 34864 7639 34882 7700
rect 34703 7594 34882 7639
rect 33699 7446 33786 7447
rect 34140 7446 34252 7465
rect 33699 7436 34151 7446
rect 33699 7347 33707 7436
rect 33778 7347 34151 7436
rect 33699 7338 34151 7347
rect 34237 7338 34253 7446
rect 36608 7427 36674 7700
rect 36731 7756 36831 7772
rect 36731 7691 36743 7756
rect 36814 7691 36831 7756
rect 36731 7679 36831 7691
rect 36731 7460 36802 7679
rect 38036 7440 38123 7911
rect 38828 7424 38914 8407
rect 43491 8394 43585 8407
rect 43136 8029 43257 8056
rect 43136 8016 43149 8029
rect 39048 7958 43149 8016
rect 39048 7441 39106 7958
rect 43136 7945 43149 7958
rect 43238 7945 43257 8029
rect 43136 7932 43257 7945
rect 43500 7839 43586 7846
rect 42859 7836 43586 7839
rect 42436 7793 42610 7811
rect 42436 7761 42458 7793
rect 39886 7409 39972 7759
rect 40148 7701 42458 7761
rect 40148 7444 40208 7701
rect 42436 7690 42458 7701
rect 42589 7690 42610 7793
rect 42436 7676 42610 7690
rect 42859 7759 43510 7836
rect 43575 7759 43586 7836
rect 42859 7758 43586 7759
rect 42204 7564 42373 7576
rect 42859 7564 42957 7758
rect 43500 7749 43586 7758
rect 42204 7438 42218 7564
rect 42355 7438 42957 7564
rect 42204 7423 42957 7438
rect 42204 7419 42373 7423
rect 33699 7333 34253 7338
rect 34140 7321 34252 7333
rect 42819 6607 42993 6614
rect 42819 6606 43602 6607
rect 42819 6600 43651 6606
rect 37916 5511 38002 6591
rect 42819 6474 42834 6600
rect 42970 6590 43651 6600
rect 42970 6512 43530 6590
rect 43610 6512 43651 6590
rect 42970 6494 43651 6512
rect 42970 6474 42993 6494
rect 42819 6454 42993 6474
rect 37887 5487 38018 5511
rect 37887 5388 37904 5487
rect 37999 5388 38018 5487
rect 37887 5372 38018 5388
rect 39886 5359 39972 6312
rect 57209 5739 57574 5773
rect 57209 5557 57242 5739
rect 53733 5480 57242 5557
rect 41140 5395 41368 5415
rect 41140 5359 41168 5395
rect 39886 5288 41168 5359
rect 41335 5288 41368 5395
rect 39886 5273 41368 5288
rect 57209 5320 57242 5480
rect 57547 5320 57574 5739
rect 57209 5279 57574 5320
rect 41140 5244 41368 5273
rect 17918 4646 18476 4749
rect 17918 4174 18015 4646
rect 18361 4578 18476 4646
rect 58325 4673 58921 4807
rect 34257 4578 34638 4580
rect 58325 4578 58446 4673
rect 18361 4511 58446 4578
rect 18361 4485 34321 4511
rect 18361 4259 28023 4485
rect 28259 4259 34321 4485
rect 18361 4239 34321 4259
rect 34580 4471 58446 4511
rect 34580 4310 42782 4471
rect 43061 4310 58446 4471
rect 34580 4239 58446 4310
rect 18361 4174 58446 4239
rect 17918 4083 18476 4174
rect 34257 4173 34638 4174
rect 58325 4114 58446 4174
rect 58860 4114 58921 4673
rect 58325 4004 58921 4114
rect 32588 3464 33088 3505
rect 56354 3492 56692 3519
rect 20027 3416 20444 3462
rect 20027 3193 20069 3416
rect 20374 3413 20444 3416
rect 32588 3413 32613 3464
rect 20374 3193 32613 3413
rect 20027 3176 32613 3193
rect 20027 3126 20444 3176
rect 32588 3090 32613 3176
rect 33033 3090 33088 3464
rect 40772 3478 56384 3492
rect 40772 3333 40784 3478
rect 40913 3333 56384 3478
rect 40772 3318 56384 3333
rect 56354 3260 56384 3318
rect 56662 3260 56692 3492
rect 56354 3217 56692 3260
rect 32588 3048 33088 3090
rect 19154 2897 19426 2933
rect 19154 2703 19172 2897
rect 19390 2848 19426 2897
rect 19390 2752 24487 2848
rect 19390 2703 19426 2752
rect 19154 2679 19426 2703
rect 40758 1825 40961 1850
rect 40758 1786 40793 1825
rect 36204 1710 40793 1786
rect 40930 1710 40961 1825
rect 36204 1704 40961 1710
rect 36204 1139 36286 1704
rect 40758 1684 40961 1704
rect 36204 1075 36211 1139
rect 36279 1075 36286 1139
rect 36204 1066 36286 1075
rect 43034 551 43146 560
rect 43034 549 43458 551
rect 43034 473 43051 549
rect 43135 547 43458 549
rect 43135 485 43376 547
rect 43448 485 43458 547
rect 43135 481 43458 485
rect 43135 473 43146 481
rect 43034 458 43146 473
rect 37238 278 37329 284
rect 40844 283 40979 302
rect 40844 278 40858 283
rect 37238 272 40858 278
rect 37238 204 37249 272
rect 37317 204 40858 272
rect 37238 200 40858 204
rect 40964 200 40979 283
rect 37238 199 40979 200
rect 37238 197 37329 199
rect 40844 182 40979 199
rect 35883 89 35985 94
rect 43040 89 43152 103
rect 35883 87 43152 89
rect 35883 84 43056 87
rect 35883 7 35893 84
rect 35976 11 43056 84
rect 43140 11 43152 87
rect 35976 7 43152 11
rect 35883 2 43152 7
rect 35883 -5 35985 2
rect 43040 -1 43152 2
rect 34108 -839 34251 -820
rect 34108 -969 34119 -839
rect 34237 -850 34251 -839
rect 35889 -850 35982 -848
rect 34237 -859 35982 -850
rect 34237 -938 35895 -859
rect 35978 -938 35982 -859
rect 34237 -946 35982 -938
rect 34237 -969 34251 -946
rect 35889 -949 35982 -946
rect 37013 -855 37113 -846
rect 37013 -933 37022 -855
rect 37101 -933 37113 -855
rect 34108 -982 34251 -969
rect 33879 -1059 34025 -1051
rect 37013 -1059 37113 -933
rect 33879 -1061 37113 -1059
rect 33879 -1160 33893 -1061
rect 34011 -1159 37113 -1061
rect 34011 -1160 34025 -1159
rect 33879 -1165 34025 -1160
rect 57144 -1680 57542 -1584
rect 57144 -1829 57206 -1680
rect 52444 -1906 57206 -1829
rect 36196 -1924 36287 -1916
rect 36196 -1996 36205 -1924
rect 36279 -1996 36287 -1924
rect 36196 -2004 36287 -1996
rect 35155 -2569 35392 -2546
rect 35155 -2707 35175 -2569
rect 35355 -2586 35392 -2569
rect 36196 -2586 36284 -2004
rect 57144 -2071 57206 -1906
rect 57480 -2071 57542 -1680
rect 57144 -2201 57542 -2071
rect 35355 -2674 36284 -2586
rect 40834 -2571 41014 -2569
rect 55980 -2571 56278 -2546
rect 40834 -2585 56278 -2571
rect 40834 -2590 56003 -2585
rect 35355 -2707 35392 -2674
rect 35155 -2732 35392 -2707
rect 40834 -2791 40849 -2590
rect 40987 -2791 56003 -2590
rect 40834 -2804 56003 -2791
rect 55980 -2807 56003 -2804
rect 56241 -2807 56278 -2585
rect 55980 -2852 56278 -2807
rect 18971 -4097 19435 -3950
rect 18971 -4640 19016 -4097
rect 19333 -4165 19435 -4097
rect 57240 -4082 57627 -3991
rect 57240 -4165 57286 -4082
rect 19333 -4569 57286 -4165
rect 19333 -4640 19435 -4569
rect 18971 -4719 19435 -4640
rect 57240 -4667 57286 -4569
rect 57576 -4667 57627 -4082
rect 57240 -4718 57627 -4667
rect 18018 -5667 18388 -5581
rect 18018 -6036 18068 -5667
rect 18326 -5855 18388 -5667
rect 18326 -5944 20728 -5855
rect 18326 -6036 18388 -5944
rect 18018 -6110 18388 -6036
rect 19088 -7733 19417 -7703
rect 19088 -8031 19101 -7733
rect 19398 -7844 19417 -7733
rect 19398 -7961 21052 -7844
rect 19398 -8031 19417 -7961
rect 19088 -8079 19417 -8031
rect 58352 -8539 58873 -8459
rect 58352 -8586 58398 -8539
rect 55478 -8618 58398 -8586
rect 55478 -8866 55495 -8618
rect 55721 -8866 58398 -8618
rect 55478 -8880 58398 -8866
rect 58352 -8967 58398 -8880
rect 58813 -8967 58873 -8539
rect 58352 -9020 58873 -8967
rect 57244 -9679 57490 -9673
rect 57211 -9726 57563 -9679
rect 57211 -9879 57237 -9726
rect 52242 -9936 57237 -9879
rect 57211 -10051 57237 -9936
rect 57490 -10051 57563 -9726
rect 57211 -10104 57563 -10051
rect 20882 -11188 55877 -10784
rect 57220 -16141 57646 -16072
rect 57220 -16311 57269 -16141
rect 53784 -16459 57269 -16311
rect 57220 -16560 57269 -16459
rect 57584 -16560 57646 -16141
rect 57220 -16623 57646 -16560
rect 41992 -16829 42276 -16807
rect 19108 -16979 19454 -16917
rect 19108 -17246 19155 -16979
rect 19388 -17066 19454 -16979
rect 41992 -17003 42022 -16829
rect 42239 -16856 43193 -16829
rect 42239 -16990 42947 -16856
rect 43146 -16990 43193 -16856
rect 42239 -17003 43193 -16990
rect 41992 -17032 43193 -17003
rect 41992 -17041 42276 -17032
rect 19388 -17147 23318 -17066
rect 19388 -17246 19454 -17147
rect 19108 -17290 19454 -17246
rect 58202 -21289 58979 -21286
rect 17773 -21340 58979 -21289
rect 17773 -21374 58283 -21340
rect 17773 -21836 17929 -21374
rect 18465 -21483 58283 -21374
rect 18465 -21527 41995 -21483
rect 18465 -21809 35912 -21527
rect 36348 -21764 41995 -21527
rect 42303 -21764 58283 -21483
rect 36348 -21809 58283 -21764
rect 18465 -21836 58283 -21809
rect 17773 -21871 58283 -21836
rect 58922 -21871 58979 -21340
rect 17773 -21942 58979 -21871
rect 17773 -21947 58961 -21942
rect 17794 -21951 18560 -21947
use CLK_div_90_mag  CLK_div_90_mag_0
timestamp 1695206022
transform 1 0 18281 0 1 301
box 3140 4330 16201 11389
use CLK_div_93_mag  CLK_div_93_mag_0
timestamp 1695206022
transform 1 0 20761 0 1 -10236
box -502 -242 21015 5340
use CLK_div_96_mag  CLK_div_96_mag_0
timestamp 1695206022
transform 1 0 21556 0 1 -3347
box 40 105 9646 6783
use CLK_div_99_mag  CLK_div_99_mag_0
timestamp 1695206022
transform 1 0 19954 0 1 -28521
box 1317 7658 17710 16746
use CLK_div_100_mag  CLK_div_100_mag_0
timestamp 1695206022
transform 1 0 43329 0 1 -2455
box -125 0 12197 5567
use CLK_div_105_mag  CLK_div_105_mag_0
timestamp 1695206022
transform 1 0 43441 0 1 4931
box -125 0 12197 5567
use CLK_div_108_new_mag  CLK_div_108_new_mag_0
timestamp 1695206022
transform 1 0 36094 0 1 -10375
box 6435 -290 19896 6076
use CLK_div_110_mag  CLK_div_110_mag_0
timestamp 1695206022
transform 1 0 42879 0 1 -18358
box -2562 -2430 13288 6270
use dec3x8_ibr_mag  dec3x8_ibr_mag_0
timestamp 1695127730
transform 1 0 35812 0 1 6609
box -402 -1051 5095 1052
use mux_8x1_ibr  mux_8x1_ibr_0
timestamp 1695306401
transform 1 0 34946 0 1 -427
box 0 -2102 4512 2102
<< labels >>
flabel via1 18060 10950 18060 10950 0 FreeSans 1600 0 0 0 CLK
port 0 nsew
flabel via1 19040 11030 19040 11030 0 FreeSans 1600 0 0 0 RST
port 1 nsew
flabel via1 35010 12010 35010 12010 0 FreeSans 1600 0 0 0 F2
port 2 nsew
flabel via1 35260 12020 35260 12020 0 FreeSans 1600 0 0 0 F1
port 3 nsew
flabel via1 35580 12020 35580 12020 0 FreeSans 1600 0 0 0 F0
port 4 nsew
flabel via1 41850 12020 41850 12020 0 FreeSans 1600 0 0 0 Vdiv
port 5 nsew
flabel metal1 37780 11070 37780 11070 0 FreeSans 1600 0 0 0 VDD
port 6 nsew
flabel metal1 39430 -23230 39430 -23230 0 FreeSans 1600 0 0 0 VSS
port 7 nsew
flabel metal2 34180 -70 34180 -70 0 FreeSans 1600 0 0 0 Vdiv90
port 8 nsew
flabel metal1 31410 1580 31410 1580 0 FreeSans 1600 0 0 0 Vdiv96
port 9 nsew
flabel metal1 35060 -5630 35060 -5630 0 FreeSans 1600 0 0 0 Vdiv93
port 10 nsew
flabel metal1 35090 -12990 35090 -12990 0 FreeSans 1600 0 0 0 Vdiv99
port 11 nsew
flabel metal1 56060 -19860 56060 -19860 0 FreeSans 1600 0 0 0 Vdiv110
port 12 nsew
flabel metal2 40890 -1630 40890 -1630 0 FreeSans 1600 0 0 0 Vdiv108
port 13 nsew
flabel metal2 43100 230 43100 230 0 FreeSans 1600 0 0 0 Vdiv100
port 14 nsew
flabel metal2 42270 6740 42270 6740 0 FreeSans 1600 0 0 0 Vdiv105
port 15 nsew
flabel metal2 36760 8080 36760 8080 0 FreeSans 1600 0 0 0 VDD90
port 16 nsew
flabel metal1 32080 2230 32080 2230 0 FreeSans 1600 0 0 0 VDD96
port 17 nsew
flabel metal2 34360 -3880 34360 -3880 0 FreeSans 1600 0 0 0 VDD93
port 18 nsew
flabel metal1 20460 -12270 20460 -12270 0 FreeSans 1600 0 0 0 VDD99
port 19 nsew
flabel metal2 41480 -11920 41480 -11920 0 FreeSans 1600 0 0 0 VDD110
port 20 nsew
flabel metal2 42500 -1740 42500 -1740 0 FreeSans 1600 0 0 0 VDD108
port 21 nsew
flabel metal2 43270 3890 43270 3890 0 FreeSans 1600 0 0 0 VDD100
port 22 nsew
flabel metal3 41370 8440 41370 8440 0 FreeSans 1600 0 0 0 VDD105
port 23 nsew
<< end >>
