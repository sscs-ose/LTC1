magic
tech gf180mcuD
magscale 1 10
timestamp 1713866589
<< metal1 >>
rect -50 14000 50 14063
rect -50 -14063 50 -14000
<< rmetal1 >>
rect -50 -14000 50 14000
<< properties >>
string gencell rm1
string library gf180mcu
string parameters w 0.5 l 140 m 1 nx 1 wmin 0.16 lmin 0.16 rho 0.076 val 21.28 dummy 0 dw 0.0 term 0.0 roverlap 0 full_metal {}
<< end >>
