magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1715 -1319 1715 1319
<< metal4 >>
rect -712 311 712 316
rect -712 283 -707 311
rect -679 283 -641 311
rect -613 283 -575 311
rect -547 283 -509 311
rect -481 283 -443 311
rect -415 283 -377 311
rect -349 283 -311 311
rect -283 283 -245 311
rect -217 283 -179 311
rect -151 283 -113 311
rect -85 283 -47 311
rect -19 283 19 311
rect 47 283 85 311
rect 113 283 151 311
rect 179 283 217 311
rect 245 283 283 311
rect 311 283 349 311
rect 377 283 415 311
rect 443 283 481 311
rect 509 283 547 311
rect 575 283 613 311
rect 641 283 679 311
rect 707 283 712 311
rect -712 245 712 283
rect -712 217 -707 245
rect -679 217 -641 245
rect -613 217 -575 245
rect -547 217 -509 245
rect -481 217 -443 245
rect -415 217 -377 245
rect -349 217 -311 245
rect -283 217 -245 245
rect -217 217 -179 245
rect -151 217 -113 245
rect -85 217 -47 245
rect -19 217 19 245
rect 47 217 85 245
rect 113 217 151 245
rect 179 217 217 245
rect 245 217 283 245
rect 311 217 349 245
rect 377 217 415 245
rect 443 217 481 245
rect 509 217 547 245
rect 575 217 613 245
rect 641 217 679 245
rect 707 217 712 245
rect -712 179 712 217
rect -712 151 -707 179
rect -679 151 -641 179
rect -613 151 -575 179
rect -547 151 -509 179
rect -481 151 -443 179
rect -415 151 -377 179
rect -349 151 -311 179
rect -283 151 -245 179
rect -217 151 -179 179
rect -151 151 -113 179
rect -85 151 -47 179
rect -19 151 19 179
rect 47 151 85 179
rect 113 151 151 179
rect 179 151 217 179
rect 245 151 283 179
rect 311 151 349 179
rect 377 151 415 179
rect 443 151 481 179
rect 509 151 547 179
rect 575 151 613 179
rect 641 151 679 179
rect 707 151 712 179
rect -712 113 712 151
rect -712 85 -707 113
rect -679 85 -641 113
rect -613 85 -575 113
rect -547 85 -509 113
rect -481 85 -443 113
rect -415 85 -377 113
rect -349 85 -311 113
rect -283 85 -245 113
rect -217 85 -179 113
rect -151 85 -113 113
rect -85 85 -47 113
rect -19 85 19 113
rect 47 85 85 113
rect 113 85 151 113
rect 179 85 217 113
rect 245 85 283 113
rect 311 85 349 113
rect 377 85 415 113
rect 443 85 481 113
rect 509 85 547 113
rect 575 85 613 113
rect 641 85 679 113
rect 707 85 712 113
rect -712 47 712 85
rect -712 19 -707 47
rect -679 19 -641 47
rect -613 19 -575 47
rect -547 19 -509 47
rect -481 19 -443 47
rect -415 19 -377 47
rect -349 19 -311 47
rect -283 19 -245 47
rect -217 19 -179 47
rect -151 19 -113 47
rect -85 19 -47 47
rect -19 19 19 47
rect 47 19 85 47
rect 113 19 151 47
rect 179 19 217 47
rect 245 19 283 47
rect 311 19 349 47
rect 377 19 415 47
rect 443 19 481 47
rect 509 19 547 47
rect 575 19 613 47
rect 641 19 679 47
rect 707 19 712 47
rect -712 -19 712 19
rect -712 -47 -707 -19
rect -679 -47 -641 -19
rect -613 -47 -575 -19
rect -547 -47 -509 -19
rect -481 -47 -443 -19
rect -415 -47 -377 -19
rect -349 -47 -311 -19
rect -283 -47 -245 -19
rect -217 -47 -179 -19
rect -151 -47 -113 -19
rect -85 -47 -47 -19
rect -19 -47 19 -19
rect 47 -47 85 -19
rect 113 -47 151 -19
rect 179 -47 217 -19
rect 245 -47 283 -19
rect 311 -47 349 -19
rect 377 -47 415 -19
rect 443 -47 481 -19
rect 509 -47 547 -19
rect 575 -47 613 -19
rect 641 -47 679 -19
rect 707 -47 712 -19
rect -712 -85 712 -47
rect -712 -113 -707 -85
rect -679 -113 -641 -85
rect -613 -113 -575 -85
rect -547 -113 -509 -85
rect -481 -113 -443 -85
rect -415 -113 -377 -85
rect -349 -113 -311 -85
rect -283 -113 -245 -85
rect -217 -113 -179 -85
rect -151 -113 -113 -85
rect -85 -113 -47 -85
rect -19 -113 19 -85
rect 47 -113 85 -85
rect 113 -113 151 -85
rect 179 -113 217 -85
rect 245 -113 283 -85
rect 311 -113 349 -85
rect 377 -113 415 -85
rect 443 -113 481 -85
rect 509 -113 547 -85
rect 575 -113 613 -85
rect 641 -113 679 -85
rect 707 -113 712 -85
rect -712 -151 712 -113
rect -712 -179 -707 -151
rect -679 -179 -641 -151
rect -613 -179 -575 -151
rect -547 -179 -509 -151
rect -481 -179 -443 -151
rect -415 -179 -377 -151
rect -349 -179 -311 -151
rect -283 -179 -245 -151
rect -217 -179 -179 -151
rect -151 -179 -113 -151
rect -85 -179 -47 -151
rect -19 -179 19 -151
rect 47 -179 85 -151
rect 113 -179 151 -151
rect 179 -179 217 -151
rect 245 -179 283 -151
rect 311 -179 349 -151
rect 377 -179 415 -151
rect 443 -179 481 -151
rect 509 -179 547 -151
rect 575 -179 613 -151
rect 641 -179 679 -151
rect 707 -179 712 -151
rect -712 -217 712 -179
rect -712 -245 -707 -217
rect -679 -245 -641 -217
rect -613 -245 -575 -217
rect -547 -245 -509 -217
rect -481 -245 -443 -217
rect -415 -245 -377 -217
rect -349 -245 -311 -217
rect -283 -245 -245 -217
rect -217 -245 -179 -217
rect -151 -245 -113 -217
rect -85 -245 -47 -217
rect -19 -245 19 -217
rect 47 -245 85 -217
rect 113 -245 151 -217
rect 179 -245 217 -217
rect 245 -245 283 -217
rect 311 -245 349 -217
rect 377 -245 415 -217
rect 443 -245 481 -217
rect 509 -245 547 -217
rect 575 -245 613 -217
rect 641 -245 679 -217
rect 707 -245 712 -217
rect -712 -283 712 -245
rect -712 -311 -707 -283
rect -679 -311 -641 -283
rect -613 -311 -575 -283
rect -547 -311 -509 -283
rect -481 -311 -443 -283
rect -415 -311 -377 -283
rect -349 -311 -311 -283
rect -283 -311 -245 -283
rect -217 -311 -179 -283
rect -151 -311 -113 -283
rect -85 -311 -47 -283
rect -19 -311 19 -283
rect 47 -311 85 -283
rect 113 -311 151 -283
rect 179 -311 217 -283
rect 245 -311 283 -283
rect 311 -311 349 -283
rect 377 -311 415 -283
rect 443 -311 481 -283
rect 509 -311 547 -283
rect 575 -311 613 -283
rect 641 -311 679 -283
rect 707 -311 712 -283
rect -712 -316 712 -311
<< via4 >>
rect -707 283 -679 311
rect -641 283 -613 311
rect -575 283 -547 311
rect -509 283 -481 311
rect -443 283 -415 311
rect -377 283 -349 311
rect -311 283 -283 311
rect -245 283 -217 311
rect -179 283 -151 311
rect -113 283 -85 311
rect -47 283 -19 311
rect 19 283 47 311
rect 85 283 113 311
rect 151 283 179 311
rect 217 283 245 311
rect 283 283 311 311
rect 349 283 377 311
rect 415 283 443 311
rect 481 283 509 311
rect 547 283 575 311
rect 613 283 641 311
rect 679 283 707 311
rect -707 217 -679 245
rect -641 217 -613 245
rect -575 217 -547 245
rect -509 217 -481 245
rect -443 217 -415 245
rect -377 217 -349 245
rect -311 217 -283 245
rect -245 217 -217 245
rect -179 217 -151 245
rect -113 217 -85 245
rect -47 217 -19 245
rect 19 217 47 245
rect 85 217 113 245
rect 151 217 179 245
rect 217 217 245 245
rect 283 217 311 245
rect 349 217 377 245
rect 415 217 443 245
rect 481 217 509 245
rect 547 217 575 245
rect 613 217 641 245
rect 679 217 707 245
rect -707 151 -679 179
rect -641 151 -613 179
rect -575 151 -547 179
rect -509 151 -481 179
rect -443 151 -415 179
rect -377 151 -349 179
rect -311 151 -283 179
rect -245 151 -217 179
rect -179 151 -151 179
rect -113 151 -85 179
rect -47 151 -19 179
rect 19 151 47 179
rect 85 151 113 179
rect 151 151 179 179
rect 217 151 245 179
rect 283 151 311 179
rect 349 151 377 179
rect 415 151 443 179
rect 481 151 509 179
rect 547 151 575 179
rect 613 151 641 179
rect 679 151 707 179
rect -707 85 -679 113
rect -641 85 -613 113
rect -575 85 -547 113
rect -509 85 -481 113
rect -443 85 -415 113
rect -377 85 -349 113
rect -311 85 -283 113
rect -245 85 -217 113
rect -179 85 -151 113
rect -113 85 -85 113
rect -47 85 -19 113
rect 19 85 47 113
rect 85 85 113 113
rect 151 85 179 113
rect 217 85 245 113
rect 283 85 311 113
rect 349 85 377 113
rect 415 85 443 113
rect 481 85 509 113
rect 547 85 575 113
rect 613 85 641 113
rect 679 85 707 113
rect -707 19 -679 47
rect -641 19 -613 47
rect -575 19 -547 47
rect -509 19 -481 47
rect -443 19 -415 47
rect -377 19 -349 47
rect -311 19 -283 47
rect -245 19 -217 47
rect -179 19 -151 47
rect -113 19 -85 47
rect -47 19 -19 47
rect 19 19 47 47
rect 85 19 113 47
rect 151 19 179 47
rect 217 19 245 47
rect 283 19 311 47
rect 349 19 377 47
rect 415 19 443 47
rect 481 19 509 47
rect 547 19 575 47
rect 613 19 641 47
rect 679 19 707 47
rect -707 -47 -679 -19
rect -641 -47 -613 -19
rect -575 -47 -547 -19
rect -509 -47 -481 -19
rect -443 -47 -415 -19
rect -377 -47 -349 -19
rect -311 -47 -283 -19
rect -245 -47 -217 -19
rect -179 -47 -151 -19
rect -113 -47 -85 -19
rect -47 -47 -19 -19
rect 19 -47 47 -19
rect 85 -47 113 -19
rect 151 -47 179 -19
rect 217 -47 245 -19
rect 283 -47 311 -19
rect 349 -47 377 -19
rect 415 -47 443 -19
rect 481 -47 509 -19
rect 547 -47 575 -19
rect 613 -47 641 -19
rect 679 -47 707 -19
rect -707 -113 -679 -85
rect -641 -113 -613 -85
rect -575 -113 -547 -85
rect -509 -113 -481 -85
rect -443 -113 -415 -85
rect -377 -113 -349 -85
rect -311 -113 -283 -85
rect -245 -113 -217 -85
rect -179 -113 -151 -85
rect -113 -113 -85 -85
rect -47 -113 -19 -85
rect 19 -113 47 -85
rect 85 -113 113 -85
rect 151 -113 179 -85
rect 217 -113 245 -85
rect 283 -113 311 -85
rect 349 -113 377 -85
rect 415 -113 443 -85
rect 481 -113 509 -85
rect 547 -113 575 -85
rect 613 -113 641 -85
rect 679 -113 707 -85
rect -707 -179 -679 -151
rect -641 -179 -613 -151
rect -575 -179 -547 -151
rect -509 -179 -481 -151
rect -443 -179 -415 -151
rect -377 -179 -349 -151
rect -311 -179 -283 -151
rect -245 -179 -217 -151
rect -179 -179 -151 -151
rect -113 -179 -85 -151
rect -47 -179 -19 -151
rect 19 -179 47 -151
rect 85 -179 113 -151
rect 151 -179 179 -151
rect 217 -179 245 -151
rect 283 -179 311 -151
rect 349 -179 377 -151
rect 415 -179 443 -151
rect 481 -179 509 -151
rect 547 -179 575 -151
rect 613 -179 641 -151
rect 679 -179 707 -151
rect -707 -245 -679 -217
rect -641 -245 -613 -217
rect -575 -245 -547 -217
rect -509 -245 -481 -217
rect -443 -245 -415 -217
rect -377 -245 -349 -217
rect -311 -245 -283 -217
rect -245 -245 -217 -217
rect -179 -245 -151 -217
rect -113 -245 -85 -217
rect -47 -245 -19 -217
rect 19 -245 47 -217
rect 85 -245 113 -217
rect 151 -245 179 -217
rect 217 -245 245 -217
rect 283 -245 311 -217
rect 349 -245 377 -217
rect 415 -245 443 -217
rect 481 -245 509 -217
rect 547 -245 575 -217
rect 613 -245 641 -217
rect 679 -245 707 -217
rect -707 -311 -679 -283
rect -641 -311 -613 -283
rect -575 -311 -547 -283
rect -509 -311 -481 -283
rect -443 -311 -415 -283
rect -377 -311 -349 -283
rect -311 -311 -283 -283
rect -245 -311 -217 -283
rect -179 -311 -151 -283
rect -113 -311 -85 -283
rect -47 -311 -19 -283
rect 19 -311 47 -283
rect 85 -311 113 -283
rect 151 -311 179 -283
rect 217 -311 245 -283
rect 283 -311 311 -283
rect 349 -311 377 -283
rect 415 -311 443 -283
rect 481 -311 509 -283
rect 547 -311 575 -283
rect 613 -311 641 -283
rect 679 -311 707 -283
<< metal5 >>
rect -715 311 715 319
rect -715 283 -707 311
rect -679 283 -641 311
rect -613 283 -575 311
rect -547 283 -509 311
rect -481 283 -443 311
rect -415 283 -377 311
rect -349 283 -311 311
rect -283 283 -245 311
rect -217 283 -179 311
rect -151 283 -113 311
rect -85 283 -47 311
rect -19 283 19 311
rect 47 283 85 311
rect 113 283 151 311
rect 179 283 217 311
rect 245 283 283 311
rect 311 283 349 311
rect 377 283 415 311
rect 443 283 481 311
rect 509 283 547 311
rect 575 283 613 311
rect 641 283 679 311
rect 707 283 715 311
rect -715 245 715 283
rect -715 217 -707 245
rect -679 217 -641 245
rect -613 217 -575 245
rect -547 217 -509 245
rect -481 217 -443 245
rect -415 217 -377 245
rect -349 217 -311 245
rect -283 217 -245 245
rect -217 217 -179 245
rect -151 217 -113 245
rect -85 217 -47 245
rect -19 217 19 245
rect 47 217 85 245
rect 113 217 151 245
rect 179 217 217 245
rect 245 217 283 245
rect 311 217 349 245
rect 377 217 415 245
rect 443 217 481 245
rect 509 217 547 245
rect 575 217 613 245
rect 641 217 679 245
rect 707 217 715 245
rect -715 179 715 217
rect -715 151 -707 179
rect -679 151 -641 179
rect -613 151 -575 179
rect -547 151 -509 179
rect -481 151 -443 179
rect -415 151 -377 179
rect -349 151 -311 179
rect -283 151 -245 179
rect -217 151 -179 179
rect -151 151 -113 179
rect -85 151 -47 179
rect -19 151 19 179
rect 47 151 85 179
rect 113 151 151 179
rect 179 151 217 179
rect 245 151 283 179
rect 311 151 349 179
rect 377 151 415 179
rect 443 151 481 179
rect 509 151 547 179
rect 575 151 613 179
rect 641 151 679 179
rect 707 151 715 179
rect -715 113 715 151
rect -715 85 -707 113
rect -679 85 -641 113
rect -613 85 -575 113
rect -547 85 -509 113
rect -481 85 -443 113
rect -415 85 -377 113
rect -349 85 -311 113
rect -283 85 -245 113
rect -217 85 -179 113
rect -151 85 -113 113
rect -85 85 -47 113
rect -19 85 19 113
rect 47 85 85 113
rect 113 85 151 113
rect 179 85 217 113
rect 245 85 283 113
rect 311 85 349 113
rect 377 85 415 113
rect 443 85 481 113
rect 509 85 547 113
rect 575 85 613 113
rect 641 85 679 113
rect 707 85 715 113
rect -715 47 715 85
rect -715 19 -707 47
rect -679 19 -641 47
rect -613 19 -575 47
rect -547 19 -509 47
rect -481 19 -443 47
rect -415 19 -377 47
rect -349 19 -311 47
rect -283 19 -245 47
rect -217 19 -179 47
rect -151 19 -113 47
rect -85 19 -47 47
rect -19 19 19 47
rect 47 19 85 47
rect 113 19 151 47
rect 179 19 217 47
rect 245 19 283 47
rect 311 19 349 47
rect 377 19 415 47
rect 443 19 481 47
rect 509 19 547 47
rect 575 19 613 47
rect 641 19 679 47
rect 707 19 715 47
rect -715 -19 715 19
rect -715 -47 -707 -19
rect -679 -47 -641 -19
rect -613 -47 -575 -19
rect -547 -47 -509 -19
rect -481 -47 -443 -19
rect -415 -47 -377 -19
rect -349 -47 -311 -19
rect -283 -47 -245 -19
rect -217 -47 -179 -19
rect -151 -47 -113 -19
rect -85 -47 -47 -19
rect -19 -47 19 -19
rect 47 -47 85 -19
rect 113 -47 151 -19
rect 179 -47 217 -19
rect 245 -47 283 -19
rect 311 -47 349 -19
rect 377 -47 415 -19
rect 443 -47 481 -19
rect 509 -47 547 -19
rect 575 -47 613 -19
rect 641 -47 679 -19
rect 707 -47 715 -19
rect -715 -85 715 -47
rect -715 -113 -707 -85
rect -679 -113 -641 -85
rect -613 -113 -575 -85
rect -547 -113 -509 -85
rect -481 -113 -443 -85
rect -415 -113 -377 -85
rect -349 -113 -311 -85
rect -283 -113 -245 -85
rect -217 -113 -179 -85
rect -151 -113 -113 -85
rect -85 -113 -47 -85
rect -19 -113 19 -85
rect 47 -113 85 -85
rect 113 -113 151 -85
rect 179 -113 217 -85
rect 245 -113 283 -85
rect 311 -113 349 -85
rect 377 -113 415 -85
rect 443 -113 481 -85
rect 509 -113 547 -85
rect 575 -113 613 -85
rect 641 -113 679 -85
rect 707 -113 715 -85
rect -715 -151 715 -113
rect -715 -179 -707 -151
rect -679 -179 -641 -151
rect -613 -179 -575 -151
rect -547 -179 -509 -151
rect -481 -179 -443 -151
rect -415 -179 -377 -151
rect -349 -179 -311 -151
rect -283 -179 -245 -151
rect -217 -179 -179 -151
rect -151 -179 -113 -151
rect -85 -179 -47 -151
rect -19 -179 19 -151
rect 47 -179 85 -151
rect 113 -179 151 -151
rect 179 -179 217 -151
rect 245 -179 283 -151
rect 311 -179 349 -151
rect 377 -179 415 -151
rect 443 -179 481 -151
rect 509 -179 547 -151
rect 575 -179 613 -151
rect 641 -179 679 -151
rect 707 -179 715 -151
rect -715 -217 715 -179
rect -715 -245 -707 -217
rect -679 -245 -641 -217
rect -613 -245 -575 -217
rect -547 -245 -509 -217
rect -481 -245 -443 -217
rect -415 -245 -377 -217
rect -349 -245 -311 -217
rect -283 -245 -245 -217
rect -217 -245 -179 -217
rect -151 -245 -113 -217
rect -85 -245 -47 -217
rect -19 -245 19 -217
rect 47 -245 85 -217
rect 113 -245 151 -217
rect 179 -245 217 -217
rect 245 -245 283 -217
rect 311 -245 349 -217
rect 377 -245 415 -217
rect 443 -245 481 -217
rect 509 -245 547 -217
rect 575 -245 613 -217
rect 641 -245 679 -217
rect 707 -245 715 -217
rect -715 -283 715 -245
rect -715 -311 -707 -283
rect -679 -311 -641 -283
rect -613 -311 -575 -283
rect -547 -311 -509 -283
rect -481 -311 -443 -283
rect -415 -311 -377 -283
rect -349 -311 -311 -283
rect -283 -311 -245 -283
rect -217 -311 -179 -283
rect -151 -311 -113 -283
rect -85 -311 -47 -283
rect -19 -311 19 -283
rect 47 -311 85 -283
rect 113 -311 151 -283
rect 179 -311 217 -283
rect 245 -311 283 -283
rect 311 -311 349 -283
rect 377 -311 415 -283
rect 443 -311 481 -283
rect 509 -311 547 -283
rect 575 -311 613 -283
rect 641 -311 679 -283
rect 707 -311 715 -283
rect -715 -319 715 -311
<< end >>
