magic
tech gf180mcuC
magscale 1 10
timestamp 1692949670
<< error_p >>
rect -3306 -3700 -3182 -3676
rect -1330 -3700 -1206 -3676
rect -3282 -3724 -3206 -3700
rect -1306 -3724 -1230 -3700
rect -2435 -4033 -2373 -3971
rect -3392 -4475 -3327 -4303
rect -3282 -4475 -3256 -4451
rect -3306 -4496 -3256 -4475
rect -3244 -4475 -3206 -4451
rect -2667 -4466 -2621 -4462
rect -2507 -4466 -2461 -4462
rect -2029 -4466 -1983 -4462
rect -1869 -4466 -1823 -4462
rect -1306 -4475 -1276 -4451
rect -3244 -4496 -3108 -4475
rect -3306 -4499 -3108 -4496
rect -1330 -4496 -1276 -4475
rect -1264 -4475 -1230 -4451
rect -1192 -4475 -1128 -4303
rect -1264 -4496 -1128 -4475
rect -1330 -4499 -1128 -4496
rect -3304 -4520 -3108 -4499
rect -1324 -4520 -1128 -4499
rect -3304 -4544 -3196 -4520
rect -1324 -4544 -1216 -4520
<< nwell >>
rect -3327 -4475 -1192 -3700
rect -3280 -4520 -3220 -4475
rect -1300 -4520 -1240 -4475
<< pdiff >>
rect -2435 -4033 -2373 -3971
<< nsubdiff >>
rect -3282 -3722 -3206 -3700
rect -3282 -3768 -3267 -3722
rect -3221 -3768 -3206 -3722
rect -3282 -3816 -3206 -3768
rect -3282 -3862 -3267 -3816
rect -3221 -3862 -3206 -3816
rect -3282 -3910 -3206 -3862
rect -3282 -3956 -3267 -3910
rect -3221 -3956 -3206 -3910
rect -3282 -4004 -3206 -3956
rect -1306 -3722 -1230 -3700
rect -1306 -3768 -1291 -3722
rect -1245 -3768 -1230 -3722
rect -1306 -3816 -1230 -3768
rect -1306 -3862 -1291 -3816
rect -1245 -3862 -1230 -3816
rect -1306 -3910 -1230 -3862
rect -1306 -3956 -1291 -3910
rect -1245 -3956 -1230 -3910
rect -3282 -4050 -3267 -4004
rect -3221 -4050 -3206 -4004
rect -1306 -4004 -1230 -3956
rect -3282 -4098 -3206 -4050
rect -3282 -4144 -3267 -4098
rect -3221 -4144 -3206 -4098
rect -3282 -4192 -3206 -4144
rect -3282 -4238 -3267 -4192
rect -3221 -4238 -3206 -4192
rect -3282 -4286 -3206 -4238
rect -3282 -4332 -3267 -4286
rect -3221 -4332 -3206 -4286
rect -3282 -4380 -3206 -4332
rect -1306 -4050 -1291 -4004
rect -1245 -4050 -1230 -4004
rect -1306 -4098 -1230 -4050
rect -1306 -4144 -1291 -4098
rect -1245 -4144 -1230 -4098
rect -1306 -4192 -1230 -4144
rect -1306 -4238 -1291 -4192
rect -1245 -4238 -1230 -4192
rect -1306 -4286 -1230 -4238
rect -1306 -4332 -1291 -4286
rect -1245 -4332 -1230 -4286
rect -3282 -4426 -3267 -4380
rect -3221 -4426 -3206 -4380
rect -3282 -4475 -3206 -4426
rect -1306 -4380 -1230 -4332
rect -1306 -4426 -1291 -4380
rect -1245 -4426 -1230 -4380
rect -1306 -4475 -1230 -4426
rect -3280 -4520 -3220 -4475
rect -1300 -4520 -1240 -4475
<< nsubdiffcont >>
rect -3267 -3768 -3221 -3722
rect -3267 -3862 -3221 -3816
rect -3267 -3956 -3221 -3910
rect -1291 -3768 -1245 -3722
rect -1291 -3862 -1245 -3816
rect -1291 -3956 -1245 -3910
rect -3267 -4050 -3221 -4004
rect -3267 -4144 -3221 -4098
rect -3267 -4238 -3221 -4192
rect -3267 -4332 -3221 -4286
rect -1291 -4050 -1245 -4004
rect -1291 -4144 -1245 -4098
rect -1291 -4238 -1245 -4192
rect -1291 -4332 -1245 -4286
rect -3267 -4426 -3221 -4380
rect -1291 -4426 -1245 -4380
<< polysilicon >>
rect -3086 -4380 -2937 -4361
rect -3086 -4426 -3068 -4380
rect -3022 -4426 -2937 -4380
rect -2673 -4402 -2617 -4361
rect -3086 -4453 -2937 -4426
rect -2688 -4420 -2601 -4402
rect -2513 -4403 -2457 -4361
rect -2033 -4403 -1977 -4361
rect -1873 -4402 -1817 -4361
rect -1553 -4381 -1396 -4361
rect -2688 -4466 -2667 -4420
rect -2621 -4466 -2601 -4420
rect -2688 -4475 -2601 -4466
rect -2529 -4420 -2442 -4403
rect -2529 -4466 -2507 -4420
rect -2461 -4466 -2442 -4420
rect -2529 -4475 -2442 -4466
rect -2048 -4420 -1961 -4403
rect -2048 -4466 -2029 -4420
rect -1983 -4466 -1961 -4420
rect -2048 -4475 -1961 -4466
rect -1889 -4420 -1802 -4402
rect -1889 -4466 -1869 -4420
rect -1823 -4466 -1802 -4420
rect -1553 -4427 -1468 -4381
rect -1422 -4427 -1396 -4381
rect -1553 -4448 -1396 -4427
rect -1889 -4475 -1802 -4466
<< polycontact >>
rect -3068 -4426 -3022 -4380
rect -2667 -4466 -2621 -4420
rect -2507 -4466 -2461 -4420
rect -2029 -4466 -1983 -4420
rect -1869 -4466 -1823 -4420
rect -1468 -4427 -1422 -4381
<< metal1 >>
rect -3293 -3722 -3195 -3700
rect -3293 -3768 -3267 -3722
rect -3221 -3768 -3195 -3722
rect -3293 -3816 -3195 -3768
rect -1317 -3722 -1219 -3700
rect -1317 -3768 -1291 -3722
rect -1245 -3768 -1219 -3722
rect -3293 -3862 -3267 -3816
rect -3221 -3862 -3195 -3816
rect -3293 -3910 -3195 -3862
rect -2607 -3822 -2524 -3808
rect -2607 -3878 -2593 -3822
rect -2537 -3878 -2524 -3822
rect -2607 -3890 -2524 -3878
rect -1965 -3822 -1882 -3809
rect -1965 -3878 -1952 -3822
rect -1896 -3878 -1882 -3822
rect -1965 -3891 -1882 -3878
rect -1317 -3816 -1219 -3768
rect -1317 -3862 -1291 -3816
rect -1245 -3862 -1219 -3816
rect -3293 -3956 -3267 -3910
rect -3221 -3956 -3195 -3910
rect -3293 -4004 -3195 -3956
rect -1317 -3910 -1219 -3862
rect -1317 -3956 -1291 -3910
rect -1245 -3956 -1219 -3910
rect -3293 -4050 -3267 -4004
rect -3221 -4050 -3195 -4004
rect -2767 -3975 -2684 -3961
rect -2767 -4031 -2753 -3975
rect -2697 -4031 -2684 -3975
rect -2767 -4043 -2684 -4031
rect -2446 -3971 -2363 -3960
rect -2446 -4033 -2435 -3971
rect -2373 -4033 -2363 -3971
rect -2446 -4042 -2363 -4033
rect -2126 -3974 -2043 -3960
rect -2126 -4030 -2112 -3974
rect -2056 -4030 -2043 -3974
rect -2126 -4042 -2043 -4030
rect -1806 -3975 -1723 -3961
rect -1806 -4031 -1792 -3975
rect -1736 -4031 -1723 -3975
rect -1806 -4043 -1723 -4031
rect -1317 -4004 -1219 -3956
rect -3293 -4098 -3195 -4050
rect -3293 -4144 -3267 -4098
rect -3221 -4144 -3195 -4098
rect -1317 -4050 -1291 -4004
rect -1245 -4050 -1219 -4004
rect -1317 -4098 -1219 -4050
rect -3293 -4192 -3195 -4144
rect -3293 -4238 -3267 -4192
rect -3221 -4238 -3195 -4192
rect -3088 -4134 -3004 -4120
rect -3088 -4190 -3074 -4134
rect -3018 -4190 -3004 -4134
rect -3088 -4204 -3004 -4190
rect -2927 -4134 -2843 -4119
rect -2927 -4190 -2913 -4134
rect -2857 -4190 -2843 -4134
rect -2927 -4203 -2843 -4190
rect -2288 -4134 -2202 -4120
rect -2288 -4190 -2274 -4134
rect -2216 -4190 -2202 -4134
rect -2288 -4204 -2202 -4190
rect -1647 -4134 -1563 -4119
rect -1647 -4190 -1633 -4134
rect -1577 -4190 -1563 -4134
rect -1647 -4203 -1563 -4190
rect -1487 -4134 -1403 -4120
rect -1487 -4190 -1473 -4134
rect -1417 -4190 -1403 -4134
rect -1487 -4204 -1403 -4190
rect -1317 -4144 -1291 -4098
rect -1245 -4121 -1219 -4098
rect -1245 -4144 -1142 -4121
rect -1317 -4192 -1142 -4144
rect -3293 -4286 -3195 -4238
rect -3293 -4332 -3267 -4286
rect -3221 -4332 -3195 -4286
rect -1317 -4238 -1291 -4192
rect -1245 -4238 -1142 -4192
rect -1317 -4268 -1142 -4238
rect -1317 -4286 -1219 -4268
rect -3293 -4380 -3195 -4332
rect -3068 -4373 -3022 -4315
rect -1468 -4369 -1422 -4315
rect -1317 -4332 -1291 -4286
rect -1245 -4332 -1219 -4286
rect -3293 -4426 -3267 -4380
rect -3221 -4426 -3195 -4380
rect -3293 -4475 -3195 -4426
rect -3080 -4380 -3010 -4373
rect -3080 -4426 -3068 -4380
rect -3022 -4426 -3010 -4380
rect -1480 -4381 -1410 -4369
rect -1745 -4407 -1644 -4386
rect -1745 -4415 -1724 -4407
rect -3080 -4439 -3010 -4426
rect -2688 -4420 -1724 -4415
rect -2688 -4466 -2667 -4420
rect -2621 -4466 -2507 -4420
rect -2461 -4466 -2029 -4420
rect -1983 -4466 -1869 -4420
rect -1823 -4463 -1724 -4420
rect -1668 -4463 -1644 -4407
rect -1480 -4427 -1468 -4381
rect -1422 -4427 -1410 -4381
rect -1480 -4439 -1410 -4427
rect -1317 -4380 -1219 -4332
rect -1317 -4426 -1291 -4380
rect -1245 -4426 -1219 -4380
rect -1823 -4466 -1644 -4463
rect -2688 -4471 -1644 -4466
rect -1745 -4475 -1644 -4471
rect -1317 -4475 -1219 -4426
rect -3280 -4520 -3220 -4475
rect -1300 -4520 -1240 -4475
<< via1 >>
rect -2593 -3878 -2537 -3822
rect -1952 -3878 -1896 -3822
rect -2753 -4031 -2697 -3975
rect -2435 -4033 -2373 -3971
rect -2112 -4030 -2056 -3974
rect -1792 -4031 -1736 -3975
rect -3074 -4190 -3018 -4134
rect -2913 -4190 -2857 -4134
rect -2274 -4190 -2216 -4134
rect -1633 -4190 -1577 -4134
rect -1473 -4190 -1417 -4134
rect -1724 -4463 -1668 -4407
<< metal2 >>
rect -3472 -3973 -3352 -3700
rect -2524 -3808 -2332 -3806
rect -2607 -3819 -2332 -3808
rect -2607 -3822 -2510 -3819
rect -2607 -3878 -2593 -3822
rect -2537 -3875 -2510 -3822
rect -2454 -3875 -2400 -3819
rect -2344 -3820 -2332 -3819
rect -1965 -3820 -1882 -3809
rect -2344 -3822 -1882 -3820
rect -2344 -3875 -1952 -3822
rect -2537 -3878 -1952 -3875
rect -1896 -3878 -1882 -3822
rect -2607 -3880 -1882 -3878
rect -2607 -3890 -2332 -3880
rect -1965 -3891 -1882 -3880
rect -2767 -3973 -2684 -3961
rect -2446 -3971 -2363 -3960
rect -2446 -3973 -2435 -3971
rect -3472 -3975 -2435 -3973
rect -3472 -4031 -2753 -3975
rect -2697 -4031 -2435 -3975
rect -3472 -4033 -2435 -4031
rect -2373 -3973 -2363 -3971
rect -2126 -3973 -2043 -3960
rect -1806 -3973 -1723 -3961
rect -2373 -3974 -1723 -3973
rect -2373 -4030 -2112 -3974
rect -2056 -3975 -1723 -3974
rect -2056 -4030 -1792 -3975
rect -2373 -4031 -1792 -4030
rect -1736 -4031 -1723 -3975
rect -2373 -4033 -1723 -4031
rect -3472 -4034 -1723 -4033
rect -3472 -4475 -3352 -4034
rect -2767 -4043 -2684 -4034
rect -2446 -4042 -2363 -4034
rect -2126 -4042 -2043 -4034
rect -1806 -4043 -1723 -4034
rect -3088 -4132 -3004 -4120
rect -2927 -4132 -2843 -4119
rect -2288 -4132 -2202 -4120
rect -2121 -4131 -1929 -4118
rect -2121 -4132 -2107 -4131
rect -3088 -4134 -2107 -4132
rect -3088 -4190 -3074 -4134
rect -3018 -4190 -2913 -4134
rect -2857 -4190 -2274 -4134
rect -2216 -4187 -2107 -4134
rect -2051 -4187 -1997 -4131
rect -1941 -4132 -1929 -4131
rect -1647 -4132 -1563 -4119
rect -1487 -4132 -1403 -4120
rect -1941 -4134 -1403 -4132
rect -1941 -4187 -1633 -4134
rect -2216 -4190 -1633 -4187
rect -1577 -4190 -1473 -4134
rect -1417 -4190 -1403 -4134
rect -3088 -4192 -1403 -4190
rect -3088 -4204 -3004 -4192
rect -2927 -4203 -2843 -4192
rect -2288 -4204 -2202 -4192
rect -2121 -4202 -1929 -4192
rect -1647 -4203 -1563 -4192
rect -1487 -4204 -1403 -4192
rect -1745 -4407 -1644 -4386
rect -1745 -4463 -1724 -4407
rect -1668 -4463 -1644 -4407
rect -1745 -4475 -1644 -4463
<< via2 >>
rect -2510 -3875 -2454 -3819
rect -2400 -3875 -2344 -3819
rect -2107 -4187 -2051 -4131
rect -1997 -4187 -1941 -4131
rect -1724 -4463 -1668 -4407
<< metal3 >>
rect -2833 -4475 -2767 -3700
rect -2458 -3806 -2392 -3700
rect -2524 -3819 -2332 -3806
rect -2524 -3875 -2510 -3819
rect -2454 -3875 -2400 -3819
rect -2344 -3875 -2332 -3819
rect -2524 -3890 -2332 -3875
rect -2458 -4475 -2392 -3890
rect -2097 -4118 -2031 -3700
rect -2121 -4131 -1929 -4118
rect -2121 -4187 -2107 -4131
rect -2051 -4187 -1997 -4131
rect -1941 -4187 -1929 -4131
rect -2121 -4202 -1929 -4187
rect -2097 -4475 -2031 -4202
rect -1726 -4386 -1660 -3700
rect -1745 -4407 -1644 -4386
rect -1745 -4463 -1724 -4407
rect -1668 -4463 -1644 -4407
rect -1745 -4475 -1644 -4463
<< end >>
