magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -5573 -1745 5573 1745
<< metal3 >>
rect -4573 740 4573 745
rect -4573 712 -4568 740
rect -4540 712 -4502 740
rect -4474 712 -4436 740
rect -4408 712 -4370 740
rect -4342 712 -4304 740
rect -4276 712 -4238 740
rect -4210 712 -4172 740
rect -4144 712 -4106 740
rect -4078 712 -4040 740
rect -4012 712 -3974 740
rect -3946 712 -3908 740
rect -3880 712 -3842 740
rect -3814 712 -3776 740
rect -3748 712 -3710 740
rect -3682 712 -3644 740
rect -3616 712 -3578 740
rect -3550 712 -3512 740
rect -3484 712 -3446 740
rect -3418 712 -3380 740
rect -3352 712 -3314 740
rect -3286 712 -3248 740
rect -3220 712 -3182 740
rect -3154 712 -3116 740
rect -3088 712 -3050 740
rect -3022 712 -2984 740
rect -2956 712 -2918 740
rect -2890 712 -2852 740
rect -2824 712 -2786 740
rect -2758 712 -2720 740
rect -2692 712 -2654 740
rect -2626 712 -2588 740
rect -2560 712 -2522 740
rect -2494 712 -2456 740
rect -2428 712 -2390 740
rect -2362 712 -2324 740
rect -2296 712 -2258 740
rect -2230 712 -2192 740
rect -2164 712 -2126 740
rect -2098 712 -2060 740
rect -2032 712 -1994 740
rect -1966 712 -1928 740
rect -1900 712 -1862 740
rect -1834 712 -1796 740
rect -1768 712 -1730 740
rect -1702 712 -1664 740
rect -1636 712 -1598 740
rect -1570 712 -1532 740
rect -1504 712 -1466 740
rect -1438 712 -1400 740
rect -1372 712 -1334 740
rect -1306 712 -1268 740
rect -1240 712 -1202 740
rect -1174 712 -1136 740
rect -1108 712 -1070 740
rect -1042 712 -1004 740
rect -976 712 -938 740
rect -910 712 -872 740
rect -844 712 -806 740
rect -778 712 -740 740
rect -712 712 -674 740
rect -646 712 -608 740
rect -580 712 -542 740
rect -514 712 -476 740
rect -448 712 -410 740
rect -382 712 -344 740
rect -316 712 -278 740
rect -250 712 -212 740
rect -184 712 -146 740
rect -118 712 -80 740
rect -52 712 -14 740
rect 14 712 52 740
rect 80 712 118 740
rect 146 712 184 740
rect 212 712 250 740
rect 278 712 316 740
rect 344 712 382 740
rect 410 712 448 740
rect 476 712 514 740
rect 542 712 580 740
rect 608 712 646 740
rect 674 712 712 740
rect 740 712 778 740
rect 806 712 844 740
rect 872 712 910 740
rect 938 712 976 740
rect 1004 712 1042 740
rect 1070 712 1108 740
rect 1136 712 1174 740
rect 1202 712 1240 740
rect 1268 712 1306 740
rect 1334 712 1372 740
rect 1400 712 1438 740
rect 1466 712 1504 740
rect 1532 712 1570 740
rect 1598 712 1636 740
rect 1664 712 1702 740
rect 1730 712 1768 740
rect 1796 712 1834 740
rect 1862 712 1900 740
rect 1928 712 1966 740
rect 1994 712 2032 740
rect 2060 712 2098 740
rect 2126 712 2164 740
rect 2192 712 2230 740
rect 2258 712 2296 740
rect 2324 712 2362 740
rect 2390 712 2428 740
rect 2456 712 2494 740
rect 2522 712 2560 740
rect 2588 712 2626 740
rect 2654 712 2692 740
rect 2720 712 2758 740
rect 2786 712 2824 740
rect 2852 712 2890 740
rect 2918 712 2956 740
rect 2984 712 3022 740
rect 3050 712 3088 740
rect 3116 712 3154 740
rect 3182 712 3220 740
rect 3248 712 3286 740
rect 3314 712 3352 740
rect 3380 712 3418 740
rect 3446 712 3484 740
rect 3512 712 3550 740
rect 3578 712 3616 740
rect 3644 712 3682 740
rect 3710 712 3748 740
rect 3776 712 3814 740
rect 3842 712 3880 740
rect 3908 712 3946 740
rect 3974 712 4012 740
rect 4040 712 4078 740
rect 4106 712 4144 740
rect 4172 712 4210 740
rect 4238 712 4276 740
rect 4304 712 4342 740
rect 4370 712 4408 740
rect 4436 712 4474 740
rect 4502 712 4540 740
rect 4568 712 4573 740
rect -4573 674 4573 712
rect -4573 646 -4568 674
rect -4540 646 -4502 674
rect -4474 646 -4436 674
rect -4408 646 -4370 674
rect -4342 646 -4304 674
rect -4276 646 -4238 674
rect -4210 646 -4172 674
rect -4144 646 -4106 674
rect -4078 646 -4040 674
rect -4012 646 -3974 674
rect -3946 646 -3908 674
rect -3880 646 -3842 674
rect -3814 646 -3776 674
rect -3748 646 -3710 674
rect -3682 646 -3644 674
rect -3616 646 -3578 674
rect -3550 646 -3512 674
rect -3484 646 -3446 674
rect -3418 646 -3380 674
rect -3352 646 -3314 674
rect -3286 646 -3248 674
rect -3220 646 -3182 674
rect -3154 646 -3116 674
rect -3088 646 -3050 674
rect -3022 646 -2984 674
rect -2956 646 -2918 674
rect -2890 646 -2852 674
rect -2824 646 -2786 674
rect -2758 646 -2720 674
rect -2692 646 -2654 674
rect -2626 646 -2588 674
rect -2560 646 -2522 674
rect -2494 646 -2456 674
rect -2428 646 -2390 674
rect -2362 646 -2324 674
rect -2296 646 -2258 674
rect -2230 646 -2192 674
rect -2164 646 -2126 674
rect -2098 646 -2060 674
rect -2032 646 -1994 674
rect -1966 646 -1928 674
rect -1900 646 -1862 674
rect -1834 646 -1796 674
rect -1768 646 -1730 674
rect -1702 646 -1664 674
rect -1636 646 -1598 674
rect -1570 646 -1532 674
rect -1504 646 -1466 674
rect -1438 646 -1400 674
rect -1372 646 -1334 674
rect -1306 646 -1268 674
rect -1240 646 -1202 674
rect -1174 646 -1136 674
rect -1108 646 -1070 674
rect -1042 646 -1004 674
rect -976 646 -938 674
rect -910 646 -872 674
rect -844 646 -806 674
rect -778 646 -740 674
rect -712 646 -674 674
rect -646 646 -608 674
rect -580 646 -542 674
rect -514 646 -476 674
rect -448 646 -410 674
rect -382 646 -344 674
rect -316 646 -278 674
rect -250 646 -212 674
rect -184 646 -146 674
rect -118 646 -80 674
rect -52 646 -14 674
rect 14 646 52 674
rect 80 646 118 674
rect 146 646 184 674
rect 212 646 250 674
rect 278 646 316 674
rect 344 646 382 674
rect 410 646 448 674
rect 476 646 514 674
rect 542 646 580 674
rect 608 646 646 674
rect 674 646 712 674
rect 740 646 778 674
rect 806 646 844 674
rect 872 646 910 674
rect 938 646 976 674
rect 1004 646 1042 674
rect 1070 646 1108 674
rect 1136 646 1174 674
rect 1202 646 1240 674
rect 1268 646 1306 674
rect 1334 646 1372 674
rect 1400 646 1438 674
rect 1466 646 1504 674
rect 1532 646 1570 674
rect 1598 646 1636 674
rect 1664 646 1702 674
rect 1730 646 1768 674
rect 1796 646 1834 674
rect 1862 646 1900 674
rect 1928 646 1966 674
rect 1994 646 2032 674
rect 2060 646 2098 674
rect 2126 646 2164 674
rect 2192 646 2230 674
rect 2258 646 2296 674
rect 2324 646 2362 674
rect 2390 646 2428 674
rect 2456 646 2494 674
rect 2522 646 2560 674
rect 2588 646 2626 674
rect 2654 646 2692 674
rect 2720 646 2758 674
rect 2786 646 2824 674
rect 2852 646 2890 674
rect 2918 646 2956 674
rect 2984 646 3022 674
rect 3050 646 3088 674
rect 3116 646 3154 674
rect 3182 646 3220 674
rect 3248 646 3286 674
rect 3314 646 3352 674
rect 3380 646 3418 674
rect 3446 646 3484 674
rect 3512 646 3550 674
rect 3578 646 3616 674
rect 3644 646 3682 674
rect 3710 646 3748 674
rect 3776 646 3814 674
rect 3842 646 3880 674
rect 3908 646 3946 674
rect 3974 646 4012 674
rect 4040 646 4078 674
rect 4106 646 4144 674
rect 4172 646 4210 674
rect 4238 646 4276 674
rect 4304 646 4342 674
rect 4370 646 4408 674
rect 4436 646 4474 674
rect 4502 646 4540 674
rect 4568 646 4573 674
rect -4573 608 4573 646
rect -4573 580 -4568 608
rect -4540 580 -4502 608
rect -4474 580 -4436 608
rect -4408 580 -4370 608
rect -4342 580 -4304 608
rect -4276 580 -4238 608
rect -4210 580 -4172 608
rect -4144 580 -4106 608
rect -4078 580 -4040 608
rect -4012 580 -3974 608
rect -3946 580 -3908 608
rect -3880 580 -3842 608
rect -3814 580 -3776 608
rect -3748 580 -3710 608
rect -3682 580 -3644 608
rect -3616 580 -3578 608
rect -3550 580 -3512 608
rect -3484 580 -3446 608
rect -3418 580 -3380 608
rect -3352 580 -3314 608
rect -3286 580 -3248 608
rect -3220 580 -3182 608
rect -3154 580 -3116 608
rect -3088 580 -3050 608
rect -3022 580 -2984 608
rect -2956 580 -2918 608
rect -2890 580 -2852 608
rect -2824 580 -2786 608
rect -2758 580 -2720 608
rect -2692 580 -2654 608
rect -2626 580 -2588 608
rect -2560 580 -2522 608
rect -2494 580 -2456 608
rect -2428 580 -2390 608
rect -2362 580 -2324 608
rect -2296 580 -2258 608
rect -2230 580 -2192 608
rect -2164 580 -2126 608
rect -2098 580 -2060 608
rect -2032 580 -1994 608
rect -1966 580 -1928 608
rect -1900 580 -1862 608
rect -1834 580 -1796 608
rect -1768 580 -1730 608
rect -1702 580 -1664 608
rect -1636 580 -1598 608
rect -1570 580 -1532 608
rect -1504 580 -1466 608
rect -1438 580 -1400 608
rect -1372 580 -1334 608
rect -1306 580 -1268 608
rect -1240 580 -1202 608
rect -1174 580 -1136 608
rect -1108 580 -1070 608
rect -1042 580 -1004 608
rect -976 580 -938 608
rect -910 580 -872 608
rect -844 580 -806 608
rect -778 580 -740 608
rect -712 580 -674 608
rect -646 580 -608 608
rect -580 580 -542 608
rect -514 580 -476 608
rect -448 580 -410 608
rect -382 580 -344 608
rect -316 580 -278 608
rect -250 580 -212 608
rect -184 580 -146 608
rect -118 580 -80 608
rect -52 580 -14 608
rect 14 580 52 608
rect 80 580 118 608
rect 146 580 184 608
rect 212 580 250 608
rect 278 580 316 608
rect 344 580 382 608
rect 410 580 448 608
rect 476 580 514 608
rect 542 580 580 608
rect 608 580 646 608
rect 674 580 712 608
rect 740 580 778 608
rect 806 580 844 608
rect 872 580 910 608
rect 938 580 976 608
rect 1004 580 1042 608
rect 1070 580 1108 608
rect 1136 580 1174 608
rect 1202 580 1240 608
rect 1268 580 1306 608
rect 1334 580 1372 608
rect 1400 580 1438 608
rect 1466 580 1504 608
rect 1532 580 1570 608
rect 1598 580 1636 608
rect 1664 580 1702 608
rect 1730 580 1768 608
rect 1796 580 1834 608
rect 1862 580 1900 608
rect 1928 580 1966 608
rect 1994 580 2032 608
rect 2060 580 2098 608
rect 2126 580 2164 608
rect 2192 580 2230 608
rect 2258 580 2296 608
rect 2324 580 2362 608
rect 2390 580 2428 608
rect 2456 580 2494 608
rect 2522 580 2560 608
rect 2588 580 2626 608
rect 2654 580 2692 608
rect 2720 580 2758 608
rect 2786 580 2824 608
rect 2852 580 2890 608
rect 2918 580 2956 608
rect 2984 580 3022 608
rect 3050 580 3088 608
rect 3116 580 3154 608
rect 3182 580 3220 608
rect 3248 580 3286 608
rect 3314 580 3352 608
rect 3380 580 3418 608
rect 3446 580 3484 608
rect 3512 580 3550 608
rect 3578 580 3616 608
rect 3644 580 3682 608
rect 3710 580 3748 608
rect 3776 580 3814 608
rect 3842 580 3880 608
rect 3908 580 3946 608
rect 3974 580 4012 608
rect 4040 580 4078 608
rect 4106 580 4144 608
rect 4172 580 4210 608
rect 4238 580 4276 608
rect 4304 580 4342 608
rect 4370 580 4408 608
rect 4436 580 4474 608
rect 4502 580 4540 608
rect 4568 580 4573 608
rect -4573 542 4573 580
rect -4573 514 -4568 542
rect -4540 514 -4502 542
rect -4474 514 -4436 542
rect -4408 514 -4370 542
rect -4342 514 -4304 542
rect -4276 514 -4238 542
rect -4210 514 -4172 542
rect -4144 514 -4106 542
rect -4078 514 -4040 542
rect -4012 514 -3974 542
rect -3946 514 -3908 542
rect -3880 514 -3842 542
rect -3814 514 -3776 542
rect -3748 514 -3710 542
rect -3682 514 -3644 542
rect -3616 514 -3578 542
rect -3550 514 -3512 542
rect -3484 514 -3446 542
rect -3418 514 -3380 542
rect -3352 514 -3314 542
rect -3286 514 -3248 542
rect -3220 514 -3182 542
rect -3154 514 -3116 542
rect -3088 514 -3050 542
rect -3022 514 -2984 542
rect -2956 514 -2918 542
rect -2890 514 -2852 542
rect -2824 514 -2786 542
rect -2758 514 -2720 542
rect -2692 514 -2654 542
rect -2626 514 -2588 542
rect -2560 514 -2522 542
rect -2494 514 -2456 542
rect -2428 514 -2390 542
rect -2362 514 -2324 542
rect -2296 514 -2258 542
rect -2230 514 -2192 542
rect -2164 514 -2126 542
rect -2098 514 -2060 542
rect -2032 514 -1994 542
rect -1966 514 -1928 542
rect -1900 514 -1862 542
rect -1834 514 -1796 542
rect -1768 514 -1730 542
rect -1702 514 -1664 542
rect -1636 514 -1598 542
rect -1570 514 -1532 542
rect -1504 514 -1466 542
rect -1438 514 -1400 542
rect -1372 514 -1334 542
rect -1306 514 -1268 542
rect -1240 514 -1202 542
rect -1174 514 -1136 542
rect -1108 514 -1070 542
rect -1042 514 -1004 542
rect -976 514 -938 542
rect -910 514 -872 542
rect -844 514 -806 542
rect -778 514 -740 542
rect -712 514 -674 542
rect -646 514 -608 542
rect -580 514 -542 542
rect -514 514 -476 542
rect -448 514 -410 542
rect -382 514 -344 542
rect -316 514 -278 542
rect -250 514 -212 542
rect -184 514 -146 542
rect -118 514 -80 542
rect -52 514 -14 542
rect 14 514 52 542
rect 80 514 118 542
rect 146 514 184 542
rect 212 514 250 542
rect 278 514 316 542
rect 344 514 382 542
rect 410 514 448 542
rect 476 514 514 542
rect 542 514 580 542
rect 608 514 646 542
rect 674 514 712 542
rect 740 514 778 542
rect 806 514 844 542
rect 872 514 910 542
rect 938 514 976 542
rect 1004 514 1042 542
rect 1070 514 1108 542
rect 1136 514 1174 542
rect 1202 514 1240 542
rect 1268 514 1306 542
rect 1334 514 1372 542
rect 1400 514 1438 542
rect 1466 514 1504 542
rect 1532 514 1570 542
rect 1598 514 1636 542
rect 1664 514 1702 542
rect 1730 514 1768 542
rect 1796 514 1834 542
rect 1862 514 1900 542
rect 1928 514 1966 542
rect 1994 514 2032 542
rect 2060 514 2098 542
rect 2126 514 2164 542
rect 2192 514 2230 542
rect 2258 514 2296 542
rect 2324 514 2362 542
rect 2390 514 2428 542
rect 2456 514 2494 542
rect 2522 514 2560 542
rect 2588 514 2626 542
rect 2654 514 2692 542
rect 2720 514 2758 542
rect 2786 514 2824 542
rect 2852 514 2890 542
rect 2918 514 2956 542
rect 2984 514 3022 542
rect 3050 514 3088 542
rect 3116 514 3154 542
rect 3182 514 3220 542
rect 3248 514 3286 542
rect 3314 514 3352 542
rect 3380 514 3418 542
rect 3446 514 3484 542
rect 3512 514 3550 542
rect 3578 514 3616 542
rect 3644 514 3682 542
rect 3710 514 3748 542
rect 3776 514 3814 542
rect 3842 514 3880 542
rect 3908 514 3946 542
rect 3974 514 4012 542
rect 4040 514 4078 542
rect 4106 514 4144 542
rect 4172 514 4210 542
rect 4238 514 4276 542
rect 4304 514 4342 542
rect 4370 514 4408 542
rect 4436 514 4474 542
rect 4502 514 4540 542
rect 4568 514 4573 542
rect -4573 476 4573 514
rect -4573 448 -4568 476
rect -4540 448 -4502 476
rect -4474 448 -4436 476
rect -4408 448 -4370 476
rect -4342 448 -4304 476
rect -4276 448 -4238 476
rect -4210 448 -4172 476
rect -4144 448 -4106 476
rect -4078 448 -4040 476
rect -4012 448 -3974 476
rect -3946 448 -3908 476
rect -3880 448 -3842 476
rect -3814 448 -3776 476
rect -3748 448 -3710 476
rect -3682 448 -3644 476
rect -3616 448 -3578 476
rect -3550 448 -3512 476
rect -3484 448 -3446 476
rect -3418 448 -3380 476
rect -3352 448 -3314 476
rect -3286 448 -3248 476
rect -3220 448 -3182 476
rect -3154 448 -3116 476
rect -3088 448 -3050 476
rect -3022 448 -2984 476
rect -2956 448 -2918 476
rect -2890 448 -2852 476
rect -2824 448 -2786 476
rect -2758 448 -2720 476
rect -2692 448 -2654 476
rect -2626 448 -2588 476
rect -2560 448 -2522 476
rect -2494 448 -2456 476
rect -2428 448 -2390 476
rect -2362 448 -2324 476
rect -2296 448 -2258 476
rect -2230 448 -2192 476
rect -2164 448 -2126 476
rect -2098 448 -2060 476
rect -2032 448 -1994 476
rect -1966 448 -1928 476
rect -1900 448 -1862 476
rect -1834 448 -1796 476
rect -1768 448 -1730 476
rect -1702 448 -1664 476
rect -1636 448 -1598 476
rect -1570 448 -1532 476
rect -1504 448 -1466 476
rect -1438 448 -1400 476
rect -1372 448 -1334 476
rect -1306 448 -1268 476
rect -1240 448 -1202 476
rect -1174 448 -1136 476
rect -1108 448 -1070 476
rect -1042 448 -1004 476
rect -976 448 -938 476
rect -910 448 -872 476
rect -844 448 -806 476
rect -778 448 -740 476
rect -712 448 -674 476
rect -646 448 -608 476
rect -580 448 -542 476
rect -514 448 -476 476
rect -448 448 -410 476
rect -382 448 -344 476
rect -316 448 -278 476
rect -250 448 -212 476
rect -184 448 -146 476
rect -118 448 -80 476
rect -52 448 -14 476
rect 14 448 52 476
rect 80 448 118 476
rect 146 448 184 476
rect 212 448 250 476
rect 278 448 316 476
rect 344 448 382 476
rect 410 448 448 476
rect 476 448 514 476
rect 542 448 580 476
rect 608 448 646 476
rect 674 448 712 476
rect 740 448 778 476
rect 806 448 844 476
rect 872 448 910 476
rect 938 448 976 476
rect 1004 448 1042 476
rect 1070 448 1108 476
rect 1136 448 1174 476
rect 1202 448 1240 476
rect 1268 448 1306 476
rect 1334 448 1372 476
rect 1400 448 1438 476
rect 1466 448 1504 476
rect 1532 448 1570 476
rect 1598 448 1636 476
rect 1664 448 1702 476
rect 1730 448 1768 476
rect 1796 448 1834 476
rect 1862 448 1900 476
rect 1928 448 1966 476
rect 1994 448 2032 476
rect 2060 448 2098 476
rect 2126 448 2164 476
rect 2192 448 2230 476
rect 2258 448 2296 476
rect 2324 448 2362 476
rect 2390 448 2428 476
rect 2456 448 2494 476
rect 2522 448 2560 476
rect 2588 448 2626 476
rect 2654 448 2692 476
rect 2720 448 2758 476
rect 2786 448 2824 476
rect 2852 448 2890 476
rect 2918 448 2956 476
rect 2984 448 3022 476
rect 3050 448 3088 476
rect 3116 448 3154 476
rect 3182 448 3220 476
rect 3248 448 3286 476
rect 3314 448 3352 476
rect 3380 448 3418 476
rect 3446 448 3484 476
rect 3512 448 3550 476
rect 3578 448 3616 476
rect 3644 448 3682 476
rect 3710 448 3748 476
rect 3776 448 3814 476
rect 3842 448 3880 476
rect 3908 448 3946 476
rect 3974 448 4012 476
rect 4040 448 4078 476
rect 4106 448 4144 476
rect 4172 448 4210 476
rect 4238 448 4276 476
rect 4304 448 4342 476
rect 4370 448 4408 476
rect 4436 448 4474 476
rect 4502 448 4540 476
rect 4568 448 4573 476
rect -4573 410 4573 448
rect -4573 382 -4568 410
rect -4540 382 -4502 410
rect -4474 382 -4436 410
rect -4408 382 -4370 410
rect -4342 382 -4304 410
rect -4276 382 -4238 410
rect -4210 382 -4172 410
rect -4144 382 -4106 410
rect -4078 382 -4040 410
rect -4012 382 -3974 410
rect -3946 382 -3908 410
rect -3880 382 -3842 410
rect -3814 382 -3776 410
rect -3748 382 -3710 410
rect -3682 382 -3644 410
rect -3616 382 -3578 410
rect -3550 382 -3512 410
rect -3484 382 -3446 410
rect -3418 382 -3380 410
rect -3352 382 -3314 410
rect -3286 382 -3248 410
rect -3220 382 -3182 410
rect -3154 382 -3116 410
rect -3088 382 -3050 410
rect -3022 382 -2984 410
rect -2956 382 -2918 410
rect -2890 382 -2852 410
rect -2824 382 -2786 410
rect -2758 382 -2720 410
rect -2692 382 -2654 410
rect -2626 382 -2588 410
rect -2560 382 -2522 410
rect -2494 382 -2456 410
rect -2428 382 -2390 410
rect -2362 382 -2324 410
rect -2296 382 -2258 410
rect -2230 382 -2192 410
rect -2164 382 -2126 410
rect -2098 382 -2060 410
rect -2032 382 -1994 410
rect -1966 382 -1928 410
rect -1900 382 -1862 410
rect -1834 382 -1796 410
rect -1768 382 -1730 410
rect -1702 382 -1664 410
rect -1636 382 -1598 410
rect -1570 382 -1532 410
rect -1504 382 -1466 410
rect -1438 382 -1400 410
rect -1372 382 -1334 410
rect -1306 382 -1268 410
rect -1240 382 -1202 410
rect -1174 382 -1136 410
rect -1108 382 -1070 410
rect -1042 382 -1004 410
rect -976 382 -938 410
rect -910 382 -872 410
rect -844 382 -806 410
rect -778 382 -740 410
rect -712 382 -674 410
rect -646 382 -608 410
rect -580 382 -542 410
rect -514 382 -476 410
rect -448 382 -410 410
rect -382 382 -344 410
rect -316 382 -278 410
rect -250 382 -212 410
rect -184 382 -146 410
rect -118 382 -80 410
rect -52 382 -14 410
rect 14 382 52 410
rect 80 382 118 410
rect 146 382 184 410
rect 212 382 250 410
rect 278 382 316 410
rect 344 382 382 410
rect 410 382 448 410
rect 476 382 514 410
rect 542 382 580 410
rect 608 382 646 410
rect 674 382 712 410
rect 740 382 778 410
rect 806 382 844 410
rect 872 382 910 410
rect 938 382 976 410
rect 1004 382 1042 410
rect 1070 382 1108 410
rect 1136 382 1174 410
rect 1202 382 1240 410
rect 1268 382 1306 410
rect 1334 382 1372 410
rect 1400 382 1438 410
rect 1466 382 1504 410
rect 1532 382 1570 410
rect 1598 382 1636 410
rect 1664 382 1702 410
rect 1730 382 1768 410
rect 1796 382 1834 410
rect 1862 382 1900 410
rect 1928 382 1966 410
rect 1994 382 2032 410
rect 2060 382 2098 410
rect 2126 382 2164 410
rect 2192 382 2230 410
rect 2258 382 2296 410
rect 2324 382 2362 410
rect 2390 382 2428 410
rect 2456 382 2494 410
rect 2522 382 2560 410
rect 2588 382 2626 410
rect 2654 382 2692 410
rect 2720 382 2758 410
rect 2786 382 2824 410
rect 2852 382 2890 410
rect 2918 382 2956 410
rect 2984 382 3022 410
rect 3050 382 3088 410
rect 3116 382 3154 410
rect 3182 382 3220 410
rect 3248 382 3286 410
rect 3314 382 3352 410
rect 3380 382 3418 410
rect 3446 382 3484 410
rect 3512 382 3550 410
rect 3578 382 3616 410
rect 3644 382 3682 410
rect 3710 382 3748 410
rect 3776 382 3814 410
rect 3842 382 3880 410
rect 3908 382 3946 410
rect 3974 382 4012 410
rect 4040 382 4078 410
rect 4106 382 4144 410
rect 4172 382 4210 410
rect 4238 382 4276 410
rect 4304 382 4342 410
rect 4370 382 4408 410
rect 4436 382 4474 410
rect 4502 382 4540 410
rect 4568 382 4573 410
rect -4573 344 4573 382
rect -4573 316 -4568 344
rect -4540 316 -4502 344
rect -4474 316 -4436 344
rect -4408 316 -4370 344
rect -4342 316 -4304 344
rect -4276 316 -4238 344
rect -4210 316 -4172 344
rect -4144 316 -4106 344
rect -4078 316 -4040 344
rect -4012 316 -3974 344
rect -3946 316 -3908 344
rect -3880 316 -3842 344
rect -3814 316 -3776 344
rect -3748 316 -3710 344
rect -3682 316 -3644 344
rect -3616 316 -3578 344
rect -3550 316 -3512 344
rect -3484 316 -3446 344
rect -3418 316 -3380 344
rect -3352 316 -3314 344
rect -3286 316 -3248 344
rect -3220 316 -3182 344
rect -3154 316 -3116 344
rect -3088 316 -3050 344
rect -3022 316 -2984 344
rect -2956 316 -2918 344
rect -2890 316 -2852 344
rect -2824 316 -2786 344
rect -2758 316 -2720 344
rect -2692 316 -2654 344
rect -2626 316 -2588 344
rect -2560 316 -2522 344
rect -2494 316 -2456 344
rect -2428 316 -2390 344
rect -2362 316 -2324 344
rect -2296 316 -2258 344
rect -2230 316 -2192 344
rect -2164 316 -2126 344
rect -2098 316 -2060 344
rect -2032 316 -1994 344
rect -1966 316 -1928 344
rect -1900 316 -1862 344
rect -1834 316 -1796 344
rect -1768 316 -1730 344
rect -1702 316 -1664 344
rect -1636 316 -1598 344
rect -1570 316 -1532 344
rect -1504 316 -1466 344
rect -1438 316 -1400 344
rect -1372 316 -1334 344
rect -1306 316 -1268 344
rect -1240 316 -1202 344
rect -1174 316 -1136 344
rect -1108 316 -1070 344
rect -1042 316 -1004 344
rect -976 316 -938 344
rect -910 316 -872 344
rect -844 316 -806 344
rect -778 316 -740 344
rect -712 316 -674 344
rect -646 316 -608 344
rect -580 316 -542 344
rect -514 316 -476 344
rect -448 316 -410 344
rect -382 316 -344 344
rect -316 316 -278 344
rect -250 316 -212 344
rect -184 316 -146 344
rect -118 316 -80 344
rect -52 316 -14 344
rect 14 316 52 344
rect 80 316 118 344
rect 146 316 184 344
rect 212 316 250 344
rect 278 316 316 344
rect 344 316 382 344
rect 410 316 448 344
rect 476 316 514 344
rect 542 316 580 344
rect 608 316 646 344
rect 674 316 712 344
rect 740 316 778 344
rect 806 316 844 344
rect 872 316 910 344
rect 938 316 976 344
rect 1004 316 1042 344
rect 1070 316 1108 344
rect 1136 316 1174 344
rect 1202 316 1240 344
rect 1268 316 1306 344
rect 1334 316 1372 344
rect 1400 316 1438 344
rect 1466 316 1504 344
rect 1532 316 1570 344
rect 1598 316 1636 344
rect 1664 316 1702 344
rect 1730 316 1768 344
rect 1796 316 1834 344
rect 1862 316 1900 344
rect 1928 316 1966 344
rect 1994 316 2032 344
rect 2060 316 2098 344
rect 2126 316 2164 344
rect 2192 316 2230 344
rect 2258 316 2296 344
rect 2324 316 2362 344
rect 2390 316 2428 344
rect 2456 316 2494 344
rect 2522 316 2560 344
rect 2588 316 2626 344
rect 2654 316 2692 344
rect 2720 316 2758 344
rect 2786 316 2824 344
rect 2852 316 2890 344
rect 2918 316 2956 344
rect 2984 316 3022 344
rect 3050 316 3088 344
rect 3116 316 3154 344
rect 3182 316 3220 344
rect 3248 316 3286 344
rect 3314 316 3352 344
rect 3380 316 3418 344
rect 3446 316 3484 344
rect 3512 316 3550 344
rect 3578 316 3616 344
rect 3644 316 3682 344
rect 3710 316 3748 344
rect 3776 316 3814 344
rect 3842 316 3880 344
rect 3908 316 3946 344
rect 3974 316 4012 344
rect 4040 316 4078 344
rect 4106 316 4144 344
rect 4172 316 4210 344
rect 4238 316 4276 344
rect 4304 316 4342 344
rect 4370 316 4408 344
rect 4436 316 4474 344
rect 4502 316 4540 344
rect 4568 316 4573 344
rect -4573 278 4573 316
rect -4573 250 -4568 278
rect -4540 250 -4502 278
rect -4474 250 -4436 278
rect -4408 250 -4370 278
rect -4342 250 -4304 278
rect -4276 250 -4238 278
rect -4210 250 -4172 278
rect -4144 250 -4106 278
rect -4078 250 -4040 278
rect -4012 250 -3974 278
rect -3946 250 -3908 278
rect -3880 250 -3842 278
rect -3814 250 -3776 278
rect -3748 250 -3710 278
rect -3682 250 -3644 278
rect -3616 250 -3578 278
rect -3550 250 -3512 278
rect -3484 250 -3446 278
rect -3418 250 -3380 278
rect -3352 250 -3314 278
rect -3286 250 -3248 278
rect -3220 250 -3182 278
rect -3154 250 -3116 278
rect -3088 250 -3050 278
rect -3022 250 -2984 278
rect -2956 250 -2918 278
rect -2890 250 -2852 278
rect -2824 250 -2786 278
rect -2758 250 -2720 278
rect -2692 250 -2654 278
rect -2626 250 -2588 278
rect -2560 250 -2522 278
rect -2494 250 -2456 278
rect -2428 250 -2390 278
rect -2362 250 -2324 278
rect -2296 250 -2258 278
rect -2230 250 -2192 278
rect -2164 250 -2126 278
rect -2098 250 -2060 278
rect -2032 250 -1994 278
rect -1966 250 -1928 278
rect -1900 250 -1862 278
rect -1834 250 -1796 278
rect -1768 250 -1730 278
rect -1702 250 -1664 278
rect -1636 250 -1598 278
rect -1570 250 -1532 278
rect -1504 250 -1466 278
rect -1438 250 -1400 278
rect -1372 250 -1334 278
rect -1306 250 -1268 278
rect -1240 250 -1202 278
rect -1174 250 -1136 278
rect -1108 250 -1070 278
rect -1042 250 -1004 278
rect -976 250 -938 278
rect -910 250 -872 278
rect -844 250 -806 278
rect -778 250 -740 278
rect -712 250 -674 278
rect -646 250 -608 278
rect -580 250 -542 278
rect -514 250 -476 278
rect -448 250 -410 278
rect -382 250 -344 278
rect -316 250 -278 278
rect -250 250 -212 278
rect -184 250 -146 278
rect -118 250 -80 278
rect -52 250 -14 278
rect 14 250 52 278
rect 80 250 118 278
rect 146 250 184 278
rect 212 250 250 278
rect 278 250 316 278
rect 344 250 382 278
rect 410 250 448 278
rect 476 250 514 278
rect 542 250 580 278
rect 608 250 646 278
rect 674 250 712 278
rect 740 250 778 278
rect 806 250 844 278
rect 872 250 910 278
rect 938 250 976 278
rect 1004 250 1042 278
rect 1070 250 1108 278
rect 1136 250 1174 278
rect 1202 250 1240 278
rect 1268 250 1306 278
rect 1334 250 1372 278
rect 1400 250 1438 278
rect 1466 250 1504 278
rect 1532 250 1570 278
rect 1598 250 1636 278
rect 1664 250 1702 278
rect 1730 250 1768 278
rect 1796 250 1834 278
rect 1862 250 1900 278
rect 1928 250 1966 278
rect 1994 250 2032 278
rect 2060 250 2098 278
rect 2126 250 2164 278
rect 2192 250 2230 278
rect 2258 250 2296 278
rect 2324 250 2362 278
rect 2390 250 2428 278
rect 2456 250 2494 278
rect 2522 250 2560 278
rect 2588 250 2626 278
rect 2654 250 2692 278
rect 2720 250 2758 278
rect 2786 250 2824 278
rect 2852 250 2890 278
rect 2918 250 2956 278
rect 2984 250 3022 278
rect 3050 250 3088 278
rect 3116 250 3154 278
rect 3182 250 3220 278
rect 3248 250 3286 278
rect 3314 250 3352 278
rect 3380 250 3418 278
rect 3446 250 3484 278
rect 3512 250 3550 278
rect 3578 250 3616 278
rect 3644 250 3682 278
rect 3710 250 3748 278
rect 3776 250 3814 278
rect 3842 250 3880 278
rect 3908 250 3946 278
rect 3974 250 4012 278
rect 4040 250 4078 278
rect 4106 250 4144 278
rect 4172 250 4210 278
rect 4238 250 4276 278
rect 4304 250 4342 278
rect 4370 250 4408 278
rect 4436 250 4474 278
rect 4502 250 4540 278
rect 4568 250 4573 278
rect -4573 212 4573 250
rect -4573 184 -4568 212
rect -4540 184 -4502 212
rect -4474 184 -4436 212
rect -4408 184 -4370 212
rect -4342 184 -4304 212
rect -4276 184 -4238 212
rect -4210 184 -4172 212
rect -4144 184 -4106 212
rect -4078 184 -4040 212
rect -4012 184 -3974 212
rect -3946 184 -3908 212
rect -3880 184 -3842 212
rect -3814 184 -3776 212
rect -3748 184 -3710 212
rect -3682 184 -3644 212
rect -3616 184 -3578 212
rect -3550 184 -3512 212
rect -3484 184 -3446 212
rect -3418 184 -3380 212
rect -3352 184 -3314 212
rect -3286 184 -3248 212
rect -3220 184 -3182 212
rect -3154 184 -3116 212
rect -3088 184 -3050 212
rect -3022 184 -2984 212
rect -2956 184 -2918 212
rect -2890 184 -2852 212
rect -2824 184 -2786 212
rect -2758 184 -2720 212
rect -2692 184 -2654 212
rect -2626 184 -2588 212
rect -2560 184 -2522 212
rect -2494 184 -2456 212
rect -2428 184 -2390 212
rect -2362 184 -2324 212
rect -2296 184 -2258 212
rect -2230 184 -2192 212
rect -2164 184 -2126 212
rect -2098 184 -2060 212
rect -2032 184 -1994 212
rect -1966 184 -1928 212
rect -1900 184 -1862 212
rect -1834 184 -1796 212
rect -1768 184 -1730 212
rect -1702 184 -1664 212
rect -1636 184 -1598 212
rect -1570 184 -1532 212
rect -1504 184 -1466 212
rect -1438 184 -1400 212
rect -1372 184 -1334 212
rect -1306 184 -1268 212
rect -1240 184 -1202 212
rect -1174 184 -1136 212
rect -1108 184 -1070 212
rect -1042 184 -1004 212
rect -976 184 -938 212
rect -910 184 -872 212
rect -844 184 -806 212
rect -778 184 -740 212
rect -712 184 -674 212
rect -646 184 -608 212
rect -580 184 -542 212
rect -514 184 -476 212
rect -448 184 -410 212
rect -382 184 -344 212
rect -316 184 -278 212
rect -250 184 -212 212
rect -184 184 -146 212
rect -118 184 -80 212
rect -52 184 -14 212
rect 14 184 52 212
rect 80 184 118 212
rect 146 184 184 212
rect 212 184 250 212
rect 278 184 316 212
rect 344 184 382 212
rect 410 184 448 212
rect 476 184 514 212
rect 542 184 580 212
rect 608 184 646 212
rect 674 184 712 212
rect 740 184 778 212
rect 806 184 844 212
rect 872 184 910 212
rect 938 184 976 212
rect 1004 184 1042 212
rect 1070 184 1108 212
rect 1136 184 1174 212
rect 1202 184 1240 212
rect 1268 184 1306 212
rect 1334 184 1372 212
rect 1400 184 1438 212
rect 1466 184 1504 212
rect 1532 184 1570 212
rect 1598 184 1636 212
rect 1664 184 1702 212
rect 1730 184 1768 212
rect 1796 184 1834 212
rect 1862 184 1900 212
rect 1928 184 1966 212
rect 1994 184 2032 212
rect 2060 184 2098 212
rect 2126 184 2164 212
rect 2192 184 2230 212
rect 2258 184 2296 212
rect 2324 184 2362 212
rect 2390 184 2428 212
rect 2456 184 2494 212
rect 2522 184 2560 212
rect 2588 184 2626 212
rect 2654 184 2692 212
rect 2720 184 2758 212
rect 2786 184 2824 212
rect 2852 184 2890 212
rect 2918 184 2956 212
rect 2984 184 3022 212
rect 3050 184 3088 212
rect 3116 184 3154 212
rect 3182 184 3220 212
rect 3248 184 3286 212
rect 3314 184 3352 212
rect 3380 184 3418 212
rect 3446 184 3484 212
rect 3512 184 3550 212
rect 3578 184 3616 212
rect 3644 184 3682 212
rect 3710 184 3748 212
rect 3776 184 3814 212
rect 3842 184 3880 212
rect 3908 184 3946 212
rect 3974 184 4012 212
rect 4040 184 4078 212
rect 4106 184 4144 212
rect 4172 184 4210 212
rect 4238 184 4276 212
rect 4304 184 4342 212
rect 4370 184 4408 212
rect 4436 184 4474 212
rect 4502 184 4540 212
rect 4568 184 4573 212
rect -4573 146 4573 184
rect -4573 118 -4568 146
rect -4540 118 -4502 146
rect -4474 118 -4436 146
rect -4408 118 -4370 146
rect -4342 118 -4304 146
rect -4276 118 -4238 146
rect -4210 118 -4172 146
rect -4144 118 -4106 146
rect -4078 118 -4040 146
rect -4012 118 -3974 146
rect -3946 118 -3908 146
rect -3880 118 -3842 146
rect -3814 118 -3776 146
rect -3748 118 -3710 146
rect -3682 118 -3644 146
rect -3616 118 -3578 146
rect -3550 118 -3512 146
rect -3484 118 -3446 146
rect -3418 118 -3380 146
rect -3352 118 -3314 146
rect -3286 118 -3248 146
rect -3220 118 -3182 146
rect -3154 118 -3116 146
rect -3088 118 -3050 146
rect -3022 118 -2984 146
rect -2956 118 -2918 146
rect -2890 118 -2852 146
rect -2824 118 -2786 146
rect -2758 118 -2720 146
rect -2692 118 -2654 146
rect -2626 118 -2588 146
rect -2560 118 -2522 146
rect -2494 118 -2456 146
rect -2428 118 -2390 146
rect -2362 118 -2324 146
rect -2296 118 -2258 146
rect -2230 118 -2192 146
rect -2164 118 -2126 146
rect -2098 118 -2060 146
rect -2032 118 -1994 146
rect -1966 118 -1928 146
rect -1900 118 -1862 146
rect -1834 118 -1796 146
rect -1768 118 -1730 146
rect -1702 118 -1664 146
rect -1636 118 -1598 146
rect -1570 118 -1532 146
rect -1504 118 -1466 146
rect -1438 118 -1400 146
rect -1372 118 -1334 146
rect -1306 118 -1268 146
rect -1240 118 -1202 146
rect -1174 118 -1136 146
rect -1108 118 -1070 146
rect -1042 118 -1004 146
rect -976 118 -938 146
rect -910 118 -872 146
rect -844 118 -806 146
rect -778 118 -740 146
rect -712 118 -674 146
rect -646 118 -608 146
rect -580 118 -542 146
rect -514 118 -476 146
rect -448 118 -410 146
rect -382 118 -344 146
rect -316 118 -278 146
rect -250 118 -212 146
rect -184 118 -146 146
rect -118 118 -80 146
rect -52 118 -14 146
rect 14 118 52 146
rect 80 118 118 146
rect 146 118 184 146
rect 212 118 250 146
rect 278 118 316 146
rect 344 118 382 146
rect 410 118 448 146
rect 476 118 514 146
rect 542 118 580 146
rect 608 118 646 146
rect 674 118 712 146
rect 740 118 778 146
rect 806 118 844 146
rect 872 118 910 146
rect 938 118 976 146
rect 1004 118 1042 146
rect 1070 118 1108 146
rect 1136 118 1174 146
rect 1202 118 1240 146
rect 1268 118 1306 146
rect 1334 118 1372 146
rect 1400 118 1438 146
rect 1466 118 1504 146
rect 1532 118 1570 146
rect 1598 118 1636 146
rect 1664 118 1702 146
rect 1730 118 1768 146
rect 1796 118 1834 146
rect 1862 118 1900 146
rect 1928 118 1966 146
rect 1994 118 2032 146
rect 2060 118 2098 146
rect 2126 118 2164 146
rect 2192 118 2230 146
rect 2258 118 2296 146
rect 2324 118 2362 146
rect 2390 118 2428 146
rect 2456 118 2494 146
rect 2522 118 2560 146
rect 2588 118 2626 146
rect 2654 118 2692 146
rect 2720 118 2758 146
rect 2786 118 2824 146
rect 2852 118 2890 146
rect 2918 118 2956 146
rect 2984 118 3022 146
rect 3050 118 3088 146
rect 3116 118 3154 146
rect 3182 118 3220 146
rect 3248 118 3286 146
rect 3314 118 3352 146
rect 3380 118 3418 146
rect 3446 118 3484 146
rect 3512 118 3550 146
rect 3578 118 3616 146
rect 3644 118 3682 146
rect 3710 118 3748 146
rect 3776 118 3814 146
rect 3842 118 3880 146
rect 3908 118 3946 146
rect 3974 118 4012 146
rect 4040 118 4078 146
rect 4106 118 4144 146
rect 4172 118 4210 146
rect 4238 118 4276 146
rect 4304 118 4342 146
rect 4370 118 4408 146
rect 4436 118 4474 146
rect 4502 118 4540 146
rect 4568 118 4573 146
rect -4573 80 4573 118
rect -4573 52 -4568 80
rect -4540 52 -4502 80
rect -4474 52 -4436 80
rect -4408 52 -4370 80
rect -4342 52 -4304 80
rect -4276 52 -4238 80
rect -4210 52 -4172 80
rect -4144 52 -4106 80
rect -4078 52 -4040 80
rect -4012 52 -3974 80
rect -3946 52 -3908 80
rect -3880 52 -3842 80
rect -3814 52 -3776 80
rect -3748 52 -3710 80
rect -3682 52 -3644 80
rect -3616 52 -3578 80
rect -3550 52 -3512 80
rect -3484 52 -3446 80
rect -3418 52 -3380 80
rect -3352 52 -3314 80
rect -3286 52 -3248 80
rect -3220 52 -3182 80
rect -3154 52 -3116 80
rect -3088 52 -3050 80
rect -3022 52 -2984 80
rect -2956 52 -2918 80
rect -2890 52 -2852 80
rect -2824 52 -2786 80
rect -2758 52 -2720 80
rect -2692 52 -2654 80
rect -2626 52 -2588 80
rect -2560 52 -2522 80
rect -2494 52 -2456 80
rect -2428 52 -2390 80
rect -2362 52 -2324 80
rect -2296 52 -2258 80
rect -2230 52 -2192 80
rect -2164 52 -2126 80
rect -2098 52 -2060 80
rect -2032 52 -1994 80
rect -1966 52 -1928 80
rect -1900 52 -1862 80
rect -1834 52 -1796 80
rect -1768 52 -1730 80
rect -1702 52 -1664 80
rect -1636 52 -1598 80
rect -1570 52 -1532 80
rect -1504 52 -1466 80
rect -1438 52 -1400 80
rect -1372 52 -1334 80
rect -1306 52 -1268 80
rect -1240 52 -1202 80
rect -1174 52 -1136 80
rect -1108 52 -1070 80
rect -1042 52 -1004 80
rect -976 52 -938 80
rect -910 52 -872 80
rect -844 52 -806 80
rect -778 52 -740 80
rect -712 52 -674 80
rect -646 52 -608 80
rect -580 52 -542 80
rect -514 52 -476 80
rect -448 52 -410 80
rect -382 52 -344 80
rect -316 52 -278 80
rect -250 52 -212 80
rect -184 52 -146 80
rect -118 52 -80 80
rect -52 52 -14 80
rect 14 52 52 80
rect 80 52 118 80
rect 146 52 184 80
rect 212 52 250 80
rect 278 52 316 80
rect 344 52 382 80
rect 410 52 448 80
rect 476 52 514 80
rect 542 52 580 80
rect 608 52 646 80
rect 674 52 712 80
rect 740 52 778 80
rect 806 52 844 80
rect 872 52 910 80
rect 938 52 976 80
rect 1004 52 1042 80
rect 1070 52 1108 80
rect 1136 52 1174 80
rect 1202 52 1240 80
rect 1268 52 1306 80
rect 1334 52 1372 80
rect 1400 52 1438 80
rect 1466 52 1504 80
rect 1532 52 1570 80
rect 1598 52 1636 80
rect 1664 52 1702 80
rect 1730 52 1768 80
rect 1796 52 1834 80
rect 1862 52 1900 80
rect 1928 52 1966 80
rect 1994 52 2032 80
rect 2060 52 2098 80
rect 2126 52 2164 80
rect 2192 52 2230 80
rect 2258 52 2296 80
rect 2324 52 2362 80
rect 2390 52 2428 80
rect 2456 52 2494 80
rect 2522 52 2560 80
rect 2588 52 2626 80
rect 2654 52 2692 80
rect 2720 52 2758 80
rect 2786 52 2824 80
rect 2852 52 2890 80
rect 2918 52 2956 80
rect 2984 52 3022 80
rect 3050 52 3088 80
rect 3116 52 3154 80
rect 3182 52 3220 80
rect 3248 52 3286 80
rect 3314 52 3352 80
rect 3380 52 3418 80
rect 3446 52 3484 80
rect 3512 52 3550 80
rect 3578 52 3616 80
rect 3644 52 3682 80
rect 3710 52 3748 80
rect 3776 52 3814 80
rect 3842 52 3880 80
rect 3908 52 3946 80
rect 3974 52 4012 80
rect 4040 52 4078 80
rect 4106 52 4144 80
rect 4172 52 4210 80
rect 4238 52 4276 80
rect 4304 52 4342 80
rect 4370 52 4408 80
rect 4436 52 4474 80
rect 4502 52 4540 80
rect 4568 52 4573 80
rect -4573 14 4573 52
rect -4573 -14 -4568 14
rect -4540 -14 -4502 14
rect -4474 -14 -4436 14
rect -4408 -14 -4370 14
rect -4342 -14 -4304 14
rect -4276 -14 -4238 14
rect -4210 -14 -4172 14
rect -4144 -14 -4106 14
rect -4078 -14 -4040 14
rect -4012 -14 -3974 14
rect -3946 -14 -3908 14
rect -3880 -14 -3842 14
rect -3814 -14 -3776 14
rect -3748 -14 -3710 14
rect -3682 -14 -3644 14
rect -3616 -14 -3578 14
rect -3550 -14 -3512 14
rect -3484 -14 -3446 14
rect -3418 -14 -3380 14
rect -3352 -14 -3314 14
rect -3286 -14 -3248 14
rect -3220 -14 -3182 14
rect -3154 -14 -3116 14
rect -3088 -14 -3050 14
rect -3022 -14 -2984 14
rect -2956 -14 -2918 14
rect -2890 -14 -2852 14
rect -2824 -14 -2786 14
rect -2758 -14 -2720 14
rect -2692 -14 -2654 14
rect -2626 -14 -2588 14
rect -2560 -14 -2522 14
rect -2494 -14 -2456 14
rect -2428 -14 -2390 14
rect -2362 -14 -2324 14
rect -2296 -14 -2258 14
rect -2230 -14 -2192 14
rect -2164 -14 -2126 14
rect -2098 -14 -2060 14
rect -2032 -14 -1994 14
rect -1966 -14 -1928 14
rect -1900 -14 -1862 14
rect -1834 -14 -1796 14
rect -1768 -14 -1730 14
rect -1702 -14 -1664 14
rect -1636 -14 -1598 14
rect -1570 -14 -1532 14
rect -1504 -14 -1466 14
rect -1438 -14 -1400 14
rect -1372 -14 -1334 14
rect -1306 -14 -1268 14
rect -1240 -14 -1202 14
rect -1174 -14 -1136 14
rect -1108 -14 -1070 14
rect -1042 -14 -1004 14
rect -976 -14 -938 14
rect -910 -14 -872 14
rect -844 -14 -806 14
rect -778 -14 -740 14
rect -712 -14 -674 14
rect -646 -14 -608 14
rect -580 -14 -542 14
rect -514 -14 -476 14
rect -448 -14 -410 14
rect -382 -14 -344 14
rect -316 -14 -278 14
rect -250 -14 -212 14
rect -184 -14 -146 14
rect -118 -14 -80 14
rect -52 -14 -14 14
rect 14 -14 52 14
rect 80 -14 118 14
rect 146 -14 184 14
rect 212 -14 250 14
rect 278 -14 316 14
rect 344 -14 382 14
rect 410 -14 448 14
rect 476 -14 514 14
rect 542 -14 580 14
rect 608 -14 646 14
rect 674 -14 712 14
rect 740 -14 778 14
rect 806 -14 844 14
rect 872 -14 910 14
rect 938 -14 976 14
rect 1004 -14 1042 14
rect 1070 -14 1108 14
rect 1136 -14 1174 14
rect 1202 -14 1240 14
rect 1268 -14 1306 14
rect 1334 -14 1372 14
rect 1400 -14 1438 14
rect 1466 -14 1504 14
rect 1532 -14 1570 14
rect 1598 -14 1636 14
rect 1664 -14 1702 14
rect 1730 -14 1768 14
rect 1796 -14 1834 14
rect 1862 -14 1900 14
rect 1928 -14 1966 14
rect 1994 -14 2032 14
rect 2060 -14 2098 14
rect 2126 -14 2164 14
rect 2192 -14 2230 14
rect 2258 -14 2296 14
rect 2324 -14 2362 14
rect 2390 -14 2428 14
rect 2456 -14 2494 14
rect 2522 -14 2560 14
rect 2588 -14 2626 14
rect 2654 -14 2692 14
rect 2720 -14 2758 14
rect 2786 -14 2824 14
rect 2852 -14 2890 14
rect 2918 -14 2956 14
rect 2984 -14 3022 14
rect 3050 -14 3088 14
rect 3116 -14 3154 14
rect 3182 -14 3220 14
rect 3248 -14 3286 14
rect 3314 -14 3352 14
rect 3380 -14 3418 14
rect 3446 -14 3484 14
rect 3512 -14 3550 14
rect 3578 -14 3616 14
rect 3644 -14 3682 14
rect 3710 -14 3748 14
rect 3776 -14 3814 14
rect 3842 -14 3880 14
rect 3908 -14 3946 14
rect 3974 -14 4012 14
rect 4040 -14 4078 14
rect 4106 -14 4144 14
rect 4172 -14 4210 14
rect 4238 -14 4276 14
rect 4304 -14 4342 14
rect 4370 -14 4408 14
rect 4436 -14 4474 14
rect 4502 -14 4540 14
rect 4568 -14 4573 14
rect -4573 -52 4573 -14
rect -4573 -80 -4568 -52
rect -4540 -80 -4502 -52
rect -4474 -80 -4436 -52
rect -4408 -80 -4370 -52
rect -4342 -80 -4304 -52
rect -4276 -80 -4238 -52
rect -4210 -80 -4172 -52
rect -4144 -80 -4106 -52
rect -4078 -80 -4040 -52
rect -4012 -80 -3974 -52
rect -3946 -80 -3908 -52
rect -3880 -80 -3842 -52
rect -3814 -80 -3776 -52
rect -3748 -80 -3710 -52
rect -3682 -80 -3644 -52
rect -3616 -80 -3578 -52
rect -3550 -80 -3512 -52
rect -3484 -80 -3446 -52
rect -3418 -80 -3380 -52
rect -3352 -80 -3314 -52
rect -3286 -80 -3248 -52
rect -3220 -80 -3182 -52
rect -3154 -80 -3116 -52
rect -3088 -80 -3050 -52
rect -3022 -80 -2984 -52
rect -2956 -80 -2918 -52
rect -2890 -80 -2852 -52
rect -2824 -80 -2786 -52
rect -2758 -80 -2720 -52
rect -2692 -80 -2654 -52
rect -2626 -80 -2588 -52
rect -2560 -80 -2522 -52
rect -2494 -80 -2456 -52
rect -2428 -80 -2390 -52
rect -2362 -80 -2324 -52
rect -2296 -80 -2258 -52
rect -2230 -80 -2192 -52
rect -2164 -80 -2126 -52
rect -2098 -80 -2060 -52
rect -2032 -80 -1994 -52
rect -1966 -80 -1928 -52
rect -1900 -80 -1862 -52
rect -1834 -80 -1796 -52
rect -1768 -80 -1730 -52
rect -1702 -80 -1664 -52
rect -1636 -80 -1598 -52
rect -1570 -80 -1532 -52
rect -1504 -80 -1466 -52
rect -1438 -80 -1400 -52
rect -1372 -80 -1334 -52
rect -1306 -80 -1268 -52
rect -1240 -80 -1202 -52
rect -1174 -80 -1136 -52
rect -1108 -80 -1070 -52
rect -1042 -80 -1004 -52
rect -976 -80 -938 -52
rect -910 -80 -872 -52
rect -844 -80 -806 -52
rect -778 -80 -740 -52
rect -712 -80 -674 -52
rect -646 -80 -608 -52
rect -580 -80 -542 -52
rect -514 -80 -476 -52
rect -448 -80 -410 -52
rect -382 -80 -344 -52
rect -316 -80 -278 -52
rect -250 -80 -212 -52
rect -184 -80 -146 -52
rect -118 -80 -80 -52
rect -52 -80 -14 -52
rect 14 -80 52 -52
rect 80 -80 118 -52
rect 146 -80 184 -52
rect 212 -80 250 -52
rect 278 -80 316 -52
rect 344 -80 382 -52
rect 410 -80 448 -52
rect 476 -80 514 -52
rect 542 -80 580 -52
rect 608 -80 646 -52
rect 674 -80 712 -52
rect 740 -80 778 -52
rect 806 -80 844 -52
rect 872 -80 910 -52
rect 938 -80 976 -52
rect 1004 -80 1042 -52
rect 1070 -80 1108 -52
rect 1136 -80 1174 -52
rect 1202 -80 1240 -52
rect 1268 -80 1306 -52
rect 1334 -80 1372 -52
rect 1400 -80 1438 -52
rect 1466 -80 1504 -52
rect 1532 -80 1570 -52
rect 1598 -80 1636 -52
rect 1664 -80 1702 -52
rect 1730 -80 1768 -52
rect 1796 -80 1834 -52
rect 1862 -80 1900 -52
rect 1928 -80 1966 -52
rect 1994 -80 2032 -52
rect 2060 -80 2098 -52
rect 2126 -80 2164 -52
rect 2192 -80 2230 -52
rect 2258 -80 2296 -52
rect 2324 -80 2362 -52
rect 2390 -80 2428 -52
rect 2456 -80 2494 -52
rect 2522 -80 2560 -52
rect 2588 -80 2626 -52
rect 2654 -80 2692 -52
rect 2720 -80 2758 -52
rect 2786 -80 2824 -52
rect 2852 -80 2890 -52
rect 2918 -80 2956 -52
rect 2984 -80 3022 -52
rect 3050 -80 3088 -52
rect 3116 -80 3154 -52
rect 3182 -80 3220 -52
rect 3248 -80 3286 -52
rect 3314 -80 3352 -52
rect 3380 -80 3418 -52
rect 3446 -80 3484 -52
rect 3512 -80 3550 -52
rect 3578 -80 3616 -52
rect 3644 -80 3682 -52
rect 3710 -80 3748 -52
rect 3776 -80 3814 -52
rect 3842 -80 3880 -52
rect 3908 -80 3946 -52
rect 3974 -80 4012 -52
rect 4040 -80 4078 -52
rect 4106 -80 4144 -52
rect 4172 -80 4210 -52
rect 4238 -80 4276 -52
rect 4304 -80 4342 -52
rect 4370 -80 4408 -52
rect 4436 -80 4474 -52
rect 4502 -80 4540 -52
rect 4568 -80 4573 -52
rect -4573 -118 4573 -80
rect -4573 -146 -4568 -118
rect -4540 -146 -4502 -118
rect -4474 -146 -4436 -118
rect -4408 -146 -4370 -118
rect -4342 -146 -4304 -118
rect -4276 -146 -4238 -118
rect -4210 -146 -4172 -118
rect -4144 -146 -4106 -118
rect -4078 -146 -4040 -118
rect -4012 -146 -3974 -118
rect -3946 -146 -3908 -118
rect -3880 -146 -3842 -118
rect -3814 -146 -3776 -118
rect -3748 -146 -3710 -118
rect -3682 -146 -3644 -118
rect -3616 -146 -3578 -118
rect -3550 -146 -3512 -118
rect -3484 -146 -3446 -118
rect -3418 -146 -3380 -118
rect -3352 -146 -3314 -118
rect -3286 -146 -3248 -118
rect -3220 -146 -3182 -118
rect -3154 -146 -3116 -118
rect -3088 -146 -3050 -118
rect -3022 -146 -2984 -118
rect -2956 -146 -2918 -118
rect -2890 -146 -2852 -118
rect -2824 -146 -2786 -118
rect -2758 -146 -2720 -118
rect -2692 -146 -2654 -118
rect -2626 -146 -2588 -118
rect -2560 -146 -2522 -118
rect -2494 -146 -2456 -118
rect -2428 -146 -2390 -118
rect -2362 -146 -2324 -118
rect -2296 -146 -2258 -118
rect -2230 -146 -2192 -118
rect -2164 -146 -2126 -118
rect -2098 -146 -2060 -118
rect -2032 -146 -1994 -118
rect -1966 -146 -1928 -118
rect -1900 -146 -1862 -118
rect -1834 -146 -1796 -118
rect -1768 -146 -1730 -118
rect -1702 -146 -1664 -118
rect -1636 -146 -1598 -118
rect -1570 -146 -1532 -118
rect -1504 -146 -1466 -118
rect -1438 -146 -1400 -118
rect -1372 -146 -1334 -118
rect -1306 -146 -1268 -118
rect -1240 -146 -1202 -118
rect -1174 -146 -1136 -118
rect -1108 -146 -1070 -118
rect -1042 -146 -1004 -118
rect -976 -146 -938 -118
rect -910 -146 -872 -118
rect -844 -146 -806 -118
rect -778 -146 -740 -118
rect -712 -146 -674 -118
rect -646 -146 -608 -118
rect -580 -146 -542 -118
rect -514 -146 -476 -118
rect -448 -146 -410 -118
rect -382 -146 -344 -118
rect -316 -146 -278 -118
rect -250 -146 -212 -118
rect -184 -146 -146 -118
rect -118 -146 -80 -118
rect -52 -146 -14 -118
rect 14 -146 52 -118
rect 80 -146 118 -118
rect 146 -146 184 -118
rect 212 -146 250 -118
rect 278 -146 316 -118
rect 344 -146 382 -118
rect 410 -146 448 -118
rect 476 -146 514 -118
rect 542 -146 580 -118
rect 608 -146 646 -118
rect 674 -146 712 -118
rect 740 -146 778 -118
rect 806 -146 844 -118
rect 872 -146 910 -118
rect 938 -146 976 -118
rect 1004 -146 1042 -118
rect 1070 -146 1108 -118
rect 1136 -146 1174 -118
rect 1202 -146 1240 -118
rect 1268 -146 1306 -118
rect 1334 -146 1372 -118
rect 1400 -146 1438 -118
rect 1466 -146 1504 -118
rect 1532 -146 1570 -118
rect 1598 -146 1636 -118
rect 1664 -146 1702 -118
rect 1730 -146 1768 -118
rect 1796 -146 1834 -118
rect 1862 -146 1900 -118
rect 1928 -146 1966 -118
rect 1994 -146 2032 -118
rect 2060 -146 2098 -118
rect 2126 -146 2164 -118
rect 2192 -146 2230 -118
rect 2258 -146 2296 -118
rect 2324 -146 2362 -118
rect 2390 -146 2428 -118
rect 2456 -146 2494 -118
rect 2522 -146 2560 -118
rect 2588 -146 2626 -118
rect 2654 -146 2692 -118
rect 2720 -146 2758 -118
rect 2786 -146 2824 -118
rect 2852 -146 2890 -118
rect 2918 -146 2956 -118
rect 2984 -146 3022 -118
rect 3050 -146 3088 -118
rect 3116 -146 3154 -118
rect 3182 -146 3220 -118
rect 3248 -146 3286 -118
rect 3314 -146 3352 -118
rect 3380 -146 3418 -118
rect 3446 -146 3484 -118
rect 3512 -146 3550 -118
rect 3578 -146 3616 -118
rect 3644 -146 3682 -118
rect 3710 -146 3748 -118
rect 3776 -146 3814 -118
rect 3842 -146 3880 -118
rect 3908 -146 3946 -118
rect 3974 -146 4012 -118
rect 4040 -146 4078 -118
rect 4106 -146 4144 -118
rect 4172 -146 4210 -118
rect 4238 -146 4276 -118
rect 4304 -146 4342 -118
rect 4370 -146 4408 -118
rect 4436 -146 4474 -118
rect 4502 -146 4540 -118
rect 4568 -146 4573 -118
rect -4573 -184 4573 -146
rect -4573 -212 -4568 -184
rect -4540 -212 -4502 -184
rect -4474 -212 -4436 -184
rect -4408 -212 -4370 -184
rect -4342 -212 -4304 -184
rect -4276 -212 -4238 -184
rect -4210 -212 -4172 -184
rect -4144 -212 -4106 -184
rect -4078 -212 -4040 -184
rect -4012 -212 -3974 -184
rect -3946 -212 -3908 -184
rect -3880 -212 -3842 -184
rect -3814 -212 -3776 -184
rect -3748 -212 -3710 -184
rect -3682 -212 -3644 -184
rect -3616 -212 -3578 -184
rect -3550 -212 -3512 -184
rect -3484 -212 -3446 -184
rect -3418 -212 -3380 -184
rect -3352 -212 -3314 -184
rect -3286 -212 -3248 -184
rect -3220 -212 -3182 -184
rect -3154 -212 -3116 -184
rect -3088 -212 -3050 -184
rect -3022 -212 -2984 -184
rect -2956 -212 -2918 -184
rect -2890 -212 -2852 -184
rect -2824 -212 -2786 -184
rect -2758 -212 -2720 -184
rect -2692 -212 -2654 -184
rect -2626 -212 -2588 -184
rect -2560 -212 -2522 -184
rect -2494 -212 -2456 -184
rect -2428 -212 -2390 -184
rect -2362 -212 -2324 -184
rect -2296 -212 -2258 -184
rect -2230 -212 -2192 -184
rect -2164 -212 -2126 -184
rect -2098 -212 -2060 -184
rect -2032 -212 -1994 -184
rect -1966 -212 -1928 -184
rect -1900 -212 -1862 -184
rect -1834 -212 -1796 -184
rect -1768 -212 -1730 -184
rect -1702 -212 -1664 -184
rect -1636 -212 -1598 -184
rect -1570 -212 -1532 -184
rect -1504 -212 -1466 -184
rect -1438 -212 -1400 -184
rect -1372 -212 -1334 -184
rect -1306 -212 -1268 -184
rect -1240 -212 -1202 -184
rect -1174 -212 -1136 -184
rect -1108 -212 -1070 -184
rect -1042 -212 -1004 -184
rect -976 -212 -938 -184
rect -910 -212 -872 -184
rect -844 -212 -806 -184
rect -778 -212 -740 -184
rect -712 -212 -674 -184
rect -646 -212 -608 -184
rect -580 -212 -542 -184
rect -514 -212 -476 -184
rect -448 -212 -410 -184
rect -382 -212 -344 -184
rect -316 -212 -278 -184
rect -250 -212 -212 -184
rect -184 -212 -146 -184
rect -118 -212 -80 -184
rect -52 -212 -14 -184
rect 14 -212 52 -184
rect 80 -212 118 -184
rect 146 -212 184 -184
rect 212 -212 250 -184
rect 278 -212 316 -184
rect 344 -212 382 -184
rect 410 -212 448 -184
rect 476 -212 514 -184
rect 542 -212 580 -184
rect 608 -212 646 -184
rect 674 -212 712 -184
rect 740 -212 778 -184
rect 806 -212 844 -184
rect 872 -212 910 -184
rect 938 -212 976 -184
rect 1004 -212 1042 -184
rect 1070 -212 1108 -184
rect 1136 -212 1174 -184
rect 1202 -212 1240 -184
rect 1268 -212 1306 -184
rect 1334 -212 1372 -184
rect 1400 -212 1438 -184
rect 1466 -212 1504 -184
rect 1532 -212 1570 -184
rect 1598 -212 1636 -184
rect 1664 -212 1702 -184
rect 1730 -212 1768 -184
rect 1796 -212 1834 -184
rect 1862 -212 1900 -184
rect 1928 -212 1966 -184
rect 1994 -212 2032 -184
rect 2060 -212 2098 -184
rect 2126 -212 2164 -184
rect 2192 -212 2230 -184
rect 2258 -212 2296 -184
rect 2324 -212 2362 -184
rect 2390 -212 2428 -184
rect 2456 -212 2494 -184
rect 2522 -212 2560 -184
rect 2588 -212 2626 -184
rect 2654 -212 2692 -184
rect 2720 -212 2758 -184
rect 2786 -212 2824 -184
rect 2852 -212 2890 -184
rect 2918 -212 2956 -184
rect 2984 -212 3022 -184
rect 3050 -212 3088 -184
rect 3116 -212 3154 -184
rect 3182 -212 3220 -184
rect 3248 -212 3286 -184
rect 3314 -212 3352 -184
rect 3380 -212 3418 -184
rect 3446 -212 3484 -184
rect 3512 -212 3550 -184
rect 3578 -212 3616 -184
rect 3644 -212 3682 -184
rect 3710 -212 3748 -184
rect 3776 -212 3814 -184
rect 3842 -212 3880 -184
rect 3908 -212 3946 -184
rect 3974 -212 4012 -184
rect 4040 -212 4078 -184
rect 4106 -212 4144 -184
rect 4172 -212 4210 -184
rect 4238 -212 4276 -184
rect 4304 -212 4342 -184
rect 4370 -212 4408 -184
rect 4436 -212 4474 -184
rect 4502 -212 4540 -184
rect 4568 -212 4573 -184
rect -4573 -250 4573 -212
rect -4573 -278 -4568 -250
rect -4540 -278 -4502 -250
rect -4474 -278 -4436 -250
rect -4408 -278 -4370 -250
rect -4342 -278 -4304 -250
rect -4276 -278 -4238 -250
rect -4210 -278 -4172 -250
rect -4144 -278 -4106 -250
rect -4078 -278 -4040 -250
rect -4012 -278 -3974 -250
rect -3946 -278 -3908 -250
rect -3880 -278 -3842 -250
rect -3814 -278 -3776 -250
rect -3748 -278 -3710 -250
rect -3682 -278 -3644 -250
rect -3616 -278 -3578 -250
rect -3550 -278 -3512 -250
rect -3484 -278 -3446 -250
rect -3418 -278 -3380 -250
rect -3352 -278 -3314 -250
rect -3286 -278 -3248 -250
rect -3220 -278 -3182 -250
rect -3154 -278 -3116 -250
rect -3088 -278 -3050 -250
rect -3022 -278 -2984 -250
rect -2956 -278 -2918 -250
rect -2890 -278 -2852 -250
rect -2824 -278 -2786 -250
rect -2758 -278 -2720 -250
rect -2692 -278 -2654 -250
rect -2626 -278 -2588 -250
rect -2560 -278 -2522 -250
rect -2494 -278 -2456 -250
rect -2428 -278 -2390 -250
rect -2362 -278 -2324 -250
rect -2296 -278 -2258 -250
rect -2230 -278 -2192 -250
rect -2164 -278 -2126 -250
rect -2098 -278 -2060 -250
rect -2032 -278 -1994 -250
rect -1966 -278 -1928 -250
rect -1900 -278 -1862 -250
rect -1834 -278 -1796 -250
rect -1768 -278 -1730 -250
rect -1702 -278 -1664 -250
rect -1636 -278 -1598 -250
rect -1570 -278 -1532 -250
rect -1504 -278 -1466 -250
rect -1438 -278 -1400 -250
rect -1372 -278 -1334 -250
rect -1306 -278 -1268 -250
rect -1240 -278 -1202 -250
rect -1174 -278 -1136 -250
rect -1108 -278 -1070 -250
rect -1042 -278 -1004 -250
rect -976 -278 -938 -250
rect -910 -278 -872 -250
rect -844 -278 -806 -250
rect -778 -278 -740 -250
rect -712 -278 -674 -250
rect -646 -278 -608 -250
rect -580 -278 -542 -250
rect -514 -278 -476 -250
rect -448 -278 -410 -250
rect -382 -278 -344 -250
rect -316 -278 -278 -250
rect -250 -278 -212 -250
rect -184 -278 -146 -250
rect -118 -278 -80 -250
rect -52 -278 -14 -250
rect 14 -278 52 -250
rect 80 -278 118 -250
rect 146 -278 184 -250
rect 212 -278 250 -250
rect 278 -278 316 -250
rect 344 -278 382 -250
rect 410 -278 448 -250
rect 476 -278 514 -250
rect 542 -278 580 -250
rect 608 -278 646 -250
rect 674 -278 712 -250
rect 740 -278 778 -250
rect 806 -278 844 -250
rect 872 -278 910 -250
rect 938 -278 976 -250
rect 1004 -278 1042 -250
rect 1070 -278 1108 -250
rect 1136 -278 1174 -250
rect 1202 -278 1240 -250
rect 1268 -278 1306 -250
rect 1334 -278 1372 -250
rect 1400 -278 1438 -250
rect 1466 -278 1504 -250
rect 1532 -278 1570 -250
rect 1598 -278 1636 -250
rect 1664 -278 1702 -250
rect 1730 -278 1768 -250
rect 1796 -278 1834 -250
rect 1862 -278 1900 -250
rect 1928 -278 1966 -250
rect 1994 -278 2032 -250
rect 2060 -278 2098 -250
rect 2126 -278 2164 -250
rect 2192 -278 2230 -250
rect 2258 -278 2296 -250
rect 2324 -278 2362 -250
rect 2390 -278 2428 -250
rect 2456 -278 2494 -250
rect 2522 -278 2560 -250
rect 2588 -278 2626 -250
rect 2654 -278 2692 -250
rect 2720 -278 2758 -250
rect 2786 -278 2824 -250
rect 2852 -278 2890 -250
rect 2918 -278 2956 -250
rect 2984 -278 3022 -250
rect 3050 -278 3088 -250
rect 3116 -278 3154 -250
rect 3182 -278 3220 -250
rect 3248 -278 3286 -250
rect 3314 -278 3352 -250
rect 3380 -278 3418 -250
rect 3446 -278 3484 -250
rect 3512 -278 3550 -250
rect 3578 -278 3616 -250
rect 3644 -278 3682 -250
rect 3710 -278 3748 -250
rect 3776 -278 3814 -250
rect 3842 -278 3880 -250
rect 3908 -278 3946 -250
rect 3974 -278 4012 -250
rect 4040 -278 4078 -250
rect 4106 -278 4144 -250
rect 4172 -278 4210 -250
rect 4238 -278 4276 -250
rect 4304 -278 4342 -250
rect 4370 -278 4408 -250
rect 4436 -278 4474 -250
rect 4502 -278 4540 -250
rect 4568 -278 4573 -250
rect -4573 -316 4573 -278
rect -4573 -344 -4568 -316
rect -4540 -344 -4502 -316
rect -4474 -344 -4436 -316
rect -4408 -344 -4370 -316
rect -4342 -344 -4304 -316
rect -4276 -344 -4238 -316
rect -4210 -344 -4172 -316
rect -4144 -344 -4106 -316
rect -4078 -344 -4040 -316
rect -4012 -344 -3974 -316
rect -3946 -344 -3908 -316
rect -3880 -344 -3842 -316
rect -3814 -344 -3776 -316
rect -3748 -344 -3710 -316
rect -3682 -344 -3644 -316
rect -3616 -344 -3578 -316
rect -3550 -344 -3512 -316
rect -3484 -344 -3446 -316
rect -3418 -344 -3380 -316
rect -3352 -344 -3314 -316
rect -3286 -344 -3248 -316
rect -3220 -344 -3182 -316
rect -3154 -344 -3116 -316
rect -3088 -344 -3050 -316
rect -3022 -344 -2984 -316
rect -2956 -344 -2918 -316
rect -2890 -344 -2852 -316
rect -2824 -344 -2786 -316
rect -2758 -344 -2720 -316
rect -2692 -344 -2654 -316
rect -2626 -344 -2588 -316
rect -2560 -344 -2522 -316
rect -2494 -344 -2456 -316
rect -2428 -344 -2390 -316
rect -2362 -344 -2324 -316
rect -2296 -344 -2258 -316
rect -2230 -344 -2192 -316
rect -2164 -344 -2126 -316
rect -2098 -344 -2060 -316
rect -2032 -344 -1994 -316
rect -1966 -344 -1928 -316
rect -1900 -344 -1862 -316
rect -1834 -344 -1796 -316
rect -1768 -344 -1730 -316
rect -1702 -344 -1664 -316
rect -1636 -344 -1598 -316
rect -1570 -344 -1532 -316
rect -1504 -344 -1466 -316
rect -1438 -344 -1400 -316
rect -1372 -344 -1334 -316
rect -1306 -344 -1268 -316
rect -1240 -344 -1202 -316
rect -1174 -344 -1136 -316
rect -1108 -344 -1070 -316
rect -1042 -344 -1004 -316
rect -976 -344 -938 -316
rect -910 -344 -872 -316
rect -844 -344 -806 -316
rect -778 -344 -740 -316
rect -712 -344 -674 -316
rect -646 -344 -608 -316
rect -580 -344 -542 -316
rect -514 -344 -476 -316
rect -448 -344 -410 -316
rect -382 -344 -344 -316
rect -316 -344 -278 -316
rect -250 -344 -212 -316
rect -184 -344 -146 -316
rect -118 -344 -80 -316
rect -52 -344 -14 -316
rect 14 -344 52 -316
rect 80 -344 118 -316
rect 146 -344 184 -316
rect 212 -344 250 -316
rect 278 -344 316 -316
rect 344 -344 382 -316
rect 410 -344 448 -316
rect 476 -344 514 -316
rect 542 -344 580 -316
rect 608 -344 646 -316
rect 674 -344 712 -316
rect 740 -344 778 -316
rect 806 -344 844 -316
rect 872 -344 910 -316
rect 938 -344 976 -316
rect 1004 -344 1042 -316
rect 1070 -344 1108 -316
rect 1136 -344 1174 -316
rect 1202 -344 1240 -316
rect 1268 -344 1306 -316
rect 1334 -344 1372 -316
rect 1400 -344 1438 -316
rect 1466 -344 1504 -316
rect 1532 -344 1570 -316
rect 1598 -344 1636 -316
rect 1664 -344 1702 -316
rect 1730 -344 1768 -316
rect 1796 -344 1834 -316
rect 1862 -344 1900 -316
rect 1928 -344 1966 -316
rect 1994 -344 2032 -316
rect 2060 -344 2098 -316
rect 2126 -344 2164 -316
rect 2192 -344 2230 -316
rect 2258 -344 2296 -316
rect 2324 -344 2362 -316
rect 2390 -344 2428 -316
rect 2456 -344 2494 -316
rect 2522 -344 2560 -316
rect 2588 -344 2626 -316
rect 2654 -344 2692 -316
rect 2720 -344 2758 -316
rect 2786 -344 2824 -316
rect 2852 -344 2890 -316
rect 2918 -344 2956 -316
rect 2984 -344 3022 -316
rect 3050 -344 3088 -316
rect 3116 -344 3154 -316
rect 3182 -344 3220 -316
rect 3248 -344 3286 -316
rect 3314 -344 3352 -316
rect 3380 -344 3418 -316
rect 3446 -344 3484 -316
rect 3512 -344 3550 -316
rect 3578 -344 3616 -316
rect 3644 -344 3682 -316
rect 3710 -344 3748 -316
rect 3776 -344 3814 -316
rect 3842 -344 3880 -316
rect 3908 -344 3946 -316
rect 3974 -344 4012 -316
rect 4040 -344 4078 -316
rect 4106 -344 4144 -316
rect 4172 -344 4210 -316
rect 4238 -344 4276 -316
rect 4304 -344 4342 -316
rect 4370 -344 4408 -316
rect 4436 -344 4474 -316
rect 4502 -344 4540 -316
rect 4568 -344 4573 -316
rect -4573 -382 4573 -344
rect -4573 -410 -4568 -382
rect -4540 -410 -4502 -382
rect -4474 -410 -4436 -382
rect -4408 -410 -4370 -382
rect -4342 -410 -4304 -382
rect -4276 -410 -4238 -382
rect -4210 -410 -4172 -382
rect -4144 -410 -4106 -382
rect -4078 -410 -4040 -382
rect -4012 -410 -3974 -382
rect -3946 -410 -3908 -382
rect -3880 -410 -3842 -382
rect -3814 -410 -3776 -382
rect -3748 -410 -3710 -382
rect -3682 -410 -3644 -382
rect -3616 -410 -3578 -382
rect -3550 -410 -3512 -382
rect -3484 -410 -3446 -382
rect -3418 -410 -3380 -382
rect -3352 -410 -3314 -382
rect -3286 -410 -3248 -382
rect -3220 -410 -3182 -382
rect -3154 -410 -3116 -382
rect -3088 -410 -3050 -382
rect -3022 -410 -2984 -382
rect -2956 -410 -2918 -382
rect -2890 -410 -2852 -382
rect -2824 -410 -2786 -382
rect -2758 -410 -2720 -382
rect -2692 -410 -2654 -382
rect -2626 -410 -2588 -382
rect -2560 -410 -2522 -382
rect -2494 -410 -2456 -382
rect -2428 -410 -2390 -382
rect -2362 -410 -2324 -382
rect -2296 -410 -2258 -382
rect -2230 -410 -2192 -382
rect -2164 -410 -2126 -382
rect -2098 -410 -2060 -382
rect -2032 -410 -1994 -382
rect -1966 -410 -1928 -382
rect -1900 -410 -1862 -382
rect -1834 -410 -1796 -382
rect -1768 -410 -1730 -382
rect -1702 -410 -1664 -382
rect -1636 -410 -1598 -382
rect -1570 -410 -1532 -382
rect -1504 -410 -1466 -382
rect -1438 -410 -1400 -382
rect -1372 -410 -1334 -382
rect -1306 -410 -1268 -382
rect -1240 -410 -1202 -382
rect -1174 -410 -1136 -382
rect -1108 -410 -1070 -382
rect -1042 -410 -1004 -382
rect -976 -410 -938 -382
rect -910 -410 -872 -382
rect -844 -410 -806 -382
rect -778 -410 -740 -382
rect -712 -410 -674 -382
rect -646 -410 -608 -382
rect -580 -410 -542 -382
rect -514 -410 -476 -382
rect -448 -410 -410 -382
rect -382 -410 -344 -382
rect -316 -410 -278 -382
rect -250 -410 -212 -382
rect -184 -410 -146 -382
rect -118 -410 -80 -382
rect -52 -410 -14 -382
rect 14 -410 52 -382
rect 80 -410 118 -382
rect 146 -410 184 -382
rect 212 -410 250 -382
rect 278 -410 316 -382
rect 344 -410 382 -382
rect 410 -410 448 -382
rect 476 -410 514 -382
rect 542 -410 580 -382
rect 608 -410 646 -382
rect 674 -410 712 -382
rect 740 -410 778 -382
rect 806 -410 844 -382
rect 872 -410 910 -382
rect 938 -410 976 -382
rect 1004 -410 1042 -382
rect 1070 -410 1108 -382
rect 1136 -410 1174 -382
rect 1202 -410 1240 -382
rect 1268 -410 1306 -382
rect 1334 -410 1372 -382
rect 1400 -410 1438 -382
rect 1466 -410 1504 -382
rect 1532 -410 1570 -382
rect 1598 -410 1636 -382
rect 1664 -410 1702 -382
rect 1730 -410 1768 -382
rect 1796 -410 1834 -382
rect 1862 -410 1900 -382
rect 1928 -410 1966 -382
rect 1994 -410 2032 -382
rect 2060 -410 2098 -382
rect 2126 -410 2164 -382
rect 2192 -410 2230 -382
rect 2258 -410 2296 -382
rect 2324 -410 2362 -382
rect 2390 -410 2428 -382
rect 2456 -410 2494 -382
rect 2522 -410 2560 -382
rect 2588 -410 2626 -382
rect 2654 -410 2692 -382
rect 2720 -410 2758 -382
rect 2786 -410 2824 -382
rect 2852 -410 2890 -382
rect 2918 -410 2956 -382
rect 2984 -410 3022 -382
rect 3050 -410 3088 -382
rect 3116 -410 3154 -382
rect 3182 -410 3220 -382
rect 3248 -410 3286 -382
rect 3314 -410 3352 -382
rect 3380 -410 3418 -382
rect 3446 -410 3484 -382
rect 3512 -410 3550 -382
rect 3578 -410 3616 -382
rect 3644 -410 3682 -382
rect 3710 -410 3748 -382
rect 3776 -410 3814 -382
rect 3842 -410 3880 -382
rect 3908 -410 3946 -382
rect 3974 -410 4012 -382
rect 4040 -410 4078 -382
rect 4106 -410 4144 -382
rect 4172 -410 4210 -382
rect 4238 -410 4276 -382
rect 4304 -410 4342 -382
rect 4370 -410 4408 -382
rect 4436 -410 4474 -382
rect 4502 -410 4540 -382
rect 4568 -410 4573 -382
rect -4573 -448 4573 -410
rect -4573 -476 -4568 -448
rect -4540 -476 -4502 -448
rect -4474 -476 -4436 -448
rect -4408 -476 -4370 -448
rect -4342 -476 -4304 -448
rect -4276 -476 -4238 -448
rect -4210 -476 -4172 -448
rect -4144 -476 -4106 -448
rect -4078 -476 -4040 -448
rect -4012 -476 -3974 -448
rect -3946 -476 -3908 -448
rect -3880 -476 -3842 -448
rect -3814 -476 -3776 -448
rect -3748 -476 -3710 -448
rect -3682 -476 -3644 -448
rect -3616 -476 -3578 -448
rect -3550 -476 -3512 -448
rect -3484 -476 -3446 -448
rect -3418 -476 -3380 -448
rect -3352 -476 -3314 -448
rect -3286 -476 -3248 -448
rect -3220 -476 -3182 -448
rect -3154 -476 -3116 -448
rect -3088 -476 -3050 -448
rect -3022 -476 -2984 -448
rect -2956 -476 -2918 -448
rect -2890 -476 -2852 -448
rect -2824 -476 -2786 -448
rect -2758 -476 -2720 -448
rect -2692 -476 -2654 -448
rect -2626 -476 -2588 -448
rect -2560 -476 -2522 -448
rect -2494 -476 -2456 -448
rect -2428 -476 -2390 -448
rect -2362 -476 -2324 -448
rect -2296 -476 -2258 -448
rect -2230 -476 -2192 -448
rect -2164 -476 -2126 -448
rect -2098 -476 -2060 -448
rect -2032 -476 -1994 -448
rect -1966 -476 -1928 -448
rect -1900 -476 -1862 -448
rect -1834 -476 -1796 -448
rect -1768 -476 -1730 -448
rect -1702 -476 -1664 -448
rect -1636 -476 -1598 -448
rect -1570 -476 -1532 -448
rect -1504 -476 -1466 -448
rect -1438 -476 -1400 -448
rect -1372 -476 -1334 -448
rect -1306 -476 -1268 -448
rect -1240 -476 -1202 -448
rect -1174 -476 -1136 -448
rect -1108 -476 -1070 -448
rect -1042 -476 -1004 -448
rect -976 -476 -938 -448
rect -910 -476 -872 -448
rect -844 -476 -806 -448
rect -778 -476 -740 -448
rect -712 -476 -674 -448
rect -646 -476 -608 -448
rect -580 -476 -542 -448
rect -514 -476 -476 -448
rect -448 -476 -410 -448
rect -382 -476 -344 -448
rect -316 -476 -278 -448
rect -250 -476 -212 -448
rect -184 -476 -146 -448
rect -118 -476 -80 -448
rect -52 -476 -14 -448
rect 14 -476 52 -448
rect 80 -476 118 -448
rect 146 -476 184 -448
rect 212 -476 250 -448
rect 278 -476 316 -448
rect 344 -476 382 -448
rect 410 -476 448 -448
rect 476 -476 514 -448
rect 542 -476 580 -448
rect 608 -476 646 -448
rect 674 -476 712 -448
rect 740 -476 778 -448
rect 806 -476 844 -448
rect 872 -476 910 -448
rect 938 -476 976 -448
rect 1004 -476 1042 -448
rect 1070 -476 1108 -448
rect 1136 -476 1174 -448
rect 1202 -476 1240 -448
rect 1268 -476 1306 -448
rect 1334 -476 1372 -448
rect 1400 -476 1438 -448
rect 1466 -476 1504 -448
rect 1532 -476 1570 -448
rect 1598 -476 1636 -448
rect 1664 -476 1702 -448
rect 1730 -476 1768 -448
rect 1796 -476 1834 -448
rect 1862 -476 1900 -448
rect 1928 -476 1966 -448
rect 1994 -476 2032 -448
rect 2060 -476 2098 -448
rect 2126 -476 2164 -448
rect 2192 -476 2230 -448
rect 2258 -476 2296 -448
rect 2324 -476 2362 -448
rect 2390 -476 2428 -448
rect 2456 -476 2494 -448
rect 2522 -476 2560 -448
rect 2588 -476 2626 -448
rect 2654 -476 2692 -448
rect 2720 -476 2758 -448
rect 2786 -476 2824 -448
rect 2852 -476 2890 -448
rect 2918 -476 2956 -448
rect 2984 -476 3022 -448
rect 3050 -476 3088 -448
rect 3116 -476 3154 -448
rect 3182 -476 3220 -448
rect 3248 -476 3286 -448
rect 3314 -476 3352 -448
rect 3380 -476 3418 -448
rect 3446 -476 3484 -448
rect 3512 -476 3550 -448
rect 3578 -476 3616 -448
rect 3644 -476 3682 -448
rect 3710 -476 3748 -448
rect 3776 -476 3814 -448
rect 3842 -476 3880 -448
rect 3908 -476 3946 -448
rect 3974 -476 4012 -448
rect 4040 -476 4078 -448
rect 4106 -476 4144 -448
rect 4172 -476 4210 -448
rect 4238 -476 4276 -448
rect 4304 -476 4342 -448
rect 4370 -476 4408 -448
rect 4436 -476 4474 -448
rect 4502 -476 4540 -448
rect 4568 -476 4573 -448
rect -4573 -514 4573 -476
rect -4573 -542 -4568 -514
rect -4540 -542 -4502 -514
rect -4474 -542 -4436 -514
rect -4408 -542 -4370 -514
rect -4342 -542 -4304 -514
rect -4276 -542 -4238 -514
rect -4210 -542 -4172 -514
rect -4144 -542 -4106 -514
rect -4078 -542 -4040 -514
rect -4012 -542 -3974 -514
rect -3946 -542 -3908 -514
rect -3880 -542 -3842 -514
rect -3814 -542 -3776 -514
rect -3748 -542 -3710 -514
rect -3682 -542 -3644 -514
rect -3616 -542 -3578 -514
rect -3550 -542 -3512 -514
rect -3484 -542 -3446 -514
rect -3418 -542 -3380 -514
rect -3352 -542 -3314 -514
rect -3286 -542 -3248 -514
rect -3220 -542 -3182 -514
rect -3154 -542 -3116 -514
rect -3088 -542 -3050 -514
rect -3022 -542 -2984 -514
rect -2956 -542 -2918 -514
rect -2890 -542 -2852 -514
rect -2824 -542 -2786 -514
rect -2758 -542 -2720 -514
rect -2692 -542 -2654 -514
rect -2626 -542 -2588 -514
rect -2560 -542 -2522 -514
rect -2494 -542 -2456 -514
rect -2428 -542 -2390 -514
rect -2362 -542 -2324 -514
rect -2296 -542 -2258 -514
rect -2230 -542 -2192 -514
rect -2164 -542 -2126 -514
rect -2098 -542 -2060 -514
rect -2032 -542 -1994 -514
rect -1966 -542 -1928 -514
rect -1900 -542 -1862 -514
rect -1834 -542 -1796 -514
rect -1768 -542 -1730 -514
rect -1702 -542 -1664 -514
rect -1636 -542 -1598 -514
rect -1570 -542 -1532 -514
rect -1504 -542 -1466 -514
rect -1438 -542 -1400 -514
rect -1372 -542 -1334 -514
rect -1306 -542 -1268 -514
rect -1240 -542 -1202 -514
rect -1174 -542 -1136 -514
rect -1108 -542 -1070 -514
rect -1042 -542 -1004 -514
rect -976 -542 -938 -514
rect -910 -542 -872 -514
rect -844 -542 -806 -514
rect -778 -542 -740 -514
rect -712 -542 -674 -514
rect -646 -542 -608 -514
rect -580 -542 -542 -514
rect -514 -542 -476 -514
rect -448 -542 -410 -514
rect -382 -542 -344 -514
rect -316 -542 -278 -514
rect -250 -542 -212 -514
rect -184 -542 -146 -514
rect -118 -542 -80 -514
rect -52 -542 -14 -514
rect 14 -542 52 -514
rect 80 -542 118 -514
rect 146 -542 184 -514
rect 212 -542 250 -514
rect 278 -542 316 -514
rect 344 -542 382 -514
rect 410 -542 448 -514
rect 476 -542 514 -514
rect 542 -542 580 -514
rect 608 -542 646 -514
rect 674 -542 712 -514
rect 740 -542 778 -514
rect 806 -542 844 -514
rect 872 -542 910 -514
rect 938 -542 976 -514
rect 1004 -542 1042 -514
rect 1070 -542 1108 -514
rect 1136 -542 1174 -514
rect 1202 -542 1240 -514
rect 1268 -542 1306 -514
rect 1334 -542 1372 -514
rect 1400 -542 1438 -514
rect 1466 -542 1504 -514
rect 1532 -542 1570 -514
rect 1598 -542 1636 -514
rect 1664 -542 1702 -514
rect 1730 -542 1768 -514
rect 1796 -542 1834 -514
rect 1862 -542 1900 -514
rect 1928 -542 1966 -514
rect 1994 -542 2032 -514
rect 2060 -542 2098 -514
rect 2126 -542 2164 -514
rect 2192 -542 2230 -514
rect 2258 -542 2296 -514
rect 2324 -542 2362 -514
rect 2390 -542 2428 -514
rect 2456 -542 2494 -514
rect 2522 -542 2560 -514
rect 2588 -542 2626 -514
rect 2654 -542 2692 -514
rect 2720 -542 2758 -514
rect 2786 -542 2824 -514
rect 2852 -542 2890 -514
rect 2918 -542 2956 -514
rect 2984 -542 3022 -514
rect 3050 -542 3088 -514
rect 3116 -542 3154 -514
rect 3182 -542 3220 -514
rect 3248 -542 3286 -514
rect 3314 -542 3352 -514
rect 3380 -542 3418 -514
rect 3446 -542 3484 -514
rect 3512 -542 3550 -514
rect 3578 -542 3616 -514
rect 3644 -542 3682 -514
rect 3710 -542 3748 -514
rect 3776 -542 3814 -514
rect 3842 -542 3880 -514
rect 3908 -542 3946 -514
rect 3974 -542 4012 -514
rect 4040 -542 4078 -514
rect 4106 -542 4144 -514
rect 4172 -542 4210 -514
rect 4238 -542 4276 -514
rect 4304 -542 4342 -514
rect 4370 -542 4408 -514
rect 4436 -542 4474 -514
rect 4502 -542 4540 -514
rect 4568 -542 4573 -514
rect -4573 -580 4573 -542
rect -4573 -608 -4568 -580
rect -4540 -608 -4502 -580
rect -4474 -608 -4436 -580
rect -4408 -608 -4370 -580
rect -4342 -608 -4304 -580
rect -4276 -608 -4238 -580
rect -4210 -608 -4172 -580
rect -4144 -608 -4106 -580
rect -4078 -608 -4040 -580
rect -4012 -608 -3974 -580
rect -3946 -608 -3908 -580
rect -3880 -608 -3842 -580
rect -3814 -608 -3776 -580
rect -3748 -608 -3710 -580
rect -3682 -608 -3644 -580
rect -3616 -608 -3578 -580
rect -3550 -608 -3512 -580
rect -3484 -608 -3446 -580
rect -3418 -608 -3380 -580
rect -3352 -608 -3314 -580
rect -3286 -608 -3248 -580
rect -3220 -608 -3182 -580
rect -3154 -608 -3116 -580
rect -3088 -608 -3050 -580
rect -3022 -608 -2984 -580
rect -2956 -608 -2918 -580
rect -2890 -608 -2852 -580
rect -2824 -608 -2786 -580
rect -2758 -608 -2720 -580
rect -2692 -608 -2654 -580
rect -2626 -608 -2588 -580
rect -2560 -608 -2522 -580
rect -2494 -608 -2456 -580
rect -2428 -608 -2390 -580
rect -2362 -608 -2324 -580
rect -2296 -608 -2258 -580
rect -2230 -608 -2192 -580
rect -2164 -608 -2126 -580
rect -2098 -608 -2060 -580
rect -2032 -608 -1994 -580
rect -1966 -608 -1928 -580
rect -1900 -608 -1862 -580
rect -1834 -608 -1796 -580
rect -1768 -608 -1730 -580
rect -1702 -608 -1664 -580
rect -1636 -608 -1598 -580
rect -1570 -608 -1532 -580
rect -1504 -608 -1466 -580
rect -1438 -608 -1400 -580
rect -1372 -608 -1334 -580
rect -1306 -608 -1268 -580
rect -1240 -608 -1202 -580
rect -1174 -608 -1136 -580
rect -1108 -608 -1070 -580
rect -1042 -608 -1004 -580
rect -976 -608 -938 -580
rect -910 -608 -872 -580
rect -844 -608 -806 -580
rect -778 -608 -740 -580
rect -712 -608 -674 -580
rect -646 -608 -608 -580
rect -580 -608 -542 -580
rect -514 -608 -476 -580
rect -448 -608 -410 -580
rect -382 -608 -344 -580
rect -316 -608 -278 -580
rect -250 -608 -212 -580
rect -184 -608 -146 -580
rect -118 -608 -80 -580
rect -52 -608 -14 -580
rect 14 -608 52 -580
rect 80 -608 118 -580
rect 146 -608 184 -580
rect 212 -608 250 -580
rect 278 -608 316 -580
rect 344 -608 382 -580
rect 410 -608 448 -580
rect 476 -608 514 -580
rect 542 -608 580 -580
rect 608 -608 646 -580
rect 674 -608 712 -580
rect 740 -608 778 -580
rect 806 -608 844 -580
rect 872 -608 910 -580
rect 938 -608 976 -580
rect 1004 -608 1042 -580
rect 1070 -608 1108 -580
rect 1136 -608 1174 -580
rect 1202 -608 1240 -580
rect 1268 -608 1306 -580
rect 1334 -608 1372 -580
rect 1400 -608 1438 -580
rect 1466 -608 1504 -580
rect 1532 -608 1570 -580
rect 1598 -608 1636 -580
rect 1664 -608 1702 -580
rect 1730 -608 1768 -580
rect 1796 -608 1834 -580
rect 1862 -608 1900 -580
rect 1928 -608 1966 -580
rect 1994 -608 2032 -580
rect 2060 -608 2098 -580
rect 2126 -608 2164 -580
rect 2192 -608 2230 -580
rect 2258 -608 2296 -580
rect 2324 -608 2362 -580
rect 2390 -608 2428 -580
rect 2456 -608 2494 -580
rect 2522 -608 2560 -580
rect 2588 -608 2626 -580
rect 2654 -608 2692 -580
rect 2720 -608 2758 -580
rect 2786 -608 2824 -580
rect 2852 -608 2890 -580
rect 2918 -608 2956 -580
rect 2984 -608 3022 -580
rect 3050 -608 3088 -580
rect 3116 -608 3154 -580
rect 3182 -608 3220 -580
rect 3248 -608 3286 -580
rect 3314 -608 3352 -580
rect 3380 -608 3418 -580
rect 3446 -608 3484 -580
rect 3512 -608 3550 -580
rect 3578 -608 3616 -580
rect 3644 -608 3682 -580
rect 3710 -608 3748 -580
rect 3776 -608 3814 -580
rect 3842 -608 3880 -580
rect 3908 -608 3946 -580
rect 3974 -608 4012 -580
rect 4040 -608 4078 -580
rect 4106 -608 4144 -580
rect 4172 -608 4210 -580
rect 4238 -608 4276 -580
rect 4304 -608 4342 -580
rect 4370 -608 4408 -580
rect 4436 -608 4474 -580
rect 4502 -608 4540 -580
rect 4568 -608 4573 -580
rect -4573 -646 4573 -608
rect -4573 -674 -4568 -646
rect -4540 -674 -4502 -646
rect -4474 -674 -4436 -646
rect -4408 -674 -4370 -646
rect -4342 -674 -4304 -646
rect -4276 -674 -4238 -646
rect -4210 -674 -4172 -646
rect -4144 -674 -4106 -646
rect -4078 -674 -4040 -646
rect -4012 -674 -3974 -646
rect -3946 -674 -3908 -646
rect -3880 -674 -3842 -646
rect -3814 -674 -3776 -646
rect -3748 -674 -3710 -646
rect -3682 -674 -3644 -646
rect -3616 -674 -3578 -646
rect -3550 -674 -3512 -646
rect -3484 -674 -3446 -646
rect -3418 -674 -3380 -646
rect -3352 -674 -3314 -646
rect -3286 -674 -3248 -646
rect -3220 -674 -3182 -646
rect -3154 -674 -3116 -646
rect -3088 -674 -3050 -646
rect -3022 -674 -2984 -646
rect -2956 -674 -2918 -646
rect -2890 -674 -2852 -646
rect -2824 -674 -2786 -646
rect -2758 -674 -2720 -646
rect -2692 -674 -2654 -646
rect -2626 -674 -2588 -646
rect -2560 -674 -2522 -646
rect -2494 -674 -2456 -646
rect -2428 -674 -2390 -646
rect -2362 -674 -2324 -646
rect -2296 -674 -2258 -646
rect -2230 -674 -2192 -646
rect -2164 -674 -2126 -646
rect -2098 -674 -2060 -646
rect -2032 -674 -1994 -646
rect -1966 -674 -1928 -646
rect -1900 -674 -1862 -646
rect -1834 -674 -1796 -646
rect -1768 -674 -1730 -646
rect -1702 -674 -1664 -646
rect -1636 -674 -1598 -646
rect -1570 -674 -1532 -646
rect -1504 -674 -1466 -646
rect -1438 -674 -1400 -646
rect -1372 -674 -1334 -646
rect -1306 -674 -1268 -646
rect -1240 -674 -1202 -646
rect -1174 -674 -1136 -646
rect -1108 -674 -1070 -646
rect -1042 -674 -1004 -646
rect -976 -674 -938 -646
rect -910 -674 -872 -646
rect -844 -674 -806 -646
rect -778 -674 -740 -646
rect -712 -674 -674 -646
rect -646 -674 -608 -646
rect -580 -674 -542 -646
rect -514 -674 -476 -646
rect -448 -674 -410 -646
rect -382 -674 -344 -646
rect -316 -674 -278 -646
rect -250 -674 -212 -646
rect -184 -674 -146 -646
rect -118 -674 -80 -646
rect -52 -674 -14 -646
rect 14 -674 52 -646
rect 80 -674 118 -646
rect 146 -674 184 -646
rect 212 -674 250 -646
rect 278 -674 316 -646
rect 344 -674 382 -646
rect 410 -674 448 -646
rect 476 -674 514 -646
rect 542 -674 580 -646
rect 608 -674 646 -646
rect 674 -674 712 -646
rect 740 -674 778 -646
rect 806 -674 844 -646
rect 872 -674 910 -646
rect 938 -674 976 -646
rect 1004 -674 1042 -646
rect 1070 -674 1108 -646
rect 1136 -674 1174 -646
rect 1202 -674 1240 -646
rect 1268 -674 1306 -646
rect 1334 -674 1372 -646
rect 1400 -674 1438 -646
rect 1466 -674 1504 -646
rect 1532 -674 1570 -646
rect 1598 -674 1636 -646
rect 1664 -674 1702 -646
rect 1730 -674 1768 -646
rect 1796 -674 1834 -646
rect 1862 -674 1900 -646
rect 1928 -674 1966 -646
rect 1994 -674 2032 -646
rect 2060 -674 2098 -646
rect 2126 -674 2164 -646
rect 2192 -674 2230 -646
rect 2258 -674 2296 -646
rect 2324 -674 2362 -646
rect 2390 -674 2428 -646
rect 2456 -674 2494 -646
rect 2522 -674 2560 -646
rect 2588 -674 2626 -646
rect 2654 -674 2692 -646
rect 2720 -674 2758 -646
rect 2786 -674 2824 -646
rect 2852 -674 2890 -646
rect 2918 -674 2956 -646
rect 2984 -674 3022 -646
rect 3050 -674 3088 -646
rect 3116 -674 3154 -646
rect 3182 -674 3220 -646
rect 3248 -674 3286 -646
rect 3314 -674 3352 -646
rect 3380 -674 3418 -646
rect 3446 -674 3484 -646
rect 3512 -674 3550 -646
rect 3578 -674 3616 -646
rect 3644 -674 3682 -646
rect 3710 -674 3748 -646
rect 3776 -674 3814 -646
rect 3842 -674 3880 -646
rect 3908 -674 3946 -646
rect 3974 -674 4012 -646
rect 4040 -674 4078 -646
rect 4106 -674 4144 -646
rect 4172 -674 4210 -646
rect 4238 -674 4276 -646
rect 4304 -674 4342 -646
rect 4370 -674 4408 -646
rect 4436 -674 4474 -646
rect 4502 -674 4540 -646
rect 4568 -674 4573 -646
rect -4573 -712 4573 -674
rect -4573 -740 -4568 -712
rect -4540 -740 -4502 -712
rect -4474 -740 -4436 -712
rect -4408 -740 -4370 -712
rect -4342 -740 -4304 -712
rect -4276 -740 -4238 -712
rect -4210 -740 -4172 -712
rect -4144 -740 -4106 -712
rect -4078 -740 -4040 -712
rect -4012 -740 -3974 -712
rect -3946 -740 -3908 -712
rect -3880 -740 -3842 -712
rect -3814 -740 -3776 -712
rect -3748 -740 -3710 -712
rect -3682 -740 -3644 -712
rect -3616 -740 -3578 -712
rect -3550 -740 -3512 -712
rect -3484 -740 -3446 -712
rect -3418 -740 -3380 -712
rect -3352 -740 -3314 -712
rect -3286 -740 -3248 -712
rect -3220 -740 -3182 -712
rect -3154 -740 -3116 -712
rect -3088 -740 -3050 -712
rect -3022 -740 -2984 -712
rect -2956 -740 -2918 -712
rect -2890 -740 -2852 -712
rect -2824 -740 -2786 -712
rect -2758 -740 -2720 -712
rect -2692 -740 -2654 -712
rect -2626 -740 -2588 -712
rect -2560 -740 -2522 -712
rect -2494 -740 -2456 -712
rect -2428 -740 -2390 -712
rect -2362 -740 -2324 -712
rect -2296 -740 -2258 -712
rect -2230 -740 -2192 -712
rect -2164 -740 -2126 -712
rect -2098 -740 -2060 -712
rect -2032 -740 -1994 -712
rect -1966 -740 -1928 -712
rect -1900 -740 -1862 -712
rect -1834 -740 -1796 -712
rect -1768 -740 -1730 -712
rect -1702 -740 -1664 -712
rect -1636 -740 -1598 -712
rect -1570 -740 -1532 -712
rect -1504 -740 -1466 -712
rect -1438 -740 -1400 -712
rect -1372 -740 -1334 -712
rect -1306 -740 -1268 -712
rect -1240 -740 -1202 -712
rect -1174 -740 -1136 -712
rect -1108 -740 -1070 -712
rect -1042 -740 -1004 -712
rect -976 -740 -938 -712
rect -910 -740 -872 -712
rect -844 -740 -806 -712
rect -778 -740 -740 -712
rect -712 -740 -674 -712
rect -646 -740 -608 -712
rect -580 -740 -542 -712
rect -514 -740 -476 -712
rect -448 -740 -410 -712
rect -382 -740 -344 -712
rect -316 -740 -278 -712
rect -250 -740 -212 -712
rect -184 -740 -146 -712
rect -118 -740 -80 -712
rect -52 -740 -14 -712
rect 14 -740 52 -712
rect 80 -740 118 -712
rect 146 -740 184 -712
rect 212 -740 250 -712
rect 278 -740 316 -712
rect 344 -740 382 -712
rect 410 -740 448 -712
rect 476 -740 514 -712
rect 542 -740 580 -712
rect 608 -740 646 -712
rect 674 -740 712 -712
rect 740 -740 778 -712
rect 806 -740 844 -712
rect 872 -740 910 -712
rect 938 -740 976 -712
rect 1004 -740 1042 -712
rect 1070 -740 1108 -712
rect 1136 -740 1174 -712
rect 1202 -740 1240 -712
rect 1268 -740 1306 -712
rect 1334 -740 1372 -712
rect 1400 -740 1438 -712
rect 1466 -740 1504 -712
rect 1532 -740 1570 -712
rect 1598 -740 1636 -712
rect 1664 -740 1702 -712
rect 1730 -740 1768 -712
rect 1796 -740 1834 -712
rect 1862 -740 1900 -712
rect 1928 -740 1966 -712
rect 1994 -740 2032 -712
rect 2060 -740 2098 -712
rect 2126 -740 2164 -712
rect 2192 -740 2230 -712
rect 2258 -740 2296 -712
rect 2324 -740 2362 -712
rect 2390 -740 2428 -712
rect 2456 -740 2494 -712
rect 2522 -740 2560 -712
rect 2588 -740 2626 -712
rect 2654 -740 2692 -712
rect 2720 -740 2758 -712
rect 2786 -740 2824 -712
rect 2852 -740 2890 -712
rect 2918 -740 2956 -712
rect 2984 -740 3022 -712
rect 3050 -740 3088 -712
rect 3116 -740 3154 -712
rect 3182 -740 3220 -712
rect 3248 -740 3286 -712
rect 3314 -740 3352 -712
rect 3380 -740 3418 -712
rect 3446 -740 3484 -712
rect 3512 -740 3550 -712
rect 3578 -740 3616 -712
rect 3644 -740 3682 -712
rect 3710 -740 3748 -712
rect 3776 -740 3814 -712
rect 3842 -740 3880 -712
rect 3908 -740 3946 -712
rect 3974 -740 4012 -712
rect 4040 -740 4078 -712
rect 4106 -740 4144 -712
rect 4172 -740 4210 -712
rect 4238 -740 4276 -712
rect 4304 -740 4342 -712
rect 4370 -740 4408 -712
rect 4436 -740 4474 -712
rect 4502 -740 4540 -712
rect 4568 -740 4573 -712
rect -4573 -745 4573 -740
<< via3 >>
rect -4568 712 -4540 740
rect -4502 712 -4474 740
rect -4436 712 -4408 740
rect -4370 712 -4342 740
rect -4304 712 -4276 740
rect -4238 712 -4210 740
rect -4172 712 -4144 740
rect -4106 712 -4078 740
rect -4040 712 -4012 740
rect -3974 712 -3946 740
rect -3908 712 -3880 740
rect -3842 712 -3814 740
rect -3776 712 -3748 740
rect -3710 712 -3682 740
rect -3644 712 -3616 740
rect -3578 712 -3550 740
rect -3512 712 -3484 740
rect -3446 712 -3418 740
rect -3380 712 -3352 740
rect -3314 712 -3286 740
rect -3248 712 -3220 740
rect -3182 712 -3154 740
rect -3116 712 -3088 740
rect -3050 712 -3022 740
rect -2984 712 -2956 740
rect -2918 712 -2890 740
rect -2852 712 -2824 740
rect -2786 712 -2758 740
rect -2720 712 -2692 740
rect -2654 712 -2626 740
rect -2588 712 -2560 740
rect -2522 712 -2494 740
rect -2456 712 -2428 740
rect -2390 712 -2362 740
rect -2324 712 -2296 740
rect -2258 712 -2230 740
rect -2192 712 -2164 740
rect -2126 712 -2098 740
rect -2060 712 -2032 740
rect -1994 712 -1966 740
rect -1928 712 -1900 740
rect -1862 712 -1834 740
rect -1796 712 -1768 740
rect -1730 712 -1702 740
rect -1664 712 -1636 740
rect -1598 712 -1570 740
rect -1532 712 -1504 740
rect -1466 712 -1438 740
rect -1400 712 -1372 740
rect -1334 712 -1306 740
rect -1268 712 -1240 740
rect -1202 712 -1174 740
rect -1136 712 -1108 740
rect -1070 712 -1042 740
rect -1004 712 -976 740
rect -938 712 -910 740
rect -872 712 -844 740
rect -806 712 -778 740
rect -740 712 -712 740
rect -674 712 -646 740
rect -608 712 -580 740
rect -542 712 -514 740
rect -476 712 -448 740
rect -410 712 -382 740
rect -344 712 -316 740
rect -278 712 -250 740
rect -212 712 -184 740
rect -146 712 -118 740
rect -80 712 -52 740
rect -14 712 14 740
rect 52 712 80 740
rect 118 712 146 740
rect 184 712 212 740
rect 250 712 278 740
rect 316 712 344 740
rect 382 712 410 740
rect 448 712 476 740
rect 514 712 542 740
rect 580 712 608 740
rect 646 712 674 740
rect 712 712 740 740
rect 778 712 806 740
rect 844 712 872 740
rect 910 712 938 740
rect 976 712 1004 740
rect 1042 712 1070 740
rect 1108 712 1136 740
rect 1174 712 1202 740
rect 1240 712 1268 740
rect 1306 712 1334 740
rect 1372 712 1400 740
rect 1438 712 1466 740
rect 1504 712 1532 740
rect 1570 712 1598 740
rect 1636 712 1664 740
rect 1702 712 1730 740
rect 1768 712 1796 740
rect 1834 712 1862 740
rect 1900 712 1928 740
rect 1966 712 1994 740
rect 2032 712 2060 740
rect 2098 712 2126 740
rect 2164 712 2192 740
rect 2230 712 2258 740
rect 2296 712 2324 740
rect 2362 712 2390 740
rect 2428 712 2456 740
rect 2494 712 2522 740
rect 2560 712 2588 740
rect 2626 712 2654 740
rect 2692 712 2720 740
rect 2758 712 2786 740
rect 2824 712 2852 740
rect 2890 712 2918 740
rect 2956 712 2984 740
rect 3022 712 3050 740
rect 3088 712 3116 740
rect 3154 712 3182 740
rect 3220 712 3248 740
rect 3286 712 3314 740
rect 3352 712 3380 740
rect 3418 712 3446 740
rect 3484 712 3512 740
rect 3550 712 3578 740
rect 3616 712 3644 740
rect 3682 712 3710 740
rect 3748 712 3776 740
rect 3814 712 3842 740
rect 3880 712 3908 740
rect 3946 712 3974 740
rect 4012 712 4040 740
rect 4078 712 4106 740
rect 4144 712 4172 740
rect 4210 712 4238 740
rect 4276 712 4304 740
rect 4342 712 4370 740
rect 4408 712 4436 740
rect 4474 712 4502 740
rect 4540 712 4568 740
rect -4568 646 -4540 674
rect -4502 646 -4474 674
rect -4436 646 -4408 674
rect -4370 646 -4342 674
rect -4304 646 -4276 674
rect -4238 646 -4210 674
rect -4172 646 -4144 674
rect -4106 646 -4078 674
rect -4040 646 -4012 674
rect -3974 646 -3946 674
rect -3908 646 -3880 674
rect -3842 646 -3814 674
rect -3776 646 -3748 674
rect -3710 646 -3682 674
rect -3644 646 -3616 674
rect -3578 646 -3550 674
rect -3512 646 -3484 674
rect -3446 646 -3418 674
rect -3380 646 -3352 674
rect -3314 646 -3286 674
rect -3248 646 -3220 674
rect -3182 646 -3154 674
rect -3116 646 -3088 674
rect -3050 646 -3022 674
rect -2984 646 -2956 674
rect -2918 646 -2890 674
rect -2852 646 -2824 674
rect -2786 646 -2758 674
rect -2720 646 -2692 674
rect -2654 646 -2626 674
rect -2588 646 -2560 674
rect -2522 646 -2494 674
rect -2456 646 -2428 674
rect -2390 646 -2362 674
rect -2324 646 -2296 674
rect -2258 646 -2230 674
rect -2192 646 -2164 674
rect -2126 646 -2098 674
rect -2060 646 -2032 674
rect -1994 646 -1966 674
rect -1928 646 -1900 674
rect -1862 646 -1834 674
rect -1796 646 -1768 674
rect -1730 646 -1702 674
rect -1664 646 -1636 674
rect -1598 646 -1570 674
rect -1532 646 -1504 674
rect -1466 646 -1438 674
rect -1400 646 -1372 674
rect -1334 646 -1306 674
rect -1268 646 -1240 674
rect -1202 646 -1174 674
rect -1136 646 -1108 674
rect -1070 646 -1042 674
rect -1004 646 -976 674
rect -938 646 -910 674
rect -872 646 -844 674
rect -806 646 -778 674
rect -740 646 -712 674
rect -674 646 -646 674
rect -608 646 -580 674
rect -542 646 -514 674
rect -476 646 -448 674
rect -410 646 -382 674
rect -344 646 -316 674
rect -278 646 -250 674
rect -212 646 -184 674
rect -146 646 -118 674
rect -80 646 -52 674
rect -14 646 14 674
rect 52 646 80 674
rect 118 646 146 674
rect 184 646 212 674
rect 250 646 278 674
rect 316 646 344 674
rect 382 646 410 674
rect 448 646 476 674
rect 514 646 542 674
rect 580 646 608 674
rect 646 646 674 674
rect 712 646 740 674
rect 778 646 806 674
rect 844 646 872 674
rect 910 646 938 674
rect 976 646 1004 674
rect 1042 646 1070 674
rect 1108 646 1136 674
rect 1174 646 1202 674
rect 1240 646 1268 674
rect 1306 646 1334 674
rect 1372 646 1400 674
rect 1438 646 1466 674
rect 1504 646 1532 674
rect 1570 646 1598 674
rect 1636 646 1664 674
rect 1702 646 1730 674
rect 1768 646 1796 674
rect 1834 646 1862 674
rect 1900 646 1928 674
rect 1966 646 1994 674
rect 2032 646 2060 674
rect 2098 646 2126 674
rect 2164 646 2192 674
rect 2230 646 2258 674
rect 2296 646 2324 674
rect 2362 646 2390 674
rect 2428 646 2456 674
rect 2494 646 2522 674
rect 2560 646 2588 674
rect 2626 646 2654 674
rect 2692 646 2720 674
rect 2758 646 2786 674
rect 2824 646 2852 674
rect 2890 646 2918 674
rect 2956 646 2984 674
rect 3022 646 3050 674
rect 3088 646 3116 674
rect 3154 646 3182 674
rect 3220 646 3248 674
rect 3286 646 3314 674
rect 3352 646 3380 674
rect 3418 646 3446 674
rect 3484 646 3512 674
rect 3550 646 3578 674
rect 3616 646 3644 674
rect 3682 646 3710 674
rect 3748 646 3776 674
rect 3814 646 3842 674
rect 3880 646 3908 674
rect 3946 646 3974 674
rect 4012 646 4040 674
rect 4078 646 4106 674
rect 4144 646 4172 674
rect 4210 646 4238 674
rect 4276 646 4304 674
rect 4342 646 4370 674
rect 4408 646 4436 674
rect 4474 646 4502 674
rect 4540 646 4568 674
rect -4568 580 -4540 608
rect -4502 580 -4474 608
rect -4436 580 -4408 608
rect -4370 580 -4342 608
rect -4304 580 -4276 608
rect -4238 580 -4210 608
rect -4172 580 -4144 608
rect -4106 580 -4078 608
rect -4040 580 -4012 608
rect -3974 580 -3946 608
rect -3908 580 -3880 608
rect -3842 580 -3814 608
rect -3776 580 -3748 608
rect -3710 580 -3682 608
rect -3644 580 -3616 608
rect -3578 580 -3550 608
rect -3512 580 -3484 608
rect -3446 580 -3418 608
rect -3380 580 -3352 608
rect -3314 580 -3286 608
rect -3248 580 -3220 608
rect -3182 580 -3154 608
rect -3116 580 -3088 608
rect -3050 580 -3022 608
rect -2984 580 -2956 608
rect -2918 580 -2890 608
rect -2852 580 -2824 608
rect -2786 580 -2758 608
rect -2720 580 -2692 608
rect -2654 580 -2626 608
rect -2588 580 -2560 608
rect -2522 580 -2494 608
rect -2456 580 -2428 608
rect -2390 580 -2362 608
rect -2324 580 -2296 608
rect -2258 580 -2230 608
rect -2192 580 -2164 608
rect -2126 580 -2098 608
rect -2060 580 -2032 608
rect -1994 580 -1966 608
rect -1928 580 -1900 608
rect -1862 580 -1834 608
rect -1796 580 -1768 608
rect -1730 580 -1702 608
rect -1664 580 -1636 608
rect -1598 580 -1570 608
rect -1532 580 -1504 608
rect -1466 580 -1438 608
rect -1400 580 -1372 608
rect -1334 580 -1306 608
rect -1268 580 -1240 608
rect -1202 580 -1174 608
rect -1136 580 -1108 608
rect -1070 580 -1042 608
rect -1004 580 -976 608
rect -938 580 -910 608
rect -872 580 -844 608
rect -806 580 -778 608
rect -740 580 -712 608
rect -674 580 -646 608
rect -608 580 -580 608
rect -542 580 -514 608
rect -476 580 -448 608
rect -410 580 -382 608
rect -344 580 -316 608
rect -278 580 -250 608
rect -212 580 -184 608
rect -146 580 -118 608
rect -80 580 -52 608
rect -14 580 14 608
rect 52 580 80 608
rect 118 580 146 608
rect 184 580 212 608
rect 250 580 278 608
rect 316 580 344 608
rect 382 580 410 608
rect 448 580 476 608
rect 514 580 542 608
rect 580 580 608 608
rect 646 580 674 608
rect 712 580 740 608
rect 778 580 806 608
rect 844 580 872 608
rect 910 580 938 608
rect 976 580 1004 608
rect 1042 580 1070 608
rect 1108 580 1136 608
rect 1174 580 1202 608
rect 1240 580 1268 608
rect 1306 580 1334 608
rect 1372 580 1400 608
rect 1438 580 1466 608
rect 1504 580 1532 608
rect 1570 580 1598 608
rect 1636 580 1664 608
rect 1702 580 1730 608
rect 1768 580 1796 608
rect 1834 580 1862 608
rect 1900 580 1928 608
rect 1966 580 1994 608
rect 2032 580 2060 608
rect 2098 580 2126 608
rect 2164 580 2192 608
rect 2230 580 2258 608
rect 2296 580 2324 608
rect 2362 580 2390 608
rect 2428 580 2456 608
rect 2494 580 2522 608
rect 2560 580 2588 608
rect 2626 580 2654 608
rect 2692 580 2720 608
rect 2758 580 2786 608
rect 2824 580 2852 608
rect 2890 580 2918 608
rect 2956 580 2984 608
rect 3022 580 3050 608
rect 3088 580 3116 608
rect 3154 580 3182 608
rect 3220 580 3248 608
rect 3286 580 3314 608
rect 3352 580 3380 608
rect 3418 580 3446 608
rect 3484 580 3512 608
rect 3550 580 3578 608
rect 3616 580 3644 608
rect 3682 580 3710 608
rect 3748 580 3776 608
rect 3814 580 3842 608
rect 3880 580 3908 608
rect 3946 580 3974 608
rect 4012 580 4040 608
rect 4078 580 4106 608
rect 4144 580 4172 608
rect 4210 580 4238 608
rect 4276 580 4304 608
rect 4342 580 4370 608
rect 4408 580 4436 608
rect 4474 580 4502 608
rect 4540 580 4568 608
rect -4568 514 -4540 542
rect -4502 514 -4474 542
rect -4436 514 -4408 542
rect -4370 514 -4342 542
rect -4304 514 -4276 542
rect -4238 514 -4210 542
rect -4172 514 -4144 542
rect -4106 514 -4078 542
rect -4040 514 -4012 542
rect -3974 514 -3946 542
rect -3908 514 -3880 542
rect -3842 514 -3814 542
rect -3776 514 -3748 542
rect -3710 514 -3682 542
rect -3644 514 -3616 542
rect -3578 514 -3550 542
rect -3512 514 -3484 542
rect -3446 514 -3418 542
rect -3380 514 -3352 542
rect -3314 514 -3286 542
rect -3248 514 -3220 542
rect -3182 514 -3154 542
rect -3116 514 -3088 542
rect -3050 514 -3022 542
rect -2984 514 -2956 542
rect -2918 514 -2890 542
rect -2852 514 -2824 542
rect -2786 514 -2758 542
rect -2720 514 -2692 542
rect -2654 514 -2626 542
rect -2588 514 -2560 542
rect -2522 514 -2494 542
rect -2456 514 -2428 542
rect -2390 514 -2362 542
rect -2324 514 -2296 542
rect -2258 514 -2230 542
rect -2192 514 -2164 542
rect -2126 514 -2098 542
rect -2060 514 -2032 542
rect -1994 514 -1966 542
rect -1928 514 -1900 542
rect -1862 514 -1834 542
rect -1796 514 -1768 542
rect -1730 514 -1702 542
rect -1664 514 -1636 542
rect -1598 514 -1570 542
rect -1532 514 -1504 542
rect -1466 514 -1438 542
rect -1400 514 -1372 542
rect -1334 514 -1306 542
rect -1268 514 -1240 542
rect -1202 514 -1174 542
rect -1136 514 -1108 542
rect -1070 514 -1042 542
rect -1004 514 -976 542
rect -938 514 -910 542
rect -872 514 -844 542
rect -806 514 -778 542
rect -740 514 -712 542
rect -674 514 -646 542
rect -608 514 -580 542
rect -542 514 -514 542
rect -476 514 -448 542
rect -410 514 -382 542
rect -344 514 -316 542
rect -278 514 -250 542
rect -212 514 -184 542
rect -146 514 -118 542
rect -80 514 -52 542
rect -14 514 14 542
rect 52 514 80 542
rect 118 514 146 542
rect 184 514 212 542
rect 250 514 278 542
rect 316 514 344 542
rect 382 514 410 542
rect 448 514 476 542
rect 514 514 542 542
rect 580 514 608 542
rect 646 514 674 542
rect 712 514 740 542
rect 778 514 806 542
rect 844 514 872 542
rect 910 514 938 542
rect 976 514 1004 542
rect 1042 514 1070 542
rect 1108 514 1136 542
rect 1174 514 1202 542
rect 1240 514 1268 542
rect 1306 514 1334 542
rect 1372 514 1400 542
rect 1438 514 1466 542
rect 1504 514 1532 542
rect 1570 514 1598 542
rect 1636 514 1664 542
rect 1702 514 1730 542
rect 1768 514 1796 542
rect 1834 514 1862 542
rect 1900 514 1928 542
rect 1966 514 1994 542
rect 2032 514 2060 542
rect 2098 514 2126 542
rect 2164 514 2192 542
rect 2230 514 2258 542
rect 2296 514 2324 542
rect 2362 514 2390 542
rect 2428 514 2456 542
rect 2494 514 2522 542
rect 2560 514 2588 542
rect 2626 514 2654 542
rect 2692 514 2720 542
rect 2758 514 2786 542
rect 2824 514 2852 542
rect 2890 514 2918 542
rect 2956 514 2984 542
rect 3022 514 3050 542
rect 3088 514 3116 542
rect 3154 514 3182 542
rect 3220 514 3248 542
rect 3286 514 3314 542
rect 3352 514 3380 542
rect 3418 514 3446 542
rect 3484 514 3512 542
rect 3550 514 3578 542
rect 3616 514 3644 542
rect 3682 514 3710 542
rect 3748 514 3776 542
rect 3814 514 3842 542
rect 3880 514 3908 542
rect 3946 514 3974 542
rect 4012 514 4040 542
rect 4078 514 4106 542
rect 4144 514 4172 542
rect 4210 514 4238 542
rect 4276 514 4304 542
rect 4342 514 4370 542
rect 4408 514 4436 542
rect 4474 514 4502 542
rect 4540 514 4568 542
rect -4568 448 -4540 476
rect -4502 448 -4474 476
rect -4436 448 -4408 476
rect -4370 448 -4342 476
rect -4304 448 -4276 476
rect -4238 448 -4210 476
rect -4172 448 -4144 476
rect -4106 448 -4078 476
rect -4040 448 -4012 476
rect -3974 448 -3946 476
rect -3908 448 -3880 476
rect -3842 448 -3814 476
rect -3776 448 -3748 476
rect -3710 448 -3682 476
rect -3644 448 -3616 476
rect -3578 448 -3550 476
rect -3512 448 -3484 476
rect -3446 448 -3418 476
rect -3380 448 -3352 476
rect -3314 448 -3286 476
rect -3248 448 -3220 476
rect -3182 448 -3154 476
rect -3116 448 -3088 476
rect -3050 448 -3022 476
rect -2984 448 -2956 476
rect -2918 448 -2890 476
rect -2852 448 -2824 476
rect -2786 448 -2758 476
rect -2720 448 -2692 476
rect -2654 448 -2626 476
rect -2588 448 -2560 476
rect -2522 448 -2494 476
rect -2456 448 -2428 476
rect -2390 448 -2362 476
rect -2324 448 -2296 476
rect -2258 448 -2230 476
rect -2192 448 -2164 476
rect -2126 448 -2098 476
rect -2060 448 -2032 476
rect -1994 448 -1966 476
rect -1928 448 -1900 476
rect -1862 448 -1834 476
rect -1796 448 -1768 476
rect -1730 448 -1702 476
rect -1664 448 -1636 476
rect -1598 448 -1570 476
rect -1532 448 -1504 476
rect -1466 448 -1438 476
rect -1400 448 -1372 476
rect -1334 448 -1306 476
rect -1268 448 -1240 476
rect -1202 448 -1174 476
rect -1136 448 -1108 476
rect -1070 448 -1042 476
rect -1004 448 -976 476
rect -938 448 -910 476
rect -872 448 -844 476
rect -806 448 -778 476
rect -740 448 -712 476
rect -674 448 -646 476
rect -608 448 -580 476
rect -542 448 -514 476
rect -476 448 -448 476
rect -410 448 -382 476
rect -344 448 -316 476
rect -278 448 -250 476
rect -212 448 -184 476
rect -146 448 -118 476
rect -80 448 -52 476
rect -14 448 14 476
rect 52 448 80 476
rect 118 448 146 476
rect 184 448 212 476
rect 250 448 278 476
rect 316 448 344 476
rect 382 448 410 476
rect 448 448 476 476
rect 514 448 542 476
rect 580 448 608 476
rect 646 448 674 476
rect 712 448 740 476
rect 778 448 806 476
rect 844 448 872 476
rect 910 448 938 476
rect 976 448 1004 476
rect 1042 448 1070 476
rect 1108 448 1136 476
rect 1174 448 1202 476
rect 1240 448 1268 476
rect 1306 448 1334 476
rect 1372 448 1400 476
rect 1438 448 1466 476
rect 1504 448 1532 476
rect 1570 448 1598 476
rect 1636 448 1664 476
rect 1702 448 1730 476
rect 1768 448 1796 476
rect 1834 448 1862 476
rect 1900 448 1928 476
rect 1966 448 1994 476
rect 2032 448 2060 476
rect 2098 448 2126 476
rect 2164 448 2192 476
rect 2230 448 2258 476
rect 2296 448 2324 476
rect 2362 448 2390 476
rect 2428 448 2456 476
rect 2494 448 2522 476
rect 2560 448 2588 476
rect 2626 448 2654 476
rect 2692 448 2720 476
rect 2758 448 2786 476
rect 2824 448 2852 476
rect 2890 448 2918 476
rect 2956 448 2984 476
rect 3022 448 3050 476
rect 3088 448 3116 476
rect 3154 448 3182 476
rect 3220 448 3248 476
rect 3286 448 3314 476
rect 3352 448 3380 476
rect 3418 448 3446 476
rect 3484 448 3512 476
rect 3550 448 3578 476
rect 3616 448 3644 476
rect 3682 448 3710 476
rect 3748 448 3776 476
rect 3814 448 3842 476
rect 3880 448 3908 476
rect 3946 448 3974 476
rect 4012 448 4040 476
rect 4078 448 4106 476
rect 4144 448 4172 476
rect 4210 448 4238 476
rect 4276 448 4304 476
rect 4342 448 4370 476
rect 4408 448 4436 476
rect 4474 448 4502 476
rect 4540 448 4568 476
rect -4568 382 -4540 410
rect -4502 382 -4474 410
rect -4436 382 -4408 410
rect -4370 382 -4342 410
rect -4304 382 -4276 410
rect -4238 382 -4210 410
rect -4172 382 -4144 410
rect -4106 382 -4078 410
rect -4040 382 -4012 410
rect -3974 382 -3946 410
rect -3908 382 -3880 410
rect -3842 382 -3814 410
rect -3776 382 -3748 410
rect -3710 382 -3682 410
rect -3644 382 -3616 410
rect -3578 382 -3550 410
rect -3512 382 -3484 410
rect -3446 382 -3418 410
rect -3380 382 -3352 410
rect -3314 382 -3286 410
rect -3248 382 -3220 410
rect -3182 382 -3154 410
rect -3116 382 -3088 410
rect -3050 382 -3022 410
rect -2984 382 -2956 410
rect -2918 382 -2890 410
rect -2852 382 -2824 410
rect -2786 382 -2758 410
rect -2720 382 -2692 410
rect -2654 382 -2626 410
rect -2588 382 -2560 410
rect -2522 382 -2494 410
rect -2456 382 -2428 410
rect -2390 382 -2362 410
rect -2324 382 -2296 410
rect -2258 382 -2230 410
rect -2192 382 -2164 410
rect -2126 382 -2098 410
rect -2060 382 -2032 410
rect -1994 382 -1966 410
rect -1928 382 -1900 410
rect -1862 382 -1834 410
rect -1796 382 -1768 410
rect -1730 382 -1702 410
rect -1664 382 -1636 410
rect -1598 382 -1570 410
rect -1532 382 -1504 410
rect -1466 382 -1438 410
rect -1400 382 -1372 410
rect -1334 382 -1306 410
rect -1268 382 -1240 410
rect -1202 382 -1174 410
rect -1136 382 -1108 410
rect -1070 382 -1042 410
rect -1004 382 -976 410
rect -938 382 -910 410
rect -872 382 -844 410
rect -806 382 -778 410
rect -740 382 -712 410
rect -674 382 -646 410
rect -608 382 -580 410
rect -542 382 -514 410
rect -476 382 -448 410
rect -410 382 -382 410
rect -344 382 -316 410
rect -278 382 -250 410
rect -212 382 -184 410
rect -146 382 -118 410
rect -80 382 -52 410
rect -14 382 14 410
rect 52 382 80 410
rect 118 382 146 410
rect 184 382 212 410
rect 250 382 278 410
rect 316 382 344 410
rect 382 382 410 410
rect 448 382 476 410
rect 514 382 542 410
rect 580 382 608 410
rect 646 382 674 410
rect 712 382 740 410
rect 778 382 806 410
rect 844 382 872 410
rect 910 382 938 410
rect 976 382 1004 410
rect 1042 382 1070 410
rect 1108 382 1136 410
rect 1174 382 1202 410
rect 1240 382 1268 410
rect 1306 382 1334 410
rect 1372 382 1400 410
rect 1438 382 1466 410
rect 1504 382 1532 410
rect 1570 382 1598 410
rect 1636 382 1664 410
rect 1702 382 1730 410
rect 1768 382 1796 410
rect 1834 382 1862 410
rect 1900 382 1928 410
rect 1966 382 1994 410
rect 2032 382 2060 410
rect 2098 382 2126 410
rect 2164 382 2192 410
rect 2230 382 2258 410
rect 2296 382 2324 410
rect 2362 382 2390 410
rect 2428 382 2456 410
rect 2494 382 2522 410
rect 2560 382 2588 410
rect 2626 382 2654 410
rect 2692 382 2720 410
rect 2758 382 2786 410
rect 2824 382 2852 410
rect 2890 382 2918 410
rect 2956 382 2984 410
rect 3022 382 3050 410
rect 3088 382 3116 410
rect 3154 382 3182 410
rect 3220 382 3248 410
rect 3286 382 3314 410
rect 3352 382 3380 410
rect 3418 382 3446 410
rect 3484 382 3512 410
rect 3550 382 3578 410
rect 3616 382 3644 410
rect 3682 382 3710 410
rect 3748 382 3776 410
rect 3814 382 3842 410
rect 3880 382 3908 410
rect 3946 382 3974 410
rect 4012 382 4040 410
rect 4078 382 4106 410
rect 4144 382 4172 410
rect 4210 382 4238 410
rect 4276 382 4304 410
rect 4342 382 4370 410
rect 4408 382 4436 410
rect 4474 382 4502 410
rect 4540 382 4568 410
rect -4568 316 -4540 344
rect -4502 316 -4474 344
rect -4436 316 -4408 344
rect -4370 316 -4342 344
rect -4304 316 -4276 344
rect -4238 316 -4210 344
rect -4172 316 -4144 344
rect -4106 316 -4078 344
rect -4040 316 -4012 344
rect -3974 316 -3946 344
rect -3908 316 -3880 344
rect -3842 316 -3814 344
rect -3776 316 -3748 344
rect -3710 316 -3682 344
rect -3644 316 -3616 344
rect -3578 316 -3550 344
rect -3512 316 -3484 344
rect -3446 316 -3418 344
rect -3380 316 -3352 344
rect -3314 316 -3286 344
rect -3248 316 -3220 344
rect -3182 316 -3154 344
rect -3116 316 -3088 344
rect -3050 316 -3022 344
rect -2984 316 -2956 344
rect -2918 316 -2890 344
rect -2852 316 -2824 344
rect -2786 316 -2758 344
rect -2720 316 -2692 344
rect -2654 316 -2626 344
rect -2588 316 -2560 344
rect -2522 316 -2494 344
rect -2456 316 -2428 344
rect -2390 316 -2362 344
rect -2324 316 -2296 344
rect -2258 316 -2230 344
rect -2192 316 -2164 344
rect -2126 316 -2098 344
rect -2060 316 -2032 344
rect -1994 316 -1966 344
rect -1928 316 -1900 344
rect -1862 316 -1834 344
rect -1796 316 -1768 344
rect -1730 316 -1702 344
rect -1664 316 -1636 344
rect -1598 316 -1570 344
rect -1532 316 -1504 344
rect -1466 316 -1438 344
rect -1400 316 -1372 344
rect -1334 316 -1306 344
rect -1268 316 -1240 344
rect -1202 316 -1174 344
rect -1136 316 -1108 344
rect -1070 316 -1042 344
rect -1004 316 -976 344
rect -938 316 -910 344
rect -872 316 -844 344
rect -806 316 -778 344
rect -740 316 -712 344
rect -674 316 -646 344
rect -608 316 -580 344
rect -542 316 -514 344
rect -476 316 -448 344
rect -410 316 -382 344
rect -344 316 -316 344
rect -278 316 -250 344
rect -212 316 -184 344
rect -146 316 -118 344
rect -80 316 -52 344
rect -14 316 14 344
rect 52 316 80 344
rect 118 316 146 344
rect 184 316 212 344
rect 250 316 278 344
rect 316 316 344 344
rect 382 316 410 344
rect 448 316 476 344
rect 514 316 542 344
rect 580 316 608 344
rect 646 316 674 344
rect 712 316 740 344
rect 778 316 806 344
rect 844 316 872 344
rect 910 316 938 344
rect 976 316 1004 344
rect 1042 316 1070 344
rect 1108 316 1136 344
rect 1174 316 1202 344
rect 1240 316 1268 344
rect 1306 316 1334 344
rect 1372 316 1400 344
rect 1438 316 1466 344
rect 1504 316 1532 344
rect 1570 316 1598 344
rect 1636 316 1664 344
rect 1702 316 1730 344
rect 1768 316 1796 344
rect 1834 316 1862 344
rect 1900 316 1928 344
rect 1966 316 1994 344
rect 2032 316 2060 344
rect 2098 316 2126 344
rect 2164 316 2192 344
rect 2230 316 2258 344
rect 2296 316 2324 344
rect 2362 316 2390 344
rect 2428 316 2456 344
rect 2494 316 2522 344
rect 2560 316 2588 344
rect 2626 316 2654 344
rect 2692 316 2720 344
rect 2758 316 2786 344
rect 2824 316 2852 344
rect 2890 316 2918 344
rect 2956 316 2984 344
rect 3022 316 3050 344
rect 3088 316 3116 344
rect 3154 316 3182 344
rect 3220 316 3248 344
rect 3286 316 3314 344
rect 3352 316 3380 344
rect 3418 316 3446 344
rect 3484 316 3512 344
rect 3550 316 3578 344
rect 3616 316 3644 344
rect 3682 316 3710 344
rect 3748 316 3776 344
rect 3814 316 3842 344
rect 3880 316 3908 344
rect 3946 316 3974 344
rect 4012 316 4040 344
rect 4078 316 4106 344
rect 4144 316 4172 344
rect 4210 316 4238 344
rect 4276 316 4304 344
rect 4342 316 4370 344
rect 4408 316 4436 344
rect 4474 316 4502 344
rect 4540 316 4568 344
rect -4568 250 -4540 278
rect -4502 250 -4474 278
rect -4436 250 -4408 278
rect -4370 250 -4342 278
rect -4304 250 -4276 278
rect -4238 250 -4210 278
rect -4172 250 -4144 278
rect -4106 250 -4078 278
rect -4040 250 -4012 278
rect -3974 250 -3946 278
rect -3908 250 -3880 278
rect -3842 250 -3814 278
rect -3776 250 -3748 278
rect -3710 250 -3682 278
rect -3644 250 -3616 278
rect -3578 250 -3550 278
rect -3512 250 -3484 278
rect -3446 250 -3418 278
rect -3380 250 -3352 278
rect -3314 250 -3286 278
rect -3248 250 -3220 278
rect -3182 250 -3154 278
rect -3116 250 -3088 278
rect -3050 250 -3022 278
rect -2984 250 -2956 278
rect -2918 250 -2890 278
rect -2852 250 -2824 278
rect -2786 250 -2758 278
rect -2720 250 -2692 278
rect -2654 250 -2626 278
rect -2588 250 -2560 278
rect -2522 250 -2494 278
rect -2456 250 -2428 278
rect -2390 250 -2362 278
rect -2324 250 -2296 278
rect -2258 250 -2230 278
rect -2192 250 -2164 278
rect -2126 250 -2098 278
rect -2060 250 -2032 278
rect -1994 250 -1966 278
rect -1928 250 -1900 278
rect -1862 250 -1834 278
rect -1796 250 -1768 278
rect -1730 250 -1702 278
rect -1664 250 -1636 278
rect -1598 250 -1570 278
rect -1532 250 -1504 278
rect -1466 250 -1438 278
rect -1400 250 -1372 278
rect -1334 250 -1306 278
rect -1268 250 -1240 278
rect -1202 250 -1174 278
rect -1136 250 -1108 278
rect -1070 250 -1042 278
rect -1004 250 -976 278
rect -938 250 -910 278
rect -872 250 -844 278
rect -806 250 -778 278
rect -740 250 -712 278
rect -674 250 -646 278
rect -608 250 -580 278
rect -542 250 -514 278
rect -476 250 -448 278
rect -410 250 -382 278
rect -344 250 -316 278
rect -278 250 -250 278
rect -212 250 -184 278
rect -146 250 -118 278
rect -80 250 -52 278
rect -14 250 14 278
rect 52 250 80 278
rect 118 250 146 278
rect 184 250 212 278
rect 250 250 278 278
rect 316 250 344 278
rect 382 250 410 278
rect 448 250 476 278
rect 514 250 542 278
rect 580 250 608 278
rect 646 250 674 278
rect 712 250 740 278
rect 778 250 806 278
rect 844 250 872 278
rect 910 250 938 278
rect 976 250 1004 278
rect 1042 250 1070 278
rect 1108 250 1136 278
rect 1174 250 1202 278
rect 1240 250 1268 278
rect 1306 250 1334 278
rect 1372 250 1400 278
rect 1438 250 1466 278
rect 1504 250 1532 278
rect 1570 250 1598 278
rect 1636 250 1664 278
rect 1702 250 1730 278
rect 1768 250 1796 278
rect 1834 250 1862 278
rect 1900 250 1928 278
rect 1966 250 1994 278
rect 2032 250 2060 278
rect 2098 250 2126 278
rect 2164 250 2192 278
rect 2230 250 2258 278
rect 2296 250 2324 278
rect 2362 250 2390 278
rect 2428 250 2456 278
rect 2494 250 2522 278
rect 2560 250 2588 278
rect 2626 250 2654 278
rect 2692 250 2720 278
rect 2758 250 2786 278
rect 2824 250 2852 278
rect 2890 250 2918 278
rect 2956 250 2984 278
rect 3022 250 3050 278
rect 3088 250 3116 278
rect 3154 250 3182 278
rect 3220 250 3248 278
rect 3286 250 3314 278
rect 3352 250 3380 278
rect 3418 250 3446 278
rect 3484 250 3512 278
rect 3550 250 3578 278
rect 3616 250 3644 278
rect 3682 250 3710 278
rect 3748 250 3776 278
rect 3814 250 3842 278
rect 3880 250 3908 278
rect 3946 250 3974 278
rect 4012 250 4040 278
rect 4078 250 4106 278
rect 4144 250 4172 278
rect 4210 250 4238 278
rect 4276 250 4304 278
rect 4342 250 4370 278
rect 4408 250 4436 278
rect 4474 250 4502 278
rect 4540 250 4568 278
rect -4568 184 -4540 212
rect -4502 184 -4474 212
rect -4436 184 -4408 212
rect -4370 184 -4342 212
rect -4304 184 -4276 212
rect -4238 184 -4210 212
rect -4172 184 -4144 212
rect -4106 184 -4078 212
rect -4040 184 -4012 212
rect -3974 184 -3946 212
rect -3908 184 -3880 212
rect -3842 184 -3814 212
rect -3776 184 -3748 212
rect -3710 184 -3682 212
rect -3644 184 -3616 212
rect -3578 184 -3550 212
rect -3512 184 -3484 212
rect -3446 184 -3418 212
rect -3380 184 -3352 212
rect -3314 184 -3286 212
rect -3248 184 -3220 212
rect -3182 184 -3154 212
rect -3116 184 -3088 212
rect -3050 184 -3022 212
rect -2984 184 -2956 212
rect -2918 184 -2890 212
rect -2852 184 -2824 212
rect -2786 184 -2758 212
rect -2720 184 -2692 212
rect -2654 184 -2626 212
rect -2588 184 -2560 212
rect -2522 184 -2494 212
rect -2456 184 -2428 212
rect -2390 184 -2362 212
rect -2324 184 -2296 212
rect -2258 184 -2230 212
rect -2192 184 -2164 212
rect -2126 184 -2098 212
rect -2060 184 -2032 212
rect -1994 184 -1966 212
rect -1928 184 -1900 212
rect -1862 184 -1834 212
rect -1796 184 -1768 212
rect -1730 184 -1702 212
rect -1664 184 -1636 212
rect -1598 184 -1570 212
rect -1532 184 -1504 212
rect -1466 184 -1438 212
rect -1400 184 -1372 212
rect -1334 184 -1306 212
rect -1268 184 -1240 212
rect -1202 184 -1174 212
rect -1136 184 -1108 212
rect -1070 184 -1042 212
rect -1004 184 -976 212
rect -938 184 -910 212
rect -872 184 -844 212
rect -806 184 -778 212
rect -740 184 -712 212
rect -674 184 -646 212
rect -608 184 -580 212
rect -542 184 -514 212
rect -476 184 -448 212
rect -410 184 -382 212
rect -344 184 -316 212
rect -278 184 -250 212
rect -212 184 -184 212
rect -146 184 -118 212
rect -80 184 -52 212
rect -14 184 14 212
rect 52 184 80 212
rect 118 184 146 212
rect 184 184 212 212
rect 250 184 278 212
rect 316 184 344 212
rect 382 184 410 212
rect 448 184 476 212
rect 514 184 542 212
rect 580 184 608 212
rect 646 184 674 212
rect 712 184 740 212
rect 778 184 806 212
rect 844 184 872 212
rect 910 184 938 212
rect 976 184 1004 212
rect 1042 184 1070 212
rect 1108 184 1136 212
rect 1174 184 1202 212
rect 1240 184 1268 212
rect 1306 184 1334 212
rect 1372 184 1400 212
rect 1438 184 1466 212
rect 1504 184 1532 212
rect 1570 184 1598 212
rect 1636 184 1664 212
rect 1702 184 1730 212
rect 1768 184 1796 212
rect 1834 184 1862 212
rect 1900 184 1928 212
rect 1966 184 1994 212
rect 2032 184 2060 212
rect 2098 184 2126 212
rect 2164 184 2192 212
rect 2230 184 2258 212
rect 2296 184 2324 212
rect 2362 184 2390 212
rect 2428 184 2456 212
rect 2494 184 2522 212
rect 2560 184 2588 212
rect 2626 184 2654 212
rect 2692 184 2720 212
rect 2758 184 2786 212
rect 2824 184 2852 212
rect 2890 184 2918 212
rect 2956 184 2984 212
rect 3022 184 3050 212
rect 3088 184 3116 212
rect 3154 184 3182 212
rect 3220 184 3248 212
rect 3286 184 3314 212
rect 3352 184 3380 212
rect 3418 184 3446 212
rect 3484 184 3512 212
rect 3550 184 3578 212
rect 3616 184 3644 212
rect 3682 184 3710 212
rect 3748 184 3776 212
rect 3814 184 3842 212
rect 3880 184 3908 212
rect 3946 184 3974 212
rect 4012 184 4040 212
rect 4078 184 4106 212
rect 4144 184 4172 212
rect 4210 184 4238 212
rect 4276 184 4304 212
rect 4342 184 4370 212
rect 4408 184 4436 212
rect 4474 184 4502 212
rect 4540 184 4568 212
rect -4568 118 -4540 146
rect -4502 118 -4474 146
rect -4436 118 -4408 146
rect -4370 118 -4342 146
rect -4304 118 -4276 146
rect -4238 118 -4210 146
rect -4172 118 -4144 146
rect -4106 118 -4078 146
rect -4040 118 -4012 146
rect -3974 118 -3946 146
rect -3908 118 -3880 146
rect -3842 118 -3814 146
rect -3776 118 -3748 146
rect -3710 118 -3682 146
rect -3644 118 -3616 146
rect -3578 118 -3550 146
rect -3512 118 -3484 146
rect -3446 118 -3418 146
rect -3380 118 -3352 146
rect -3314 118 -3286 146
rect -3248 118 -3220 146
rect -3182 118 -3154 146
rect -3116 118 -3088 146
rect -3050 118 -3022 146
rect -2984 118 -2956 146
rect -2918 118 -2890 146
rect -2852 118 -2824 146
rect -2786 118 -2758 146
rect -2720 118 -2692 146
rect -2654 118 -2626 146
rect -2588 118 -2560 146
rect -2522 118 -2494 146
rect -2456 118 -2428 146
rect -2390 118 -2362 146
rect -2324 118 -2296 146
rect -2258 118 -2230 146
rect -2192 118 -2164 146
rect -2126 118 -2098 146
rect -2060 118 -2032 146
rect -1994 118 -1966 146
rect -1928 118 -1900 146
rect -1862 118 -1834 146
rect -1796 118 -1768 146
rect -1730 118 -1702 146
rect -1664 118 -1636 146
rect -1598 118 -1570 146
rect -1532 118 -1504 146
rect -1466 118 -1438 146
rect -1400 118 -1372 146
rect -1334 118 -1306 146
rect -1268 118 -1240 146
rect -1202 118 -1174 146
rect -1136 118 -1108 146
rect -1070 118 -1042 146
rect -1004 118 -976 146
rect -938 118 -910 146
rect -872 118 -844 146
rect -806 118 -778 146
rect -740 118 -712 146
rect -674 118 -646 146
rect -608 118 -580 146
rect -542 118 -514 146
rect -476 118 -448 146
rect -410 118 -382 146
rect -344 118 -316 146
rect -278 118 -250 146
rect -212 118 -184 146
rect -146 118 -118 146
rect -80 118 -52 146
rect -14 118 14 146
rect 52 118 80 146
rect 118 118 146 146
rect 184 118 212 146
rect 250 118 278 146
rect 316 118 344 146
rect 382 118 410 146
rect 448 118 476 146
rect 514 118 542 146
rect 580 118 608 146
rect 646 118 674 146
rect 712 118 740 146
rect 778 118 806 146
rect 844 118 872 146
rect 910 118 938 146
rect 976 118 1004 146
rect 1042 118 1070 146
rect 1108 118 1136 146
rect 1174 118 1202 146
rect 1240 118 1268 146
rect 1306 118 1334 146
rect 1372 118 1400 146
rect 1438 118 1466 146
rect 1504 118 1532 146
rect 1570 118 1598 146
rect 1636 118 1664 146
rect 1702 118 1730 146
rect 1768 118 1796 146
rect 1834 118 1862 146
rect 1900 118 1928 146
rect 1966 118 1994 146
rect 2032 118 2060 146
rect 2098 118 2126 146
rect 2164 118 2192 146
rect 2230 118 2258 146
rect 2296 118 2324 146
rect 2362 118 2390 146
rect 2428 118 2456 146
rect 2494 118 2522 146
rect 2560 118 2588 146
rect 2626 118 2654 146
rect 2692 118 2720 146
rect 2758 118 2786 146
rect 2824 118 2852 146
rect 2890 118 2918 146
rect 2956 118 2984 146
rect 3022 118 3050 146
rect 3088 118 3116 146
rect 3154 118 3182 146
rect 3220 118 3248 146
rect 3286 118 3314 146
rect 3352 118 3380 146
rect 3418 118 3446 146
rect 3484 118 3512 146
rect 3550 118 3578 146
rect 3616 118 3644 146
rect 3682 118 3710 146
rect 3748 118 3776 146
rect 3814 118 3842 146
rect 3880 118 3908 146
rect 3946 118 3974 146
rect 4012 118 4040 146
rect 4078 118 4106 146
rect 4144 118 4172 146
rect 4210 118 4238 146
rect 4276 118 4304 146
rect 4342 118 4370 146
rect 4408 118 4436 146
rect 4474 118 4502 146
rect 4540 118 4568 146
rect -4568 52 -4540 80
rect -4502 52 -4474 80
rect -4436 52 -4408 80
rect -4370 52 -4342 80
rect -4304 52 -4276 80
rect -4238 52 -4210 80
rect -4172 52 -4144 80
rect -4106 52 -4078 80
rect -4040 52 -4012 80
rect -3974 52 -3946 80
rect -3908 52 -3880 80
rect -3842 52 -3814 80
rect -3776 52 -3748 80
rect -3710 52 -3682 80
rect -3644 52 -3616 80
rect -3578 52 -3550 80
rect -3512 52 -3484 80
rect -3446 52 -3418 80
rect -3380 52 -3352 80
rect -3314 52 -3286 80
rect -3248 52 -3220 80
rect -3182 52 -3154 80
rect -3116 52 -3088 80
rect -3050 52 -3022 80
rect -2984 52 -2956 80
rect -2918 52 -2890 80
rect -2852 52 -2824 80
rect -2786 52 -2758 80
rect -2720 52 -2692 80
rect -2654 52 -2626 80
rect -2588 52 -2560 80
rect -2522 52 -2494 80
rect -2456 52 -2428 80
rect -2390 52 -2362 80
rect -2324 52 -2296 80
rect -2258 52 -2230 80
rect -2192 52 -2164 80
rect -2126 52 -2098 80
rect -2060 52 -2032 80
rect -1994 52 -1966 80
rect -1928 52 -1900 80
rect -1862 52 -1834 80
rect -1796 52 -1768 80
rect -1730 52 -1702 80
rect -1664 52 -1636 80
rect -1598 52 -1570 80
rect -1532 52 -1504 80
rect -1466 52 -1438 80
rect -1400 52 -1372 80
rect -1334 52 -1306 80
rect -1268 52 -1240 80
rect -1202 52 -1174 80
rect -1136 52 -1108 80
rect -1070 52 -1042 80
rect -1004 52 -976 80
rect -938 52 -910 80
rect -872 52 -844 80
rect -806 52 -778 80
rect -740 52 -712 80
rect -674 52 -646 80
rect -608 52 -580 80
rect -542 52 -514 80
rect -476 52 -448 80
rect -410 52 -382 80
rect -344 52 -316 80
rect -278 52 -250 80
rect -212 52 -184 80
rect -146 52 -118 80
rect -80 52 -52 80
rect -14 52 14 80
rect 52 52 80 80
rect 118 52 146 80
rect 184 52 212 80
rect 250 52 278 80
rect 316 52 344 80
rect 382 52 410 80
rect 448 52 476 80
rect 514 52 542 80
rect 580 52 608 80
rect 646 52 674 80
rect 712 52 740 80
rect 778 52 806 80
rect 844 52 872 80
rect 910 52 938 80
rect 976 52 1004 80
rect 1042 52 1070 80
rect 1108 52 1136 80
rect 1174 52 1202 80
rect 1240 52 1268 80
rect 1306 52 1334 80
rect 1372 52 1400 80
rect 1438 52 1466 80
rect 1504 52 1532 80
rect 1570 52 1598 80
rect 1636 52 1664 80
rect 1702 52 1730 80
rect 1768 52 1796 80
rect 1834 52 1862 80
rect 1900 52 1928 80
rect 1966 52 1994 80
rect 2032 52 2060 80
rect 2098 52 2126 80
rect 2164 52 2192 80
rect 2230 52 2258 80
rect 2296 52 2324 80
rect 2362 52 2390 80
rect 2428 52 2456 80
rect 2494 52 2522 80
rect 2560 52 2588 80
rect 2626 52 2654 80
rect 2692 52 2720 80
rect 2758 52 2786 80
rect 2824 52 2852 80
rect 2890 52 2918 80
rect 2956 52 2984 80
rect 3022 52 3050 80
rect 3088 52 3116 80
rect 3154 52 3182 80
rect 3220 52 3248 80
rect 3286 52 3314 80
rect 3352 52 3380 80
rect 3418 52 3446 80
rect 3484 52 3512 80
rect 3550 52 3578 80
rect 3616 52 3644 80
rect 3682 52 3710 80
rect 3748 52 3776 80
rect 3814 52 3842 80
rect 3880 52 3908 80
rect 3946 52 3974 80
rect 4012 52 4040 80
rect 4078 52 4106 80
rect 4144 52 4172 80
rect 4210 52 4238 80
rect 4276 52 4304 80
rect 4342 52 4370 80
rect 4408 52 4436 80
rect 4474 52 4502 80
rect 4540 52 4568 80
rect -4568 -14 -4540 14
rect -4502 -14 -4474 14
rect -4436 -14 -4408 14
rect -4370 -14 -4342 14
rect -4304 -14 -4276 14
rect -4238 -14 -4210 14
rect -4172 -14 -4144 14
rect -4106 -14 -4078 14
rect -4040 -14 -4012 14
rect -3974 -14 -3946 14
rect -3908 -14 -3880 14
rect -3842 -14 -3814 14
rect -3776 -14 -3748 14
rect -3710 -14 -3682 14
rect -3644 -14 -3616 14
rect -3578 -14 -3550 14
rect -3512 -14 -3484 14
rect -3446 -14 -3418 14
rect -3380 -14 -3352 14
rect -3314 -14 -3286 14
rect -3248 -14 -3220 14
rect -3182 -14 -3154 14
rect -3116 -14 -3088 14
rect -3050 -14 -3022 14
rect -2984 -14 -2956 14
rect -2918 -14 -2890 14
rect -2852 -14 -2824 14
rect -2786 -14 -2758 14
rect -2720 -14 -2692 14
rect -2654 -14 -2626 14
rect -2588 -14 -2560 14
rect -2522 -14 -2494 14
rect -2456 -14 -2428 14
rect -2390 -14 -2362 14
rect -2324 -14 -2296 14
rect -2258 -14 -2230 14
rect -2192 -14 -2164 14
rect -2126 -14 -2098 14
rect -2060 -14 -2032 14
rect -1994 -14 -1966 14
rect -1928 -14 -1900 14
rect -1862 -14 -1834 14
rect -1796 -14 -1768 14
rect -1730 -14 -1702 14
rect -1664 -14 -1636 14
rect -1598 -14 -1570 14
rect -1532 -14 -1504 14
rect -1466 -14 -1438 14
rect -1400 -14 -1372 14
rect -1334 -14 -1306 14
rect -1268 -14 -1240 14
rect -1202 -14 -1174 14
rect -1136 -14 -1108 14
rect -1070 -14 -1042 14
rect -1004 -14 -976 14
rect -938 -14 -910 14
rect -872 -14 -844 14
rect -806 -14 -778 14
rect -740 -14 -712 14
rect -674 -14 -646 14
rect -608 -14 -580 14
rect -542 -14 -514 14
rect -476 -14 -448 14
rect -410 -14 -382 14
rect -344 -14 -316 14
rect -278 -14 -250 14
rect -212 -14 -184 14
rect -146 -14 -118 14
rect -80 -14 -52 14
rect -14 -14 14 14
rect 52 -14 80 14
rect 118 -14 146 14
rect 184 -14 212 14
rect 250 -14 278 14
rect 316 -14 344 14
rect 382 -14 410 14
rect 448 -14 476 14
rect 514 -14 542 14
rect 580 -14 608 14
rect 646 -14 674 14
rect 712 -14 740 14
rect 778 -14 806 14
rect 844 -14 872 14
rect 910 -14 938 14
rect 976 -14 1004 14
rect 1042 -14 1070 14
rect 1108 -14 1136 14
rect 1174 -14 1202 14
rect 1240 -14 1268 14
rect 1306 -14 1334 14
rect 1372 -14 1400 14
rect 1438 -14 1466 14
rect 1504 -14 1532 14
rect 1570 -14 1598 14
rect 1636 -14 1664 14
rect 1702 -14 1730 14
rect 1768 -14 1796 14
rect 1834 -14 1862 14
rect 1900 -14 1928 14
rect 1966 -14 1994 14
rect 2032 -14 2060 14
rect 2098 -14 2126 14
rect 2164 -14 2192 14
rect 2230 -14 2258 14
rect 2296 -14 2324 14
rect 2362 -14 2390 14
rect 2428 -14 2456 14
rect 2494 -14 2522 14
rect 2560 -14 2588 14
rect 2626 -14 2654 14
rect 2692 -14 2720 14
rect 2758 -14 2786 14
rect 2824 -14 2852 14
rect 2890 -14 2918 14
rect 2956 -14 2984 14
rect 3022 -14 3050 14
rect 3088 -14 3116 14
rect 3154 -14 3182 14
rect 3220 -14 3248 14
rect 3286 -14 3314 14
rect 3352 -14 3380 14
rect 3418 -14 3446 14
rect 3484 -14 3512 14
rect 3550 -14 3578 14
rect 3616 -14 3644 14
rect 3682 -14 3710 14
rect 3748 -14 3776 14
rect 3814 -14 3842 14
rect 3880 -14 3908 14
rect 3946 -14 3974 14
rect 4012 -14 4040 14
rect 4078 -14 4106 14
rect 4144 -14 4172 14
rect 4210 -14 4238 14
rect 4276 -14 4304 14
rect 4342 -14 4370 14
rect 4408 -14 4436 14
rect 4474 -14 4502 14
rect 4540 -14 4568 14
rect -4568 -80 -4540 -52
rect -4502 -80 -4474 -52
rect -4436 -80 -4408 -52
rect -4370 -80 -4342 -52
rect -4304 -80 -4276 -52
rect -4238 -80 -4210 -52
rect -4172 -80 -4144 -52
rect -4106 -80 -4078 -52
rect -4040 -80 -4012 -52
rect -3974 -80 -3946 -52
rect -3908 -80 -3880 -52
rect -3842 -80 -3814 -52
rect -3776 -80 -3748 -52
rect -3710 -80 -3682 -52
rect -3644 -80 -3616 -52
rect -3578 -80 -3550 -52
rect -3512 -80 -3484 -52
rect -3446 -80 -3418 -52
rect -3380 -80 -3352 -52
rect -3314 -80 -3286 -52
rect -3248 -80 -3220 -52
rect -3182 -80 -3154 -52
rect -3116 -80 -3088 -52
rect -3050 -80 -3022 -52
rect -2984 -80 -2956 -52
rect -2918 -80 -2890 -52
rect -2852 -80 -2824 -52
rect -2786 -80 -2758 -52
rect -2720 -80 -2692 -52
rect -2654 -80 -2626 -52
rect -2588 -80 -2560 -52
rect -2522 -80 -2494 -52
rect -2456 -80 -2428 -52
rect -2390 -80 -2362 -52
rect -2324 -80 -2296 -52
rect -2258 -80 -2230 -52
rect -2192 -80 -2164 -52
rect -2126 -80 -2098 -52
rect -2060 -80 -2032 -52
rect -1994 -80 -1966 -52
rect -1928 -80 -1900 -52
rect -1862 -80 -1834 -52
rect -1796 -80 -1768 -52
rect -1730 -80 -1702 -52
rect -1664 -80 -1636 -52
rect -1598 -80 -1570 -52
rect -1532 -80 -1504 -52
rect -1466 -80 -1438 -52
rect -1400 -80 -1372 -52
rect -1334 -80 -1306 -52
rect -1268 -80 -1240 -52
rect -1202 -80 -1174 -52
rect -1136 -80 -1108 -52
rect -1070 -80 -1042 -52
rect -1004 -80 -976 -52
rect -938 -80 -910 -52
rect -872 -80 -844 -52
rect -806 -80 -778 -52
rect -740 -80 -712 -52
rect -674 -80 -646 -52
rect -608 -80 -580 -52
rect -542 -80 -514 -52
rect -476 -80 -448 -52
rect -410 -80 -382 -52
rect -344 -80 -316 -52
rect -278 -80 -250 -52
rect -212 -80 -184 -52
rect -146 -80 -118 -52
rect -80 -80 -52 -52
rect -14 -80 14 -52
rect 52 -80 80 -52
rect 118 -80 146 -52
rect 184 -80 212 -52
rect 250 -80 278 -52
rect 316 -80 344 -52
rect 382 -80 410 -52
rect 448 -80 476 -52
rect 514 -80 542 -52
rect 580 -80 608 -52
rect 646 -80 674 -52
rect 712 -80 740 -52
rect 778 -80 806 -52
rect 844 -80 872 -52
rect 910 -80 938 -52
rect 976 -80 1004 -52
rect 1042 -80 1070 -52
rect 1108 -80 1136 -52
rect 1174 -80 1202 -52
rect 1240 -80 1268 -52
rect 1306 -80 1334 -52
rect 1372 -80 1400 -52
rect 1438 -80 1466 -52
rect 1504 -80 1532 -52
rect 1570 -80 1598 -52
rect 1636 -80 1664 -52
rect 1702 -80 1730 -52
rect 1768 -80 1796 -52
rect 1834 -80 1862 -52
rect 1900 -80 1928 -52
rect 1966 -80 1994 -52
rect 2032 -80 2060 -52
rect 2098 -80 2126 -52
rect 2164 -80 2192 -52
rect 2230 -80 2258 -52
rect 2296 -80 2324 -52
rect 2362 -80 2390 -52
rect 2428 -80 2456 -52
rect 2494 -80 2522 -52
rect 2560 -80 2588 -52
rect 2626 -80 2654 -52
rect 2692 -80 2720 -52
rect 2758 -80 2786 -52
rect 2824 -80 2852 -52
rect 2890 -80 2918 -52
rect 2956 -80 2984 -52
rect 3022 -80 3050 -52
rect 3088 -80 3116 -52
rect 3154 -80 3182 -52
rect 3220 -80 3248 -52
rect 3286 -80 3314 -52
rect 3352 -80 3380 -52
rect 3418 -80 3446 -52
rect 3484 -80 3512 -52
rect 3550 -80 3578 -52
rect 3616 -80 3644 -52
rect 3682 -80 3710 -52
rect 3748 -80 3776 -52
rect 3814 -80 3842 -52
rect 3880 -80 3908 -52
rect 3946 -80 3974 -52
rect 4012 -80 4040 -52
rect 4078 -80 4106 -52
rect 4144 -80 4172 -52
rect 4210 -80 4238 -52
rect 4276 -80 4304 -52
rect 4342 -80 4370 -52
rect 4408 -80 4436 -52
rect 4474 -80 4502 -52
rect 4540 -80 4568 -52
rect -4568 -146 -4540 -118
rect -4502 -146 -4474 -118
rect -4436 -146 -4408 -118
rect -4370 -146 -4342 -118
rect -4304 -146 -4276 -118
rect -4238 -146 -4210 -118
rect -4172 -146 -4144 -118
rect -4106 -146 -4078 -118
rect -4040 -146 -4012 -118
rect -3974 -146 -3946 -118
rect -3908 -146 -3880 -118
rect -3842 -146 -3814 -118
rect -3776 -146 -3748 -118
rect -3710 -146 -3682 -118
rect -3644 -146 -3616 -118
rect -3578 -146 -3550 -118
rect -3512 -146 -3484 -118
rect -3446 -146 -3418 -118
rect -3380 -146 -3352 -118
rect -3314 -146 -3286 -118
rect -3248 -146 -3220 -118
rect -3182 -146 -3154 -118
rect -3116 -146 -3088 -118
rect -3050 -146 -3022 -118
rect -2984 -146 -2956 -118
rect -2918 -146 -2890 -118
rect -2852 -146 -2824 -118
rect -2786 -146 -2758 -118
rect -2720 -146 -2692 -118
rect -2654 -146 -2626 -118
rect -2588 -146 -2560 -118
rect -2522 -146 -2494 -118
rect -2456 -146 -2428 -118
rect -2390 -146 -2362 -118
rect -2324 -146 -2296 -118
rect -2258 -146 -2230 -118
rect -2192 -146 -2164 -118
rect -2126 -146 -2098 -118
rect -2060 -146 -2032 -118
rect -1994 -146 -1966 -118
rect -1928 -146 -1900 -118
rect -1862 -146 -1834 -118
rect -1796 -146 -1768 -118
rect -1730 -146 -1702 -118
rect -1664 -146 -1636 -118
rect -1598 -146 -1570 -118
rect -1532 -146 -1504 -118
rect -1466 -146 -1438 -118
rect -1400 -146 -1372 -118
rect -1334 -146 -1306 -118
rect -1268 -146 -1240 -118
rect -1202 -146 -1174 -118
rect -1136 -146 -1108 -118
rect -1070 -146 -1042 -118
rect -1004 -146 -976 -118
rect -938 -146 -910 -118
rect -872 -146 -844 -118
rect -806 -146 -778 -118
rect -740 -146 -712 -118
rect -674 -146 -646 -118
rect -608 -146 -580 -118
rect -542 -146 -514 -118
rect -476 -146 -448 -118
rect -410 -146 -382 -118
rect -344 -146 -316 -118
rect -278 -146 -250 -118
rect -212 -146 -184 -118
rect -146 -146 -118 -118
rect -80 -146 -52 -118
rect -14 -146 14 -118
rect 52 -146 80 -118
rect 118 -146 146 -118
rect 184 -146 212 -118
rect 250 -146 278 -118
rect 316 -146 344 -118
rect 382 -146 410 -118
rect 448 -146 476 -118
rect 514 -146 542 -118
rect 580 -146 608 -118
rect 646 -146 674 -118
rect 712 -146 740 -118
rect 778 -146 806 -118
rect 844 -146 872 -118
rect 910 -146 938 -118
rect 976 -146 1004 -118
rect 1042 -146 1070 -118
rect 1108 -146 1136 -118
rect 1174 -146 1202 -118
rect 1240 -146 1268 -118
rect 1306 -146 1334 -118
rect 1372 -146 1400 -118
rect 1438 -146 1466 -118
rect 1504 -146 1532 -118
rect 1570 -146 1598 -118
rect 1636 -146 1664 -118
rect 1702 -146 1730 -118
rect 1768 -146 1796 -118
rect 1834 -146 1862 -118
rect 1900 -146 1928 -118
rect 1966 -146 1994 -118
rect 2032 -146 2060 -118
rect 2098 -146 2126 -118
rect 2164 -146 2192 -118
rect 2230 -146 2258 -118
rect 2296 -146 2324 -118
rect 2362 -146 2390 -118
rect 2428 -146 2456 -118
rect 2494 -146 2522 -118
rect 2560 -146 2588 -118
rect 2626 -146 2654 -118
rect 2692 -146 2720 -118
rect 2758 -146 2786 -118
rect 2824 -146 2852 -118
rect 2890 -146 2918 -118
rect 2956 -146 2984 -118
rect 3022 -146 3050 -118
rect 3088 -146 3116 -118
rect 3154 -146 3182 -118
rect 3220 -146 3248 -118
rect 3286 -146 3314 -118
rect 3352 -146 3380 -118
rect 3418 -146 3446 -118
rect 3484 -146 3512 -118
rect 3550 -146 3578 -118
rect 3616 -146 3644 -118
rect 3682 -146 3710 -118
rect 3748 -146 3776 -118
rect 3814 -146 3842 -118
rect 3880 -146 3908 -118
rect 3946 -146 3974 -118
rect 4012 -146 4040 -118
rect 4078 -146 4106 -118
rect 4144 -146 4172 -118
rect 4210 -146 4238 -118
rect 4276 -146 4304 -118
rect 4342 -146 4370 -118
rect 4408 -146 4436 -118
rect 4474 -146 4502 -118
rect 4540 -146 4568 -118
rect -4568 -212 -4540 -184
rect -4502 -212 -4474 -184
rect -4436 -212 -4408 -184
rect -4370 -212 -4342 -184
rect -4304 -212 -4276 -184
rect -4238 -212 -4210 -184
rect -4172 -212 -4144 -184
rect -4106 -212 -4078 -184
rect -4040 -212 -4012 -184
rect -3974 -212 -3946 -184
rect -3908 -212 -3880 -184
rect -3842 -212 -3814 -184
rect -3776 -212 -3748 -184
rect -3710 -212 -3682 -184
rect -3644 -212 -3616 -184
rect -3578 -212 -3550 -184
rect -3512 -212 -3484 -184
rect -3446 -212 -3418 -184
rect -3380 -212 -3352 -184
rect -3314 -212 -3286 -184
rect -3248 -212 -3220 -184
rect -3182 -212 -3154 -184
rect -3116 -212 -3088 -184
rect -3050 -212 -3022 -184
rect -2984 -212 -2956 -184
rect -2918 -212 -2890 -184
rect -2852 -212 -2824 -184
rect -2786 -212 -2758 -184
rect -2720 -212 -2692 -184
rect -2654 -212 -2626 -184
rect -2588 -212 -2560 -184
rect -2522 -212 -2494 -184
rect -2456 -212 -2428 -184
rect -2390 -212 -2362 -184
rect -2324 -212 -2296 -184
rect -2258 -212 -2230 -184
rect -2192 -212 -2164 -184
rect -2126 -212 -2098 -184
rect -2060 -212 -2032 -184
rect -1994 -212 -1966 -184
rect -1928 -212 -1900 -184
rect -1862 -212 -1834 -184
rect -1796 -212 -1768 -184
rect -1730 -212 -1702 -184
rect -1664 -212 -1636 -184
rect -1598 -212 -1570 -184
rect -1532 -212 -1504 -184
rect -1466 -212 -1438 -184
rect -1400 -212 -1372 -184
rect -1334 -212 -1306 -184
rect -1268 -212 -1240 -184
rect -1202 -212 -1174 -184
rect -1136 -212 -1108 -184
rect -1070 -212 -1042 -184
rect -1004 -212 -976 -184
rect -938 -212 -910 -184
rect -872 -212 -844 -184
rect -806 -212 -778 -184
rect -740 -212 -712 -184
rect -674 -212 -646 -184
rect -608 -212 -580 -184
rect -542 -212 -514 -184
rect -476 -212 -448 -184
rect -410 -212 -382 -184
rect -344 -212 -316 -184
rect -278 -212 -250 -184
rect -212 -212 -184 -184
rect -146 -212 -118 -184
rect -80 -212 -52 -184
rect -14 -212 14 -184
rect 52 -212 80 -184
rect 118 -212 146 -184
rect 184 -212 212 -184
rect 250 -212 278 -184
rect 316 -212 344 -184
rect 382 -212 410 -184
rect 448 -212 476 -184
rect 514 -212 542 -184
rect 580 -212 608 -184
rect 646 -212 674 -184
rect 712 -212 740 -184
rect 778 -212 806 -184
rect 844 -212 872 -184
rect 910 -212 938 -184
rect 976 -212 1004 -184
rect 1042 -212 1070 -184
rect 1108 -212 1136 -184
rect 1174 -212 1202 -184
rect 1240 -212 1268 -184
rect 1306 -212 1334 -184
rect 1372 -212 1400 -184
rect 1438 -212 1466 -184
rect 1504 -212 1532 -184
rect 1570 -212 1598 -184
rect 1636 -212 1664 -184
rect 1702 -212 1730 -184
rect 1768 -212 1796 -184
rect 1834 -212 1862 -184
rect 1900 -212 1928 -184
rect 1966 -212 1994 -184
rect 2032 -212 2060 -184
rect 2098 -212 2126 -184
rect 2164 -212 2192 -184
rect 2230 -212 2258 -184
rect 2296 -212 2324 -184
rect 2362 -212 2390 -184
rect 2428 -212 2456 -184
rect 2494 -212 2522 -184
rect 2560 -212 2588 -184
rect 2626 -212 2654 -184
rect 2692 -212 2720 -184
rect 2758 -212 2786 -184
rect 2824 -212 2852 -184
rect 2890 -212 2918 -184
rect 2956 -212 2984 -184
rect 3022 -212 3050 -184
rect 3088 -212 3116 -184
rect 3154 -212 3182 -184
rect 3220 -212 3248 -184
rect 3286 -212 3314 -184
rect 3352 -212 3380 -184
rect 3418 -212 3446 -184
rect 3484 -212 3512 -184
rect 3550 -212 3578 -184
rect 3616 -212 3644 -184
rect 3682 -212 3710 -184
rect 3748 -212 3776 -184
rect 3814 -212 3842 -184
rect 3880 -212 3908 -184
rect 3946 -212 3974 -184
rect 4012 -212 4040 -184
rect 4078 -212 4106 -184
rect 4144 -212 4172 -184
rect 4210 -212 4238 -184
rect 4276 -212 4304 -184
rect 4342 -212 4370 -184
rect 4408 -212 4436 -184
rect 4474 -212 4502 -184
rect 4540 -212 4568 -184
rect -4568 -278 -4540 -250
rect -4502 -278 -4474 -250
rect -4436 -278 -4408 -250
rect -4370 -278 -4342 -250
rect -4304 -278 -4276 -250
rect -4238 -278 -4210 -250
rect -4172 -278 -4144 -250
rect -4106 -278 -4078 -250
rect -4040 -278 -4012 -250
rect -3974 -278 -3946 -250
rect -3908 -278 -3880 -250
rect -3842 -278 -3814 -250
rect -3776 -278 -3748 -250
rect -3710 -278 -3682 -250
rect -3644 -278 -3616 -250
rect -3578 -278 -3550 -250
rect -3512 -278 -3484 -250
rect -3446 -278 -3418 -250
rect -3380 -278 -3352 -250
rect -3314 -278 -3286 -250
rect -3248 -278 -3220 -250
rect -3182 -278 -3154 -250
rect -3116 -278 -3088 -250
rect -3050 -278 -3022 -250
rect -2984 -278 -2956 -250
rect -2918 -278 -2890 -250
rect -2852 -278 -2824 -250
rect -2786 -278 -2758 -250
rect -2720 -278 -2692 -250
rect -2654 -278 -2626 -250
rect -2588 -278 -2560 -250
rect -2522 -278 -2494 -250
rect -2456 -278 -2428 -250
rect -2390 -278 -2362 -250
rect -2324 -278 -2296 -250
rect -2258 -278 -2230 -250
rect -2192 -278 -2164 -250
rect -2126 -278 -2098 -250
rect -2060 -278 -2032 -250
rect -1994 -278 -1966 -250
rect -1928 -278 -1900 -250
rect -1862 -278 -1834 -250
rect -1796 -278 -1768 -250
rect -1730 -278 -1702 -250
rect -1664 -278 -1636 -250
rect -1598 -278 -1570 -250
rect -1532 -278 -1504 -250
rect -1466 -278 -1438 -250
rect -1400 -278 -1372 -250
rect -1334 -278 -1306 -250
rect -1268 -278 -1240 -250
rect -1202 -278 -1174 -250
rect -1136 -278 -1108 -250
rect -1070 -278 -1042 -250
rect -1004 -278 -976 -250
rect -938 -278 -910 -250
rect -872 -278 -844 -250
rect -806 -278 -778 -250
rect -740 -278 -712 -250
rect -674 -278 -646 -250
rect -608 -278 -580 -250
rect -542 -278 -514 -250
rect -476 -278 -448 -250
rect -410 -278 -382 -250
rect -344 -278 -316 -250
rect -278 -278 -250 -250
rect -212 -278 -184 -250
rect -146 -278 -118 -250
rect -80 -278 -52 -250
rect -14 -278 14 -250
rect 52 -278 80 -250
rect 118 -278 146 -250
rect 184 -278 212 -250
rect 250 -278 278 -250
rect 316 -278 344 -250
rect 382 -278 410 -250
rect 448 -278 476 -250
rect 514 -278 542 -250
rect 580 -278 608 -250
rect 646 -278 674 -250
rect 712 -278 740 -250
rect 778 -278 806 -250
rect 844 -278 872 -250
rect 910 -278 938 -250
rect 976 -278 1004 -250
rect 1042 -278 1070 -250
rect 1108 -278 1136 -250
rect 1174 -278 1202 -250
rect 1240 -278 1268 -250
rect 1306 -278 1334 -250
rect 1372 -278 1400 -250
rect 1438 -278 1466 -250
rect 1504 -278 1532 -250
rect 1570 -278 1598 -250
rect 1636 -278 1664 -250
rect 1702 -278 1730 -250
rect 1768 -278 1796 -250
rect 1834 -278 1862 -250
rect 1900 -278 1928 -250
rect 1966 -278 1994 -250
rect 2032 -278 2060 -250
rect 2098 -278 2126 -250
rect 2164 -278 2192 -250
rect 2230 -278 2258 -250
rect 2296 -278 2324 -250
rect 2362 -278 2390 -250
rect 2428 -278 2456 -250
rect 2494 -278 2522 -250
rect 2560 -278 2588 -250
rect 2626 -278 2654 -250
rect 2692 -278 2720 -250
rect 2758 -278 2786 -250
rect 2824 -278 2852 -250
rect 2890 -278 2918 -250
rect 2956 -278 2984 -250
rect 3022 -278 3050 -250
rect 3088 -278 3116 -250
rect 3154 -278 3182 -250
rect 3220 -278 3248 -250
rect 3286 -278 3314 -250
rect 3352 -278 3380 -250
rect 3418 -278 3446 -250
rect 3484 -278 3512 -250
rect 3550 -278 3578 -250
rect 3616 -278 3644 -250
rect 3682 -278 3710 -250
rect 3748 -278 3776 -250
rect 3814 -278 3842 -250
rect 3880 -278 3908 -250
rect 3946 -278 3974 -250
rect 4012 -278 4040 -250
rect 4078 -278 4106 -250
rect 4144 -278 4172 -250
rect 4210 -278 4238 -250
rect 4276 -278 4304 -250
rect 4342 -278 4370 -250
rect 4408 -278 4436 -250
rect 4474 -278 4502 -250
rect 4540 -278 4568 -250
rect -4568 -344 -4540 -316
rect -4502 -344 -4474 -316
rect -4436 -344 -4408 -316
rect -4370 -344 -4342 -316
rect -4304 -344 -4276 -316
rect -4238 -344 -4210 -316
rect -4172 -344 -4144 -316
rect -4106 -344 -4078 -316
rect -4040 -344 -4012 -316
rect -3974 -344 -3946 -316
rect -3908 -344 -3880 -316
rect -3842 -344 -3814 -316
rect -3776 -344 -3748 -316
rect -3710 -344 -3682 -316
rect -3644 -344 -3616 -316
rect -3578 -344 -3550 -316
rect -3512 -344 -3484 -316
rect -3446 -344 -3418 -316
rect -3380 -344 -3352 -316
rect -3314 -344 -3286 -316
rect -3248 -344 -3220 -316
rect -3182 -344 -3154 -316
rect -3116 -344 -3088 -316
rect -3050 -344 -3022 -316
rect -2984 -344 -2956 -316
rect -2918 -344 -2890 -316
rect -2852 -344 -2824 -316
rect -2786 -344 -2758 -316
rect -2720 -344 -2692 -316
rect -2654 -344 -2626 -316
rect -2588 -344 -2560 -316
rect -2522 -344 -2494 -316
rect -2456 -344 -2428 -316
rect -2390 -344 -2362 -316
rect -2324 -344 -2296 -316
rect -2258 -344 -2230 -316
rect -2192 -344 -2164 -316
rect -2126 -344 -2098 -316
rect -2060 -344 -2032 -316
rect -1994 -344 -1966 -316
rect -1928 -344 -1900 -316
rect -1862 -344 -1834 -316
rect -1796 -344 -1768 -316
rect -1730 -344 -1702 -316
rect -1664 -344 -1636 -316
rect -1598 -344 -1570 -316
rect -1532 -344 -1504 -316
rect -1466 -344 -1438 -316
rect -1400 -344 -1372 -316
rect -1334 -344 -1306 -316
rect -1268 -344 -1240 -316
rect -1202 -344 -1174 -316
rect -1136 -344 -1108 -316
rect -1070 -344 -1042 -316
rect -1004 -344 -976 -316
rect -938 -344 -910 -316
rect -872 -344 -844 -316
rect -806 -344 -778 -316
rect -740 -344 -712 -316
rect -674 -344 -646 -316
rect -608 -344 -580 -316
rect -542 -344 -514 -316
rect -476 -344 -448 -316
rect -410 -344 -382 -316
rect -344 -344 -316 -316
rect -278 -344 -250 -316
rect -212 -344 -184 -316
rect -146 -344 -118 -316
rect -80 -344 -52 -316
rect -14 -344 14 -316
rect 52 -344 80 -316
rect 118 -344 146 -316
rect 184 -344 212 -316
rect 250 -344 278 -316
rect 316 -344 344 -316
rect 382 -344 410 -316
rect 448 -344 476 -316
rect 514 -344 542 -316
rect 580 -344 608 -316
rect 646 -344 674 -316
rect 712 -344 740 -316
rect 778 -344 806 -316
rect 844 -344 872 -316
rect 910 -344 938 -316
rect 976 -344 1004 -316
rect 1042 -344 1070 -316
rect 1108 -344 1136 -316
rect 1174 -344 1202 -316
rect 1240 -344 1268 -316
rect 1306 -344 1334 -316
rect 1372 -344 1400 -316
rect 1438 -344 1466 -316
rect 1504 -344 1532 -316
rect 1570 -344 1598 -316
rect 1636 -344 1664 -316
rect 1702 -344 1730 -316
rect 1768 -344 1796 -316
rect 1834 -344 1862 -316
rect 1900 -344 1928 -316
rect 1966 -344 1994 -316
rect 2032 -344 2060 -316
rect 2098 -344 2126 -316
rect 2164 -344 2192 -316
rect 2230 -344 2258 -316
rect 2296 -344 2324 -316
rect 2362 -344 2390 -316
rect 2428 -344 2456 -316
rect 2494 -344 2522 -316
rect 2560 -344 2588 -316
rect 2626 -344 2654 -316
rect 2692 -344 2720 -316
rect 2758 -344 2786 -316
rect 2824 -344 2852 -316
rect 2890 -344 2918 -316
rect 2956 -344 2984 -316
rect 3022 -344 3050 -316
rect 3088 -344 3116 -316
rect 3154 -344 3182 -316
rect 3220 -344 3248 -316
rect 3286 -344 3314 -316
rect 3352 -344 3380 -316
rect 3418 -344 3446 -316
rect 3484 -344 3512 -316
rect 3550 -344 3578 -316
rect 3616 -344 3644 -316
rect 3682 -344 3710 -316
rect 3748 -344 3776 -316
rect 3814 -344 3842 -316
rect 3880 -344 3908 -316
rect 3946 -344 3974 -316
rect 4012 -344 4040 -316
rect 4078 -344 4106 -316
rect 4144 -344 4172 -316
rect 4210 -344 4238 -316
rect 4276 -344 4304 -316
rect 4342 -344 4370 -316
rect 4408 -344 4436 -316
rect 4474 -344 4502 -316
rect 4540 -344 4568 -316
rect -4568 -410 -4540 -382
rect -4502 -410 -4474 -382
rect -4436 -410 -4408 -382
rect -4370 -410 -4342 -382
rect -4304 -410 -4276 -382
rect -4238 -410 -4210 -382
rect -4172 -410 -4144 -382
rect -4106 -410 -4078 -382
rect -4040 -410 -4012 -382
rect -3974 -410 -3946 -382
rect -3908 -410 -3880 -382
rect -3842 -410 -3814 -382
rect -3776 -410 -3748 -382
rect -3710 -410 -3682 -382
rect -3644 -410 -3616 -382
rect -3578 -410 -3550 -382
rect -3512 -410 -3484 -382
rect -3446 -410 -3418 -382
rect -3380 -410 -3352 -382
rect -3314 -410 -3286 -382
rect -3248 -410 -3220 -382
rect -3182 -410 -3154 -382
rect -3116 -410 -3088 -382
rect -3050 -410 -3022 -382
rect -2984 -410 -2956 -382
rect -2918 -410 -2890 -382
rect -2852 -410 -2824 -382
rect -2786 -410 -2758 -382
rect -2720 -410 -2692 -382
rect -2654 -410 -2626 -382
rect -2588 -410 -2560 -382
rect -2522 -410 -2494 -382
rect -2456 -410 -2428 -382
rect -2390 -410 -2362 -382
rect -2324 -410 -2296 -382
rect -2258 -410 -2230 -382
rect -2192 -410 -2164 -382
rect -2126 -410 -2098 -382
rect -2060 -410 -2032 -382
rect -1994 -410 -1966 -382
rect -1928 -410 -1900 -382
rect -1862 -410 -1834 -382
rect -1796 -410 -1768 -382
rect -1730 -410 -1702 -382
rect -1664 -410 -1636 -382
rect -1598 -410 -1570 -382
rect -1532 -410 -1504 -382
rect -1466 -410 -1438 -382
rect -1400 -410 -1372 -382
rect -1334 -410 -1306 -382
rect -1268 -410 -1240 -382
rect -1202 -410 -1174 -382
rect -1136 -410 -1108 -382
rect -1070 -410 -1042 -382
rect -1004 -410 -976 -382
rect -938 -410 -910 -382
rect -872 -410 -844 -382
rect -806 -410 -778 -382
rect -740 -410 -712 -382
rect -674 -410 -646 -382
rect -608 -410 -580 -382
rect -542 -410 -514 -382
rect -476 -410 -448 -382
rect -410 -410 -382 -382
rect -344 -410 -316 -382
rect -278 -410 -250 -382
rect -212 -410 -184 -382
rect -146 -410 -118 -382
rect -80 -410 -52 -382
rect -14 -410 14 -382
rect 52 -410 80 -382
rect 118 -410 146 -382
rect 184 -410 212 -382
rect 250 -410 278 -382
rect 316 -410 344 -382
rect 382 -410 410 -382
rect 448 -410 476 -382
rect 514 -410 542 -382
rect 580 -410 608 -382
rect 646 -410 674 -382
rect 712 -410 740 -382
rect 778 -410 806 -382
rect 844 -410 872 -382
rect 910 -410 938 -382
rect 976 -410 1004 -382
rect 1042 -410 1070 -382
rect 1108 -410 1136 -382
rect 1174 -410 1202 -382
rect 1240 -410 1268 -382
rect 1306 -410 1334 -382
rect 1372 -410 1400 -382
rect 1438 -410 1466 -382
rect 1504 -410 1532 -382
rect 1570 -410 1598 -382
rect 1636 -410 1664 -382
rect 1702 -410 1730 -382
rect 1768 -410 1796 -382
rect 1834 -410 1862 -382
rect 1900 -410 1928 -382
rect 1966 -410 1994 -382
rect 2032 -410 2060 -382
rect 2098 -410 2126 -382
rect 2164 -410 2192 -382
rect 2230 -410 2258 -382
rect 2296 -410 2324 -382
rect 2362 -410 2390 -382
rect 2428 -410 2456 -382
rect 2494 -410 2522 -382
rect 2560 -410 2588 -382
rect 2626 -410 2654 -382
rect 2692 -410 2720 -382
rect 2758 -410 2786 -382
rect 2824 -410 2852 -382
rect 2890 -410 2918 -382
rect 2956 -410 2984 -382
rect 3022 -410 3050 -382
rect 3088 -410 3116 -382
rect 3154 -410 3182 -382
rect 3220 -410 3248 -382
rect 3286 -410 3314 -382
rect 3352 -410 3380 -382
rect 3418 -410 3446 -382
rect 3484 -410 3512 -382
rect 3550 -410 3578 -382
rect 3616 -410 3644 -382
rect 3682 -410 3710 -382
rect 3748 -410 3776 -382
rect 3814 -410 3842 -382
rect 3880 -410 3908 -382
rect 3946 -410 3974 -382
rect 4012 -410 4040 -382
rect 4078 -410 4106 -382
rect 4144 -410 4172 -382
rect 4210 -410 4238 -382
rect 4276 -410 4304 -382
rect 4342 -410 4370 -382
rect 4408 -410 4436 -382
rect 4474 -410 4502 -382
rect 4540 -410 4568 -382
rect -4568 -476 -4540 -448
rect -4502 -476 -4474 -448
rect -4436 -476 -4408 -448
rect -4370 -476 -4342 -448
rect -4304 -476 -4276 -448
rect -4238 -476 -4210 -448
rect -4172 -476 -4144 -448
rect -4106 -476 -4078 -448
rect -4040 -476 -4012 -448
rect -3974 -476 -3946 -448
rect -3908 -476 -3880 -448
rect -3842 -476 -3814 -448
rect -3776 -476 -3748 -448
rect -3710 -476 -3682 -448
rect -3644 -476 -3616 -448
rect -3578 -476 -3550 -448
rect -3512 -476 -3484 -448
rect -3446 -476 -3418 -448
rect -3380 -476 -3352 -448
rect -3314 -476 -3286 -448
rect -3248 -476 -3220 -448
rect -3182 -476 -3154 -448
rect -3116 -476 -3088 -448
rect -3050 -476 -3022 -448
rect -2984 -476 -2956 -448
rect -2918 -476 -2890 -448
rect -2852 -476 -2824 -448
rect -2786 -476 -2758 -448
rect -2720 -476 -2692 -448
rect -2654 -476 -2626 -448
rect -2588 -476 -2560 -448
rect -2522 -476 -2494 -448
rect -2456 -476 -2428 -448
rect -2390 -476 -2362 -448
rect -2324 -476 -2296 -448
rect -2258 -476 -2230 -448
rect -2192 -476 -2164 -448
rect -2126 -476 -2098 -448
rect -2060 -476 -2032 -448
rect -1994 -476 -1966 -448
rect -1928 -476 -1900 -448
rect -1862 -476 -1834 -448
rect -1796 -476 -1768 -448
rect -1730 -476 -1702 -448
rect -1664 -476 -1636 -448
rect -1598 -476 -1570 -448
rect -1532 -476 -1504 -448
rect -1466 -476 -1438 -448
rect -1400 -476 -1372 -448
rect -1334 -476 -1306 -448
rect -1268 -476 -1240 -448
rect -1202 -476 -1174 -448
rect -1136 -476 -1108 -448
rect -1070 -476 -1042 -448
rect -1004 -476 -976 -448
rect -938 -476 -910 -448
rect -872 -476 -844 -448
rect -806 -476 -778 -448
rect -740 -476 -712 -448
rect -674 -476 -646 -448
rect -608 -476 -580 -448
rect -542 -476 -514 -448
rect -476 -476 -448 -448
rect -410 -476 -382 -448
rect -344 -476 -316 -448
rect -278 -476 -250 -448
rect -212 -476 -184 -448
rect -146 -476 -118 -448
rect -80 -476 -52 -448
rect -14 -476 14 -448
rect 52 -476 80 -448
rect 118 -476 146 -448
rect 184 -476 212 -448
rect 250 -476 278 -448
rect 316 -476 344 -448
rect 382 -476 410 -448
rect 448 -476 476 -448
rect 514 -476 542 -448
rect 580 -476 608 -448
rect 646 -476 674 -448
rect 712 -476 740 -448
rect 778 -476 806 -448
rect 844 -476 872 -448
rect 910 -476 938 -448
rect 976 -476 1004 -448
rect 1042 -476 1070 -448
rect 1108 -476 1136 -448
rect 1174 -476 1202 -448
rect 1240 -476 1268 -448
rect 1306 -476 1334 -448
rect 1372 -476 1400 -448
rect 1438 -476 1466 -448
rect 1504 -476 1532 -448
rect 1570 -476 1598 -448
rect 1636 -476 1664 -448
rect 1702 -476 1730 -448
rect 1768 -476 1796 -448
rect 1834 -476 1862 -448
rect 1900 -476 1928 -448
rect 1966 -476 1994 -448
rect 2032 -476 2060 -448
rect 2098 -476 2126 -448
rect 2164 -476 2192 -448
rect 2230 -476 2258 -448
rect 2296 -476 2324 -448
rect 2362 -476 2390 -448
rect 2428 -476 2456 -448
rect 2494 -476 2522 -448
rect 2560 -476 2588 -448
rect 2626 -476 2654 -448
rect 2692 -476 2720 -448
rect 2758 -476 2786 -448
rect 2824 -476 2852 -448
rect 2890 -476 2918 -448
rect 2956 -476 2984 -448
rect 3022 -476 3050 -448
rect 3088 -476 3116 -448
rect 3154 -476 3182 -448
rect 3220 -476 3248 -448
rect 3286 -476 3314 -448
rect 3352 -476 3380 -448
rect 3418 -476 3446 -448
rect 3484 -476 3512 -448
rect 3550 -476 3578 -448
rect 3616 -476 3644 -448
rect 3682 -476 3710 -448
rect 3748 -476 3776 -448
rect 3814 -476 3842 -448
rect 3880 -476 3908 -448
rect 3946 -476 3974 -448
rect 4012 -476 4040 -448
rect 4078 -476 4106 -448
rect 4144 -476 4172 -448
rect 4210 -476 4238 -448
rect 4276 -476 4304 -448
rect 4342 -476 4370 -448
rect 4408 -476 4436 -448
rect 4474 -476 4502 -448
rect 4540 -476 4568 -448
rect -4568 -542 -4540 -514
rect -4502 -542 -4474 -514
rect -4436 -542 -4408 -514
rect -4370 -542 -4342 -514
rect -4304 -542 -4276 -514
rect -4238 -542 -4210 -514
rect -4172 -542 -4144 -514
rect -4106 -542 -4078 -514
rect -4040 -542 -4012 -514
rect -3974 -542 -3946 -514
rect -3908 -542 -3880 -514
rect -3842 -542 -3814 -514
rect -3776 -542 -3748 -514
rect -3710 -542 -3682 -514
rect -3644 -542 -3616 -514
rect -3578 -542 -3550 -514
rect -3512 -542 -3484 -514
rect -3446 -542 -3418 -514
rect -3380 -542 -3352 -514
rect -3314 -542 -3286 -514
rect -3248 -542 -3220 -514
rect -3182 -542 -3154 -514
rect -3116 -542 -3088 -514
rect -3050 -542 -3022 -514
rect -2984 -542 -2956 -514
rect -2918 -542 -2890 -514
rect -2852 -542 -2824 -514
rect -2786 -542 -2758 -514
rect -2720 -542 -2692 -514
rect -2654 -542 -2626 -514
rect -2588 -542 -2560 -514
rect -2522 -542 -2494 -514
rect -2456 -542 -2428 -514
rect -2390 -542 -2362 -514
rect -2324 -542 -2296 -514
rect -2258 -542 -2230 -514
rect -2192 -542 -2164 -514
rect -2126 -542 -2098 -514
rect -2060 -542 -2032 -514
rect -1994 -542 -1966 -514
rect -1928 -542 -1900 -514
rect -1862 -542 -1834 -514
rect -1796 -542 -1768 -514
rect -1730 -542 -1702 -514
rect -1664 -542 -1636 -514
rect -1598 -542 -1570 -514
rect -1532 -542 -1504 -514
rect -1466 -542 -1438 -514
rect -1400 -542 -1372 -514
rect -1334 -542 -1306 -514
rect -1268 -542 -1240 -514
rect -1202 -542 -1174 -514
rect -1136 -542 -1108 -514
rect -1070 -542 -1042 -514
rect -1004 -542 -976 -514
rect -938 -542 -910 -514
rect -872 -542 -844 -514
rect -806 -542 -778 -514
rect -740 -542 -712 -514
rect -674 -542 -646 -514
rect -608 -542 -580 -514
rect -542 -542 -514 -514
rect -476 -542 -448 -514
rect -410 -542 -382 -514
rect -344 -542 -316 -514
rect -278 -542 -250 -514
rect -212 -542 -184 -514
rect -146 -542 -118 -514
rect -80 -542 -52 -514
rect -14 -542 14 -514
rect 52 -542 80 -514
rect 118 -542 146 -514
rect 184 -542 212 -514
rect 250 -542 278 -514
rect 316 -542 344 -514
rect 382 -542 410 -514
rect 448 -542 476 -514
rect 514 -542 542 -514
rect 580 -542 608 -514
rect 646 -542 674 -514
rect 712 -542 740 -514
rect 778 -542 806 -514
rect 844 -542 872 -514
rect 910 -542 938 -514
rect 976 -542 1004 -514
rect 1042 -542 1070 -514
rect 1108 -542 1136 -514
rect 1174 -542 1202 -514
rect 1240 -542 1268 -514
rect 1306 -542 1334 -514
rect 1372 -542 1400 -514
rect 1438 -542 1466 -514
rect 1504 -542 1532 -514
rect 1570 -542 1598 -514
rect 1636 -542 1664 -514
rect 1702 -542 1730 -514
rect 1768 -542 1796 -514
rect 1834 -542 1862 -514
rect 1900 -542 1928 -514
rect 1966 -542 1994 -514
rect 2032 -542 2060 -514
rect 2098 -542 2126 -514
rect 2164 -542 2192 -514
rect 2230 -542 2258 -514
rect 2296 -542 2324 -514
rect 2362 -542 2390 -514
rect 2428 -542 2456 -514
rect 2494 -542 2522 -514
rect 2560 -542 2588 -514
rect 2626 -542 2654 -514
rect 2692 -542 2720 -514
rect 2758 -542 2786 -514
rect 2824 -542 2852 -514
rect 2890 -542 2918 -514
rect 2956 -542 2984 -514
rect 3022 -542 3050 -514
rect 3088 -542 3116 -514
rect 3154 -542 3182 -514
rect 3220 -542 3248 -514
rect 3286 -542 3314 -514
rect 3352 -542 3380 -514
rect 3418 -542 3446 -514
rect 3484 -542 3512 -514
rect 3550 -542 3578 -514
rect 3616 -542 3644 -514
rect 3682 -542 3710 -514
rect 3748 -542 3776 -514
rect 3814 -542 3842 -514
rect 3880 -542 3908 -514
rect 3946 -542 3974 -514
rect 4012 -542 4040 -514
rect 4078 -542 4106 -514
rect 4144 -542 4172 -514
rect 4210 -542 4238 -514
rect 4276 -542 4304 -514
rect 4342 -542 4370 -514
rect 4408 -542 4436 -514
rect 4474 -542 4502 -514
rect 4540 -542 4568 -514
rect -4568 -608 -4540 -580
rect -4502 -608 -4474 -580
rect -4436 -608 -4408 -580
rect -4370 -608 -4342 -580
rect -4304 -608 -4276 -580
rect -4238 -608 -4210 -580
rect -4172 -608 -4144 -580
rect -4106 -608 -4078 -580
rect -4040 -608 -4012 -580
rect -3974 -608 -3946 -580
rect -3908 -608 -3880 -580
rect -3842 -608 -3814 -580
rect -3776 -608 -3748 -580
rect -3710 -608 -3682 -580
rect -3644 -608 -3616 -580
rect -3578 -608 -3550 -580
rect -3512 -608 -3484 -580
rect -3446 -608 -3418 -580
rect -3380 -608 -3352 -580
rect -3314 -608 -3286 -580
rect -3248 -608 -3220 -580
rect -3182 -608 -3154 -580
rect -3116 -608 -3088 -580
rect -3050 -608 -3022 -580
rect -2984 -608 -2956 -580
rect -2918 -608 -2890 -580
rect -2852 -608 -2824 -580
rect -2786 -608 -2758 -580
rect -2720 -608 -2692 -580
rect -2654 -608 -2626 -580
rect -2588 -608 -2560 -580
rect -2522 -608 -2494 -580
rect -2456 -608 -2428 -580
rect -2390 -608 -2362 -580
rect -2324 -608 -2296 -580
rect -2258 -608 -2230 -580
rect -2192 -608 -2164 -580
rect -2126 -608 -2098 -580
rect -2060 -608 -2032 -580
rect -1994 -608 -1966 -580
rect -1928 -608 -1900 -580
rect -1862 -608 -1834 -580
rect -1796 -608 -1768 -580
rect -1730 -608 -1702 -580
rect -1664 -608 -1636 -580
rect -1598 -608 -1570 -580
rect -1532 -608 -1504 -580
rect -1466 -608 -1438 -580
rect -1400 -608 -1372 -580
rect -1334 -608 -1306 -580
rect -1268 -608 -1240 -580
rect -1202 -608 -1174 -580
rect -1136 -608 -1108 -580
rect -1070 -608 -1042 -580
rect -1004 -608 -976 -580
rect -938 -608 -910 -580
rect -872 -608 -844 -580
rect -806 -608 -778 -580
rect -740 -608 -712 -580
rect -674 -608 -646 -580
rect -608 -608 -580 -580
rect -542 -608 -514 -580
rect -476 -608 -448 -580
rect -410 -608 -382 -580
rect -344 -608 -316 -580
rect -278 -608 -250 -580
rect -212 -608 -184 -580
rect -146 -608 -118 -580
rect -80 -608 -52 -580
rect -14 -608 14 -580
rect 52 -608 80 -580
rect 118 -608 146 -580
rect 184 -608 212 -580
rect 250 -608 278 -580
rect 316 -608 344 -580
rect 382 -608 410 -580
rect 448 -608 476 -580
rect 514 -608 542 -580
rect 580 -608 608 -580
rect 646 -608 674 -580
rect 712 -608 740 -580
rect 778 -608 806 -580
rect 844 -608 872 -580
rect 910 -608 938 -580
rect 976 -608 1004 -580
rect 1042 -608 1070 -580
rect 1108 -608 1136 -580
rect 1174 -608 1202 -580
rect 1240 -608 1268 -580
rect 1306 -608 1334 -580
rect 1372 -608 1400 -580
rect 1438 -608 1466 -580
rect 1504 -608 1532 -580
rect 1570 -608 1598 -580
rect 1636 -608 1664 -580
rect 1702 -608 1730 -580
rect 1768 -608 1796 -580
rect 1834 -608 1862 -580
rect 1900 -608 1928 -580
rect 1966 -608 1994 -580
rect 2032 -608 2060 -580
rect 2098 -608 2126 -580
rect 2164 -608 2192 -580
rect 2230 -608 2258 -580
rect 2296 -608 2324 -580
rect 2362 -608 2390 -580
rect 2428 -608 2456 -580
rect 2494 -608 2522 -580
rect 2560 -608 2588 -580
rect 2626 -608 2654 -580
rect 2692 -608 2720 -580
rect 2758 -608 2786 -580
rect 2824 -608 2852 -580
rect 2890 -608 2918 -580
rect 2956 -608 2984 -580
rect 3022 -608 3050 -580
rect 3088 -608 3116 -580
rect 3154 -608 3182 -580
rect 3220 -608 3248 -580
rect 3286 -608 3314 -580
rect 3352 -608 3380 -580
rect 3418 -608 3446 -580
rect 3484 -608 3512 -580
rect 3550 -608 3578 -580
rect 3616 -608 3644 -580
rect 3682 -608 3710 -580
rect 3748 -608 3776 -580
rect 3814 -608 3842 -580
rect 3880 -608 3908 -580
rect 3946 -608 3974 -580
rect 4012 -608 4040 -580
rect 4078 -608 4106 -580
rect 4144 -608 4172 -580
rect 4210 -608 4238 -580
rect 4276 -608 4304 -580
rect 4342 -608 4370 -580
rect 4408 -608 4436 -580
rect 4474 -608 4502 -580
rect 4540 -608 4568 -580
rect -4568 -674 -4540 -646
rect -4502 -674 -4474 -646
rect -4436 -674 -4408 -646
rect -4370 -674 -4342 -646
rect -4304 -674 -4276 -646
rect -4238 -674 -4210 -646
rect -4172 -674 -4144 -646
rect -4106 -674 -4078 -646
rect -4040 -674 -4012 -646
rect -3974 -674 -3946 -646
rect -3908 -674 -3880 -646
rect -3842 -674 -3814 -646
rect -3776 -674 -3748 -646
rect -3710 -674 -3682 -646
rect -3644 -674 -3616 -646
rect -3578 -674 -3550 -646
rect -3512 -674 -3484 -646
rect -3446 -674 -3418 -646
rect -3380 -674 -3352 -646
rect -3314 -674 -3286 -646
rect -3248 -674 -3220 -646
rect -3182 -674 -3154 -646
rect -3116 -674 -3088 -646
rect -3050 -674 -3022 -646
rect -2984 -674 -2956 -646
rect -2918 -674 -2890 -646
rect -2852 -674 -2824 -646
rect -2786 -674 -2758 -646
rect -2720 -674 -2692 -646
rect -2654 -674 -2626 -646
rect -2588 -674 -2560 -646
rect -2522 -674 -2494 -646
rect -2456 -674 -2428 -646
rect -2390 -674 -2362 -646
rect -2324 -674 -2296 -646
rect -2258 -674 -2230 -646
rect -2192 -674 -2164 -646
rect -2126 -674 -2098 -646
rect -2060 -674 -2032 -646
rect -1994 -674 -1966 -646
rect -1928 -674 -1900 -646
rect -1862 -674 -1834 -646
rect -1796 -674 -1768 -646
rect -1730 -674 -1702 -646
rect -1664 -674 -1636 -646
rect -1598 -674 -1570 -646
rect -1532 -674 -1504 -646
rect -1466 -674 -1438 -646
rect -1400 -674 -1372 -646
rect -1334 -674 -1306 -646
rect -1268 -674 -1240 -646
rect -1202 -674 -1174 -646
rect -1136 -674 -1108 -646
rect -1070 -674 -1042 -646
rect -1004 -674 -976 -646
rect -938 -674 -910 -646
rect -872 -674 -844 -646
rect -806 -674 -778 -646
rect -740 -674 -712 -646
rect -674 -674 -646 -646
rect -608 -674 -580 -646
rect -542 -674 -514 -646
rect -476 -674 -448 -646
rect -410 -674 -382 -646
rect -344 -674 -316 -646
rect -278 -674 -250 -646
rect -212 -674 -184 -646
rect -146 -674 -118 -646
rect -80 -674 -52 -646
rect -14 -674 14 -646
rect 52 -674 80 -646
rect 118 -674 146 -646
rect 184 -674 212 -646
rect 250 -674 278 -646
rect 316 -674 344 -646
rect 382 -674 410 -646
rect 448 -674 476 -646
rect 514 -674 542 -646
rect 580 -674 608 -646
rect 646 -674 674 -646
rect 712 -674 740 -646
rect 778 -674 806 -646
rect 844 -674 872 -646
rect 910 -674 938 -646
rect 976 -674 1004 -646
rect 1042 -674 1070 -646
rect 1108 -674 1136 -646
rect 1174 -674 1202 -646
rect 1240 -674 1268 -646
rect 1306 -674 1334 -646
rect 1372 -674 1400 -646
rect 1438 -674 1466 -646
rect 1504 -674 1532 -646
rect 1570 -674 1598 -646
rect 1636 -674 1664 -646
rect 1702 -674 1730 -646
rect 1768 -674 1796 -646
rect 1834 -674 1862 -646
rect 1900 -674 1928 -646
rect 1966 -674 1994 -646
rect 2032 -674 2060 -646
rect 2098 -674 2126 -646
rect 2164 -674 2192 -646
rect 2230 -674 2258 -646
rect 2296 -674 2324 -646
rect 2362 -674 2390 -646
rect 2428 -674 2456 -646
rect 2494 -674 2522 -646
rect 2560 -674 2588 -646
rect 2626 -674 2654 -646
rect 2692 -674 2720 -646
rect 2758 -674 2786 -646
rect 2824 -674 2852 -646
rect 2890 -674 2918 -646
rect 2956 -674 2984 -646
rect 3022 -674 3050 -646
rect 3088 -674 3116 -646
rect 3154 -674 3182 -646
rect 3220 -674 3248 -646
rect 3286 -674 3314 -646
rect 3352 -674 3380 -646
rect 3418 -674 3446 -646
rect 3484 -674 3512 -646
rect 3550 -674 3578 -646
rect 3616 -674 3644 -646
rect 3682 -674 3710 -646
rect 3748 -674 3776 -646
rect 3814 -674 3842 -646
rect 3880 -674 3908 -646
rect 3946 -674 3974 -646
rect 4012 -674 4040 -646
rect 4078 -674 4106 -646
rect 4144 -674 4172 -646
rect 4210 -674 4238 -646
rect 4276 -674 4304 -646
rect 4342 -674 4370 -646
rect 4408 -674 4436 -646
rect 4474 -674 4502 -646
rect 4540 -674 4568 -646
rect -4568 -740 -4540 -712
rect -4502 -740 -4474 -712
rect -4436 -740 -4408 -712
rect -4370 -740 -4342 -712
rect -4304 -740 -4276 -712
rect -4238 -740 -4210 -712
rect -4172 -740 -4144 -712
rect -4106 -740 -4078 -712
rect -4040 -740 -4012 -712
rect -3974 -740 -3946 -712
rect -3908 -740 -3880 -712
rect -3842 -740 -3814 -712
rect -3776 -740 -3748 -712
rect -3710 -740 -3682 -712
rect -3644 -740 -3616 -712
rect -3578 -740 -3550 -712
rect -3512 -740 -3484 -712
rect -3446 -740 -3418 -712
rect -3380 -740 -3352 -712
rect -3314 -740 -3286 -712
rect -3248 -740 -3220 -712
rect -3182 -740 -3154 -712
rect -3116 -740 -3088 -712
rect -3050 -740 -3022 -712
rect -2984 -740 -2956 -712
rect -2918 -740 -2890 -712
rect -2852 -740 -2824 -712
rect -2786 -740 -2758 -712
rect -2720 -740 -2692 -712
rect -2654 -740 -2626 -712
rect -2588 -740 -2560 -712
rect -2522 -740 -2494 -712
rect -2456 -740 -2428 -712
rect -2390 -740 -2362 -712
rect -2324 -740 -2296 -712
rect -2258 -740 -2230 -712
rect -2192 -740 -2164 -712
rect -2126 -740 -2098 -712
rect -2060 -740 -2032 -712
rect -1994 -740 -1966 -712
rect -1928 -740 -1900 -712
rect -1862 -740 -1834 -712
rect -1796 -740 -1768 -712
rect -1730 -740 -1702 -712
rect -1664 -740 -1636 -712
rect -1598 -740 -1570 -712
rect -1532 -740 -1504 -712
rect -1466 -740 -1438 -712
rect -1400 -740 -1372 -712
rect -1334 -740 -1306 -712
rect -1268 -740 -1240 -712
rect -1202 -740 -1174 -712
rect -1136 -740 -1108 -712
rect -1070 -740 -1042 -712
rect -1004 -740 -976 -712
rect -938 -740 -910 -712
rect -872 -740 -844 -712
rect -806 -740 -778 -712
rect -740 -740 -712 -712
rect -674 -740 -646 -712
rect -608 -740 -580 -712
rect -542 -740 -514 -712
rect -476 -740 -448 -712
rect -410 -740 -382 -712
rect -344 -740 -316 -712
rect -278 -740 -250 -712
rect -212 -740 -184 -712
rect -146 -740 -118 -712
rect -80 -740 -52 -712
rect -14 -740 14 -712
rect 52 -740 80 -712
rect 118 -740 146 -712
rect 184 -740 212 -712
rect 250 -740 278 -712
rect 316 -740 344 -712
rect 382 -740 410 -712
rect 448 -740 476 -712
rect 514 -740 542 -712
rect 580 -740 608 -712
rect 646 -740 674 -712
rect 712 -740 740 -712
rect 778 -740 806 -712
rect 844 -740 872 -712
rect 910 -740 938 -712
rect 976 -740 1004 -712
rect 1042 -740 1070 -712
rect 1108 -740 1136 -712
rect 1174 -740 1202 -712
rect 1240 -740 1268 -712
rect 1306 -740 1334 -712
rect 1372 -740 1400 -712
rect 1438 -740 1466 -712
rect 1504 -740 1532 -712
rect 1570 -740 1598 -712
rect 1636 -740 1664 -712
rect 1702 -740 1730 -712
rect 1768 -740 1796 -712
rect 1834 -740 1862 -712
rect 1900 -740 1928 -712
rect 1966 -740 1994 -712
rect 2032 -740 2060 -712
rect 2098 -740 2126 -712
rect 2164 -740 2192 -712
rect 2230 -740 2258 -712
rect 2296 -740 2324 -712
rect 2362 -740 2390 -712
rect 2428 -740 2456 -712
rect 2494 -740 2522 -712
rect 2560 -740 2588 -712
rect 2626 -740 2654 -712
rect 2692 -740 2720 -712
rect 2758 -740 2786 -712
rect 2824 -740 2852 -712
rect 2890 -740 2918 -712
rect 2956 -740 2984 -712
rect 3022 -740 3050 -712
rect 3088 -740 3116 -712
rect 3154 -740 3182 -712
rect 3220 -740 3248 -712
rect 3286 -740 3314 -712
rect 3352 -740 3380 -712
rect 3418 -740 3446 -712
rect 3484 -740 3512 -712
rect 3550 -740 3578 -712
rect 3616 -740 3644 -712
rect 3682 -740 3710 -712
rect 3748 -740 3776 -712
rect 3814 -740 3842 -712
rect 3880 -740 3908 -712
rect 3946 -740 3974 -712
rect 4012 -740 4040 -712
rect 4078 -740 4106 -712
rect 4144 -740 4172 -712
rect 4210 -740 4238 -712
rect 4276 -740 4304 -712
rect 4342 -740 4370 -712
rect 4408 -740 4436 -712
rect 4474 -740 4502 -712
rect 4540 -740 4568 -712
<< metal4 >>
rect -4573 740 4573 745
rect -4573 712 -4568 740
rect -4540 712 -4502 740
rect -4474 712 -4436 740
rect -4408 712 -4370 740
rect -4342 712 -4304 740
rect -4276 712 -4238 740
rect -4210 712 -4172 740
rect -4144 712 -4106 740
rect -4078 712 -4040 740
rect -4012 712 -3974 740
rect -3946 712 -3908 740
rect -3880 712 -3842 740
rect -3814 712 -3776 740
rect -3748 712 -3710 740
rect -3682 712 -3644 740
rect -3616 712 -3578 740
rect -3550 712 -3512 740
rect -3484 712 -3446 740
rect -3418 712 -3380 740
rect -3352 712 -3314 740
rect -3286 712 -3248 740
rect -3220 712 -3182 740
rect -3154 712 -3116 740
rect -3088 712 -3050 740
rect -3022 712 -2984 740
rect -2956 712 -2918 740
rect -2890 712 -2852 740
rect -2824 712 -2786 740
rect -2758 712 -2720 740
rect -2692 712 -2654 740
rect -2626 712 -2588 740
rect -2560 712 -2522 740
rect -2494 712 -2456 740
rect -2428 712 -2390 740
rect -2362 712 -2324 740
rect -2296 712 -2258 740
rect -2230 712 -2192 740
rect -2164 712 -2126 740
rect -2098 712 -2060 740
rect -2032 712 -1994 740
rect -1966 712 -1928 740
rect -1900 712 -1862 740
rect -1834 712 -1796 740
rect -1768 712 -1730 740
rect -1702 712 -1664 740
rect -1636 712 -1598 740
rect -1570 712 -1532 740
rect -1504 712 -1466 740
rect -1438 712 -1400 740
rect -1372 712 -1334 740
rect -1306 712 -1268 740
rect -1240 712 -1202 740
rect -1174 712 -1136 740
rect -1108 712 -1070 740
rect -1042 712 -1004 740
rect -976 712 -938 740
rect -910 712 -872 740
rect -844 712 -806 740
rect -778 712 -740 740
rect -712 712 -674 740
rect -646 712 -608 740
rect -580 712 -542 740
rect -514 712 -476 740
rect -448 712 -410 740
rect -382 712 -344 740
rect -316 712 -278 740
rect -250 712 -212 740
rect -184 712 -146 740
rect -118 712 -80 740
rect -52 712 -14 740
rect 14 712 52 740
rect 80 712 118 740
rect 146 712 184 740
rect 212 712 250 740
rect 278 712 316 740
rect 344 712 382 740
rect 410 712 448 740
rect 476 712 514 740
rect 542 712 580 740
rect 608 712 646 740
rect 674 712 712 740
rect 740 712 778 740
rect 806 712 844 740
rect 872 712 910 740
rect 938 712 976 740
rect 1004 712 1042 740
rect 1070 712 1108 740
rect 1136 712 1174 740
rect 1202 712 1240 740
rect 1268 712 1306 740
rect 1334 712 1372 740
rect 1400 712 1438 740
rect 1466 712 1504 740
rect 1532 712 1570 740
rect 1598 712 1636 740
rect 1664 712 1702 740
rect 1730 712 1768 740
rect 1796 712 1834 740
rect 1862 712 1900 740
rect 1928 712 1966 740
rect 1994 712 2032 740
rect 2060 712 2098 740
rect 2126 712 2164 740
rect 2192 712 2230 740
rect 2258 712 2296 740
rect 2324 712 2362 740
rect 2390 712 2428 740
rect 2456 712 2494 740
rect 2522 712 2560 740
rect 2588 712 2626 740
rect 2654 712 2692 740
rect 2720 712 2758 740
rect 2786 712 2824 740
rect 2852 712 2890 740
rect 2918 712 2956 740
rect 2984 712 3022 740
rect 3050 712 3088 740
rect 3116 712 3154 740
rect 3182 712 3220 740
rect 3248 712 3286 740
rect 3314 712 3352 740
rect 3380 712 3418 740
rect 3446 712 3484 740
rect 3512 712 3550 740
rect 3578 712 3616 740
rect 3644 712 3682 740
rect 3710 712 3748 740
rect 3776 712 3814 740
rect 3842 712 3880 740
rect 3908 712 3946 740
rect 3974 712 4012 740
rect 4040 712 4078 740
rect 4106 712 4144 740
rect 4172 712 4210 740
rect 4238 712 4276 740
rect 4304 712 4342 740
rect 4370 712 4408 740
rect 4436 712 4474 740
rect 4502 712 4540 740
rect 4568 712 4573 740
rect -4573 674 4573 712
rect -4573 646 -4568 674
rect -4540 646 -4502 674
rect -4474 646 -4436 674
rect -4408 646 -4370 674
rect -4342 646 -4304 674
rect -4276 646 -4238 674
rect -4210 646 -4172 674
rect -4144 646 -4106 674
rect -4078 646 -4040 674
rect -4012 646 -3974 674
rect -3946 646 -3908 674
rect -3880 646 -3842 674
rect -3814 646 -3776 674
rect -3748 646 -3710 674
rect -3682 646 -3644 674
rect -3616 646 -3578 674
rect -3550 646 -3512 674
rect -3484 646 -3446 674
rect -3418 646 -3380 674
rect -3352 646 -3314 674
rect -3286 646 -3248 674
rect -3220 646 -3182 674
rect -3154 646 -3116 674
rect -3088 646 -3050 674
rect -3022 646 -2984 674
rect -2956 646 -2918 674
rect -2890 646 -2852 674
rect -2824 646 -2786 674
rect -2758 646 -2720 674
rect -2692 646 -2654 674
rect -2626 646 -2588 674
rect -2560 646 -2522 674
rect -2494 646 -2456 674
rect -2428 646 -2390 674
rect -2362 646 -2324 674
rect -2296 646 -2258 674
rect -2230 646 -2192 674
rect -2164 646 -2126 674
rect -2098 646 -2060 674
rect -2032 646 -1994 674
rect -1966 646 -1928 674
rect -1900 646 -1862 674
rect -1834 646 -1796 674
rect -1768 646 -1730 674
rect -1702 646 -1664 674
rect -1636 646 -1598 674
rect -1570 646 -1532 674
rect -1504 646 -1466 674
rect -1438 646 -1400 674
rect -1372 646 -1334 674
rect -1306 646 -1268 674
rect -1240 646 -1202 674
rect -1174 646 -1136 674
rect -1108 646 -1070 674
rect -1042 646 -1004 674
rect -976 646 -938 674
rect -910 646 -872 674
rect -844 646 -806 674
rect -778 646 -740 674
rect -712 646 -674 674
rect -646 646 -608 674
rect -580 646 -542 674
rect -514 646 -476 674
rect -448 646 -410 674
rect -382 646 -344 674
rect -316 646 -278 674
rect -250 646 -212 674
rect -184 646 -146 674
rect -118 646 -80 674
rect -52 646 -14 674
rect 14 646 52 674
rect 80 646 118 674
rect 146 646 184 674
rect 212 646 250 674
rect 278 646 316 674
rect 344 646 382 674
rect 410 646 448 674
rect 476 646 514 674
rect 542 646 580 674
rect 608 646 646 674
rect 674 646 712 674
rect 740 646 778 674
rect 806 646 844 674
rect 872 646 910 674
rect 938 646 976 674
rect 1004 646 1042 674
rect 1070 646 1108 674
rect 1136 646 1174 674
rect 1202 646 1240 674
rect 1268 646 1306 674
rect 1334 646 1372 674
rect 1400 646 1438 674
rect 1466 646 1504 674
rect 1532 646 1570 674
rect 1598 646 1636 674
rect 1664 646 1702 674
rect 1730 646 1768 674
rect 1796 646 1834 674
rect 1862 646 1900 674
rect 1928 646 1966 674
rect 1994 646 2032 674
rect 2060 646 2098 674
rect 2126 646 2164 674
rect 2192 646 2230 674
rect 2258 646 2296 674
rect 2324 646 2362 674
rect 2390 646 2428 674
rect 2456 646 2494 674
rect 2522 646 2560 674
rect 2588 646 2626 674
rect 2654 646 2692 674
rect 2720 646 2758 674
rect 2786 646 2824 674
rect 2852 646 2890 674
rect 2918 646 2956 674
rect 2984 646 3022 674
rect 3050 646 3088 674
rect 3116 646 3154 674
rect 3182 646 3220 674
rect 3248 646 3286 674
rect 3314 646 3352 674
rect 3380 646 3418 674
rect 3446 646 3484 674
rect 3512 646 3550 674
rect 3578 646 3616 674
rect 3644 646 3682 674
rect 3710 646 3748 674
rect 3776 646 3814 674
rect 3842 646 3880 674
rect 3908 646 3946 674
rect 3974 646 4012 674
rect 4040 646 4078 674
rect 4106 646 4144 674
rect 4172 646 4210 674
rect 4238 646 4276 674
rect 4304 646 4342 674
rect 4370 646 4408 674
rect 4436 646 4474 674
rect 4502 646 4540 674
rect 4568 646 4573 674
rect -4573 608 4573 646
rect -4573 580 -4568 608
rect -4540 580 -4502 608
rect -4474 580 -4436 608
rect -4408 580 -4370 608
rect -4342 580 -4304 608
rect -4276 580 -4238 608
rect -4210 580 -4172 608
rect -4144 580 -4106 608
rect -4078 580 -4040 608
rect -4012 580 -3974 608
rect -3946 580 -3908 608
rect -3880 580 -3842 608
rect -3814 580 -3776 608
rect -3748 580 -3710 608
rect -3682 580 -3644 608
rect -3616 580 -3578 608
rect -3550 580 -3512 608
rect -3484 580 -3446 608
rect -3418 580 -3380 608
rect -3352 580 -3314 608
rect -3286 580 -3248 608
rect -3220 580 -3182 608
rect -3154 580 -3116 608
rect -3088 580 -3050 608
rect -3022 580 -2984 608
rect -2956 580 -2918 608
rect -2890 580 -2852 608
rect -2824 580 -2786 608
rect -2758 580 -2720 608
rect -2692 580 -2654 608
rect -2626 580 -2588 608
rect -2560 580 -2522 608
rect -2494 580 -2456 608
rect -2428 580 -2390 608
rect -2362 580 -2324 608
rect -2296 580 -2258 608
rect -2230 580 -2192 608
rect -2164 580 -2126 608
rect -2098 580 -2060 608
rect -2032 580 -1994 608
rect -1966 580 -1928 608
rect -1900 580 -1862 608
rect -1834 580 -1796 608
rect -1768 580 -1730 608
rect -1702 580 -1664 608
rect -1636 580 -1598 608
rect -1570 580 -1532 608
rect -1504 580 -1466 608
rect -1438 580 -1400 608
rect -1372 580 -1334 608
rect -1306 580 -1268 608
rect -1240 580 -1202 608
rect -1174 580 -1136 608
rect -1108 580 -1070 608
rect -1042 580 -1004 608
rect -976 580 -938 608
rect -910 580 -872 608
rect -844 580 -806 608
rect -778 580 -740 608
rect -712 580 -674 608
rect -646 580 -608 608
rect -580 580 -542 608
rect -514 580 -476 608
rect -448 580 -410 608
rect -382 580 -344 608
rect -316 580 -278 608
rect -250 580 -212 608
rect -184 580 -146 608
rect -118 580 -80 608
rect -52 580 -14 608
rect 14 580 52 608
rect 80 580 118 608
rect 146 580 184 608
rect 212 580 250 608
rect 278 580 316 608
rect 344 580 382 608
rect 410 580 448 608
rect 476 580 514 608
rect 542 580 580 608
rect 608 580 646 608
rect 674 580 712 608
rect 740 580 778 608
rect 806 580 844 608
rect 872 580 910 608
rect 938 580 976 608
rect 1004 580 1042 608
rect 1070 580 1108 608
rect 1136 580 1174 608
rect 1202 580 1240 608
rect 1268 580 1306 608
rect 1334 580 1372 608
rect 1400 580 1438 608
rect 1466 580 1504 608
rect 1532 580 1570 608
rect 1598 580 1636 608
rect 1664 580 1702 608
rect 1730 580 1768 608
rect 1796 580 1834 608
rect 1862 580 1900 608
rect 1928 580 1966 608
rect 1994 580 2032 608
rect 2060 580 2098 608
rect 2126 580 2164 608
rect 2192 580 2230 608
rect 2258 580 2296 608
rect 2324 580 2362 608
rect 2390 580 2428 608
rect 2456 580 2494 608
rect 2522 580 2560 608
rect 2588 580 2626 608
rect 2654 580 2692 608
rect 2720 580 2758 608
rect 2786 580 2824 608
rect 2852 580 2890 608
rect 2918 580 2956 608
rect 2984 580 3022 608
rect 3050 580 3088 608
rect 3116 580 3154 608
rect 3182 580 3220 608
rect 3248 580 3286 608
rect 3314 580 3352 608
rect 3380 580 3418 608
rect 3446 580 3484 608
rect 3512 580 3550 608
rect 3578 580 3616 608
rect 3644 580 3682 608
rect 3710 580 3748 608
rect 3776 580 3814 608
rect 3842 580 3880 608
rect 3908 580 3946 608
rect 3974 580 4012 608
rect 4040 580 4078 608
rect 4106 580 4144 608
rect 4172 580 4210 608
rect 4238 580 4276 608
rect 4304 580 4342 608
rect 4370 580 4408 608
rect 4436 580 4474 608
rect 4502 580 4540 608
rect 4568 580 4573 608
rect -4573 542 4573 580
rect -4573 514 -4568 542
rect -4540 514 -4502 542
rect -4474 514 -4436 542
rect -4408 514 -4370 542
rect -4342 514 -4304 542
rect -4276 514 -4238 542
rect -4210 514 -4172 542
rect -4144 514 -4106 542
rect -4078 514 -4040 542
rect -4012 514 -3974 542
rect -3946 514 -3908 542
rect -3880 514 -3842 542
rect -3814 514 -3776 542
rect -3748 514 -3710 542
rect -3682 514 -3644 542
rect -3616 514 -3578 542
rect -3550 514 -3512 542
rect -3484 514 -3446 542
rect -3418 514 -3380 542
rect -3352 514 -3314 542
rect -3286 514 -3248 542
rect -3220 514 -3182 542
rect -3154 514 -3116 542
rect -3088 514 -3050 542
rect -3022 514 -2984 542
rect -2956 514 -2918 542
rect -2890 514 -2852 542
rect -2824 514 -2786 542
rect -2758 514 -2720 542
rect -2692 514 -2654 542
rect -2626 514 -2588 542
rect -2560 514 -2522 542
rect -2494 514 -2456 542
rect -2428 514 -2390 542
rect -2362 514 -2324 542
rect -2296 514 -2258 542
rect -2230 514 -2192 542
rect -2164 514 -2126 542
rect -2098 514 -2060 542
rect -2032 514 -1994 542
rect -1966 514 -1928 542
rect -1900 514 -1862 542
rect -1834 514 -1796 542
rect -1768 514 -1730 542
rect -1702 514 -1664 542
rect -1636 514 -1598 542
rect -1570 514 -1532 542
rect -1504 514 -1466 542
rect -1438 514 -1400 542
rect -1372 514 -1334 542
rect -1306 514 -1268 542
rect -1240 514 -1202 542
rect -1174 514 -1136 542
rect -1108 514 -1070 542
rect -1042 514 -1004 542
rect -976 514 -938 542
rect -910 514 -872 542
rect -844 514 -806 542
rect -778 514 -740 542
rect -712 514 -674 542
rect -646 514 -608 542
rect -580 514 -542 542
rect -514 514 -476 542
rect -448 514 -410 542
rect -382 514 -344 542
rect -316 514 -278 542
rect -250 514 -212 542
rect -184 514 -146 542
rect -118 514 -80 542
rect -52 514 -14 542
rect 14 514 52 542
rect 80 514 118 542
rect 146 514 184 542
rect 212 514 250 542
rect 278 514 316 542
rect 344 514 382 542
rect 410 514 448 542
rect 476 514 514 542
rect 542 514 580 542
rect 608 514 646 542
rect 674 514 712 542
rect 740 514 778 542
rect 806 514 844 542
rect 872 514 910 542
rect 938 514 976 542
rect 1004 514 1042 542
rect 1070 514 1108 542
rect 1136 514 1174 542
rect 1202 514 1240 542
rect 1268 514 1306 542
rect 1334 514 1372 542
rect 1400 514 1438 542
rect 1466 514 1504 542
rect 1532 514 1570 542
rect 1598 514 1636 542
rect 1664 514 1702 542
rect 1730 514 1768 542
rect 1796 514 1834 542
rect 1862 514 1900 542
rect 1928 514 1966 542
rect 1994 514 2032 542
rect 2060 514 2098 542
rect 2126 514 2164 542
rect 2192 514 2230 542
rect 2258 514 2296 542
rect 2324 514 2362 542
rect 2390 514 2428 542
rect 2456 514 2494 542
rect 2522 514 2560 542
rect 2588 514 2626 542
rect 2654 514 2692 542
rect 2720 514 2758 542
rect 2786 514 2824 542
rect 2852 514 2890 542
rect 2918 514 2956 542
rect 2984 514 3022 542
rect 3050 514 3088 542
rect 3116 514 3154 542
rect 3182 514 3220 542
rect 3248 514 3286 542
rect 3314 514 3352 542
rect 3380 514 3418 542
rect 3446 514 3484 542
rect 3512 514 3550 542
rect 3578 514 3616 542
rect 3644 514 3682 542
rect 3710 514 3748 542
rect 3776 514 3814 542
rect 3842 514 3880 542
rect 3908 514 3946 542
rect 3974 514 4012 542
rect 4040 514 4078 542
rect 4106 514 4144 542
rect 4172 514 4210 542
rect 4238 514 4276 542
rect 4304 514 4342 542
rect 4370 514 4408 542
rect 4436 514 4474 542
rect 4502 514 4540 542
rect 4568 514 4573 542
rect -4573 476 4573 514
rect -4573 448 -4568 476
rect -4540 448 -4502 476
rect -4474 448 -4436 476
rect -4408 448 -4370 476
rect -4342 448 -4304 476
rect -4276 448 -4238 476
rect -4210 448 -4172 476
rect -4144 448 -4106 476
rect -4078 448 -4040 476
rect -4012 448 -3974 476
rect -3946 448 -3908 476
rect -3880 448 -3842 476
rect -3814 448 -3776 476
rect -3748 448 -3710 476
rect -3682 448 -3644 476
rect -3616 448 -3578 476
rect -3550 448 -3512 476
rect -3484 448 -3446 476
rect -3418 448 -3380 476
rect -3352 448 -3314 476
rect -3286 448 -3248 476
rect -3220 448 -3182 476
rect -3154 448 -3116 476
rect -3088 448 -3050 476
rect -3022 448 -2984 476
rect -2956 448 -2918 476
rect -2890 448 -2852 476
rect -2824 448 -2786 476
rect -2758 448 -2720 476
rect -2692 448 -2654 476
rect -2626 448 -2588 476
rect -2560 448 -2522 476
rect -2494 448 -2456 476
rect -2428 448 -2390 476
rect -2362 448 -2324 476
rect -2296 448 -2258 476
rect -2230 448 -2192 476
rect -2164 448 -2126 476
rect -2098 448 -2060 476
rect -2032 448 -1994 476
rect -1966 448 -1928 476
rect -1900 448 -1862 476
rect -1834 448 -1796 476
rect -1768 448 -1730 476
rect -1702 448 -1664 476
rect -1636 448 -1598 476
rect -1570 448 -1532 476
rect -1504 448 -1466 476
rect -1438 448 -1400 476
rect -1372 448 -1334 476
rect -1306 448 -1268 476
rect -1240 448 -1202 476
rect -1174 448 -1136 476
rect -1108 448 -1070 476
rect -1042 448 -1004 476
rect -976 448 -938 476
rect -910 448 -872 476
rect -844 448 -806 476
rect -778 448 -740 476
rect -712 448 -674 476
rect -646 448 -608 476
rect -580 448 -542 476
rect -514 448 -476 476
rect -448 448 -410 476
rect -382 448 -344 476
rect -316 448 -278 476
rect -250 448 -212 476
rect -184 448 -146 476
rect -118 448 -80 476
rect -52 448 -14 476
rect 14 448 52 476
rect 80 448 118 476
rect 146 448 184 476
rect 212 448 250 476
rect 278 448 316 476
rect 344 448 382 476
rect 410 448 448 476
rect 476 448 514 476
rect 542 448 580 476
rect 608 448 646 476
rect 674 448 712 476
rect 740 448 778 476
rect 806 448 844 476
rect 872 448 910 476
rect 938 448 976 476
rect 1004 448 1042 476
rect 1070 448 1108 476
rect 1136 448 1174 476
rect 1202 448 1240 476
rect 1268 448 1306 476
rect 1334 448 1372 476
rect 1400 448 1438 476
rect 1466 448 1504 476
rect 1532 448 1570 476
rect 1598 448 1636 476
rect 1664 448 1702 476
rect 1730 448 1768 476
rect 1796 448 1834 476
rect 1862 448 1900 476
rect 1928 448 1966 476
rect 1994 448 2032 476
rect 2060 448 2098 476
rect 2126 448 2164 476
rect 2192 448 2230 476
rect 2258 448 2296 476
rect 2324 448 2362 476
rect 2390 448 2428 476
rect 2456 448 2494 476
rect 2522 448 2560 476
rect 2588 448 2626 476
rect 2654 448 2692 476
rect 2720 448 2758 476
rect 2786 448 2824 476
rect 2852 448 2890 476
rect 2918 448 2956 476
rect 2984 448 3022 476
rect 3050 448 3088 476
rect 3116 448 3154 476
rect 3182 448 3220 476
rect 3248 448 3286 476
rect 3314 448 3352 476
rect 3380 448 3418 476
rect 3446 448 3484 476
rect 3512 448 3550 476
rect 3578 448 3616 476
rect 3644 448 3682 476
rect 3710 448 3748 476
rect 3776 448 3814 476
rect 3842 448 3880 476
rect 3908 448 3946 476
rect 3974 448 4012 476
rect 4040 448 4078 476
rect 4106 448 4144 476
rect 4172 448 4210 476
rect 4238 448 4276 476
rect 4304 448 4342 476
rect 4370 448 4408 476
rect 4436 448 4474 476
rect 4502 448 4540 476
rect 4568 448 4573 476
rect -4573 410 4573 448
rect -4573 382 -4568 410
rect -4540 382 -4502 410
rect -4474 382 -4436 410
rect -4408 382 -4370 410
rect -4342 382 -4304 410
rect -4276 382 -4238 410
rect -4210 382 -4172 410
rect -4144 382 -4106 410
rect -4078 382 -4040 410
rect -4012 382 -3974 410
rect -3946 382 -3908 410
rect -3880 382 -3842 410
rect -3814 382 -3776 410
rect -3748 382 -3710 410
rect -3682 382 -3644 410
rect -3616 382 -3578 410
rect -3550 382 -3512 410
rect -3484 382 -3446 410
rect -3418 382 -3380 410
rect -3352 382 -3314 410
rect -3286 382 -3248 410
rect -3220 382 -3182 410
rect -3154 382 -3116 410
rect -3088 382 -3050 410
rect -3022 382 -2984 410
rect -2956 382 -2918 410
rect -2890 382 -2852 410
rect -2824 382 -2786 410
rect -2758 382 -2720 410
rect -2692 382 -2654 410
rect -2626 382 -2588 410
rect -2560 382 -2522 410
rect -2494 382 -2456 410
rect -2428 382 -2390 410
rect -2362 382 -2324 410
rect -2296 382 -2258 410
rect -2230 382 -2192 410
rect -2164 382 -2126 410
rect -2098 382 -2060 410
rect -2032 382 -1994 410
rect -1966 382 -1928 410
rect -1900 382 -1862 410
rect -1834 382 -1796 410
rect -1768 382 -1730 410
rect -1702 382 -1664 410
rect -1636 382 -1598 410
rect -1570 382 -1532 410
rect -1504 382 -1466 410
rect -1438 382 -1400 410
rect -1372 382 -1334 410
rect -1306 382 -1268 410
rect -1240 382 -1202 410
rect -1174 382 -1136 410
rect -1108 382 -1070 410
rect -1042 382 -1004 410
rect -976 382 -938 410
rect -910 382 -872 410
rect -844 382 -806 410
rect -778 382 -740 410
rect -712 382 -674 410
rect -646 382 -608 410
rect -580 382 -542 410
rect -514 382 -476 410
rect -448 382 -410 410
rect -382 382 -344 410
rect -316 382 -278 410
rect -250 382 -212 410
rect -184 382 -146 410
rect -118 382 -80 410
rect -52 382 -14 410
rect 14 382 52 410
rect 80 382 118 410
rect 146 382 184 410
rect 212 382 250 410
rect 278 382 316 410
rect 344 382 382 410
rect 410 382 448 410
rect 476 382 514 410
rect 542 382 580 410
rect 608 382 646 410
rect 674 382 712 410
rect 740 382 778 410
rect 806 382 844 410
rect 872 382 910 410
rect 938 382 976 410
rect 1004 382 1042 410
rect 1070 382 1108 410
rect 1136 382 1174 410
rect 1202 382 1240 410
rect 1268 382 1306 410
rect 1334 382 1372 410
rect 1400 382 1438 410
rect 1466 382 1504 410
rect 1532 382 1570 410
rect 1598 382 1636 410
rect 1664 382 1702 410
rect 1730 382 1768 410
rect 1796 382 1834 410
rect 1862 382 1900 410
rect 1928 382 1966 410
rect 1994 382 2032 410
rect 2060 382 2098 410
rect 2126 382 2164 410
rect 2192 382 2230 410
rect 2258 382 2296 410
rect 2324 382 2362 410
rect 2390 382 2428 410
rect 2456 382 2494 410
rect 2522 382 2560 410
rect 2588 382 2626 410
rect 2654 382 2692 410
rect 2720 382 2758 410
rect 2786 382 2824 410
rect 2852 382 2890 410
rect 2918 382 2956 410
rect 2984 382 3022 410
rect 3050 382 3088 410
rect 3116 382 3154 410
rect 3182 382 3220 410
rect 3248 382 3286 410
rect 3314 382 3352 410
rect 3380 382 3418 410
rect 3446 382 3484 410
rect 3512 382 3550 410
rect 3578 382 3616 410
rect 3644 382 3682 410
rect 3710 382 3748 410
rect 3776 382 3814 410
rect 3842 382 3880 410
rect 3908 382 3946 410
rect 3974 382 4012 410
rect 4040 382 4078 410
rect 4106 382 4144 410
rect 4172 382 4210 410
rect 4238 382 4276 410
rect 4304 382 4342 410
rect 4370 382 4408 410
rect 4436 382 4474 410
rect 4502 382 4540 410
rect 4568 382 4573 410
rect -4573 344 4573 382
rect -4573 316 -4568 344
rect -4540 316 -4502 344
rect -4474 316 -4436 344
rect -4408 316 -4370 344
rect -4342 316 -4304 344
rect -4276 316 -4238 344
rect -4210 316 -4172 344
rect -4144 316 -4106 344
rect -4078 316 -4040 344
rect -4012 316 -3974 344
rect -3946 316 -3908 344
rect -3880 316 -3842 344
rect -3814 316 -3776 344
rect -3748 316 -3710 344
rect -3682 316 -3644 344
rect -3616 316 -3578 344
rect -3550 316 -3512 344
rect -3484 316 -3446 344
rect -3418 316 -3380 344
rect -3352 316 -3314 344
rect -3286 316 -3248 344
rect -3220 316 -3182 344
rect -3154 316 -3116 344
rect -3088 316 -3050 344
rect -3022 316 -2984 344
rect -2956 316 -2918 344
rect -2890 316 -2852 344
rect -2824 316 -2786 344
rect -2758 316 -2720 344
rect -2692 316 -2654 344
rect -2626 316 -2588 344
rect -2560 316 -2522 344
rect -2494 316 -2456 344
rect -2428 316 -2390 344
rect -2362 316 -2324 344
rect -2296 316 -2258 344
rect -2230 316 -2192 344
rect -2164 316 -2126 344
rect -2098 316 -2060 344
rect -2032 316 -1994 344
rect -1966 316 -1928 344
rect -1900 316 -1862 344
rect -1834 316 -1796 344
rect -1768 316 -1730 344
rect -1702 316 -1664 344
rect -1636 316 -1598 344
rect -1570 316 -1532 344
rect -1504 316 -1466 344
rect -1438 316 -1400 344
rect -1372 316 -1334 344
rect -1306 316 -1268 344
rect -1240 316 -1202 344
rect -1174 316 -1136 344
rect -1108 316 -1070 344
rect -1042 316 -1004 344
rect -976 316 -938 344
rect -910 316 -872 344
rect -844 316 -806 344
rect -778 316 -740 344
rect -712 316 -674 344
rect -646 316 -608 344
rect -580 316 -542 344
rect -514 316 -476 344
rect -448 316 -410 344
rect -382 316 -344 344
rect -316 316 -278 344
rect -250 316 -212 344
rect -184 316 -146 344
rect -118 316 -80 344
rect -52 316 -14 344
rect 14 316 52 344
rect 80 316 118 344
rect 146 316 184 344
rect 212 316 250 344
rect 278 316 316 344
rect 344 316 382 344
rect 410 316 448 344
rect 476 316 514 344
rect 542 316 580 344
rect 608 316 646 344
rect 674 316 712 344
rect 740 316 778 344
rect 806 316 844 344
rect 872 316 910 344
rect 938 316 976 344
rect 1004 316 1042 344
rect 1070 316 1108 344
rect 1136 316 1174 344
rect 1202 316 1240 344
rect 1268 316 1306 344
rect 1334 316 1372 344
rect 1400 316 1438 344
rect 1466 316 1504 344
rect 1532 316 1570 344
rect 1598 316 1636 344
rect 1664 316 1702 344
rect 1730 316 1768 344
rect 1796 316 1834 344
rect 1862 316 1900 344
rect 1928 316 1966 344
rect 1994 316 2032 344
rect 2060 316 2098 344
rect 2126 316 2164 344
rect 2192 316 2230 344
rect 2258 316 2296 344
rect 2324 316 2362 344
rect 2390 316 2428 344
rect 2456 316 2494 344
rect 2522 316 2560 344
rect 2588 316 2626 344
rect 2654 316 2692 344
rect 2720 316 2758 344
rect 2786 316 2824 344
rect 2852 316 2890 344
rect 2918 316 2956 344
rect 2984 316 3022 344
rect 3050 316 3088 344
rect 3116 316 3154 344
rect 3182 316 3220 344
rect 3248 316 3286 344
rect 3314 316 3352 344
rect 3380 316 3418 344
rect 3446 316 3484 344
rect 3512 316 3550 344
rect 3578 316 3616 344
rect 3644 316 3682 344
rect 3710 316 3748 344
rect 3776 316 3814 344
rect 3842 316 3880 344
rect 3908 316 3946 344
rect 3974 316 4012 344
rect 4040 316 4078 344
rect 4106 316 4144 344
rect 4172 316 4210 344
rect 4238 316 4276 344
rect 4304 316 4342 344
rect 4370 316 4408 344
rect 4436 316 4474 344
rect 4502 316 4540 344
rect 4568 316 4573 344
rect -4573 278 4573 316
rect -4573 250 -4568 278
rect -4540 250 -4502 278
rect -4474 250 -4436 278
rect -4408 250 -4370 278
rect -4342 250 -4304 278
rect -4276 250 -4238 278
rect -4210 250 -4172 278
rect -4144 250 -4106 278
rect -4078 250 -4040 278
rect -4012 250 -3974 278
rect -3946 250 -3908 278
rect -3880 250 -3842 278
rect -3814 250 -3776 278
rect -3748 250 -3710 278
rect -3682 250 -3644 278
rect -3616 250 -3578 278
rect -3550 250 -3512 278
rect -3484 250 -3446 278
rect -3418 250 -3380 278
rect -3352 250 -3314 278
rect -3286 250 -3248 278
rect -3220 250 -3182 278
rect -3154 250 -3116 278
rect -3088 250 -3050 278
rect -3022 250 -2984 278
rect -2956 250 -2918 278
rect -2890 250 -2852 278
rect -2824 250 -2786 278
rect -2758 250 -2720 278
rect -2692 250 -2654 278
rect -2626 250 -2588 278
rect -2560 250 -2522 278
rect -2494 250 -2456 278
rect -2428 250 -2390 278
rect -2362 250 -2324 278
rect -2296 250 -2258 278
rect -2230 250 -2192 278
rect -2164 250 -2126 278
rect -2098 250 -2060 278
rect -2032 250 -1994 278
rect -1966 250 -1928 278
rect -1900 250 -1862 278
rect -1834 250 -1796 278
rect -1768 250 -1730 278
rect -1702 250 -1664 278
rect -1636 250 -1598 278
rect -1570 250 -1532 278
rect -1504 250 -1466 278
rect -1438 250 -1400 278
rect -1372 250 -1334 278
rect -1306 250 -1268 278
rect -1240 250 -1202 278
rect -1174 250 -1136 278
rect -1108 250 -1070 278
rect -1042 250 -1004 278
rect -976 250 -938 278
rect -910 250 -872 278
rect -844 250 -806 278
rect -778 250 -740 278
rect -712 250 -674 278
rect -646 250 -608 278
rect -580 250 -542 278
rect -514 250 -476 278
rect -448 250 -410 278
rect -382 250 -344 278
rect -316 250 -278 278
rect -250 250 -212 278
rect -184 250 -146 278
rect -118 250 -80 278
rect -52 250 -14 278
rect 14 250 52 278
rect 80 250 118 278
rect 146 250 184 278
rect 212 250 250 278
rect 278 250 316 278
rect 344 250 382 278
rect 410 250 448 278
rect 476 250 514 278
rect 542 250 580 278
rect 608 250 646 278
rect 674 250 712 278
rect 740 250 778 278
rect 806 250 844 278
rect 872 250 910 278
rect 938 250 976 278
rect 1004 250 1042 278
rect 1070 250 1108 278
rect 1136 250 1174 278
rect 1202 250 1240 278
rect 1268 250 1306 278
rect 1334 250 1372 278
rect 1400 250 1438 278
rect 1466 250 1504 278
rect 1532 250 1570 278
rect 1598 250 1636 278
rect 1664 250 1702 278
rect 1730 250 1768 278
rect 1796 250 1834 278
rect 1862 250 1900 278
rect 1928 250 1966 278
rect 1994 250 2032 278
rect 2060 250 2098 278
rect 2126 250 2164 278
rect 2192 250 2230 278
rect 2258 250 2296 278
rect 2324 250 2362 278
rect 2390 250 2428 278
rect 2456 250 2494 278
rect 2522 250 2560 278
rect 2588 250 2626 278
rect 2654 250 2692 278
rect 2720 250 2758 278
rect 2786 250 2824 278
rect 2852 250 2890 278
rect 2918 250 2956 278
rect 2984 250 3022 278
rect 3050 250 3088 278
rect 3116 250 3154 278
rect 3182 250 3220 278
rect 3248 250 3286 278
rect 3314 250 3352 278
rect 3380 250 3418 278
rect 3446 250 3484 278
rect 3512 250 3550 278
rect 3578 250 3616 278
rect 3644 250 3682 278
rect 3710 250 3748 278
rect 3776 250 3814 278
rect 3842 250 3880 278
rect 3908 250 3946 278
rect 3974 250 4012 278
rect 4040 250 4078 278
rect 4106 250 4144 278
rect 4172 250 4210 278
rect 4238 250 4276 278
rect 4304 250 4342 278
rect 4370 250 4408 278
rect 4436 250 4474 278
rect 4502 250 4540 278
rect 4568 250 4573 278
rect -4573 212 4573 250
rect -4573 184 -4568 212
rect -4540 184 -4502 212
rect -4474 184 -4436 212
rect -4408 184 -4370 212
rect -4342 184 -4304 212
rect -4276 184 -4238 212
rect -4210 184 -4172 212
rect -4144 184 -4106 212
rect -4078 184 -4040 212
rect -4012 184 -3974 212
rect -3946 184 -3908 212
rect -3880 184 -3842 212
rect -3814 184 -3776 212
rect -3748 184 -3710 212
rect -3682 184 -3644 212
rect -3616 184 -3578 212
rect -3550 184 -3512 212
rect -3484 184 -3446 212
rect -3418 184 -3380 212
rect -3352 184 -3314 212
rect -3286 184 -3248 212
rect -3220 184 -3182 212
rect -3154 184 -3116 212
rect -3088 184 -3050 212
rect -3022 184 -2984 212
rect -2956 184 -2918 212
rect -2890 184 -2852 212
rect -2824 184 -2786 212
rect -2758 184 -2720 212
rect -2692 184 -2654 212
rect -2626 184 -2588 212
rect -2560 184 -2522 212
rect -2494 184 -2456 212
rect -2428 184 -2390 212
rect -2362 184 -2324 212
rect -2296 184 -2258 212
rect -2230 184 -2192 212
rect -2164 184 -2126 212
rect -2098 184 -2060 212
rect -2032 184 -1994 212
rect -1966 184 -1928 212
rect -1900 184 -1862 212
rect -1834 184 -1796 212
rect -1768 184 -1730 212
rect -1702 184 -1664 212
rect -1636 184 -1598 212
rect -1570 184 -1532 212
rect -1504 184 -1466 212
rect -1438 184 -1400 212
rect -1372 184 -1334 212
rect -1306 184 -1268 212
rect -1240 184 -1202 212
rect -1174 184 -1136 212
rect -1108 184 -1070 212
rect -1042 184 -1004 212
rect -976 184 -938 212
rect -910 184 -872 212
rect -844 184 -806 212
rect -778 184 -740 212
rect -712 184 -674 212
rect -646 184 -608 212
rect -580 184 -542 212
rect -514 184 -476 212
rect -448 184 -410 212
rect -382 184 -344 212
rect -316 184 -278 212
rect -250 184 -212 212
rect -184 184 -146 212
rect -118 184 -80 212
rect -52 184 -14 212
rect 14 184 52 212
rect 80 184 118 212
rect 146 184 184 212
rect 212 184 250 212
rect 278 184 316 212
rect 344 184 382 212
rect 410 184 448 212
rect 476 184 514 212
rect 542 184 580 212
rect 608 184 646 212
rect 674 184 712 212
rect 740 184 778 212
rect 806 184 844 212
rect 872 184 910 212
rect 938 184 976 212
rect 1004 184 1042 212
rect 1070 184 1108 212
rect 1136 184 1174 212
rect 1202 184 1240 212
rect 1268 184 1306 212
rect 1334 184 1372 212
rect 1400 184 1438 212
rect 1466 184 1504 212
rect 1532 184 1570 212
rect 1598 184 1636 212
rect 1664 184 1702 212
rect 1730 184 1768 212
rect 1796 184 1834 212
rect 1862 184 1900 212
rect 1928 184 1966 212
rect 1994 184 2032 212
rect 2060 184 2098 212
rect 2126 184 2164 212
rect 2192 184 2230 212
rect 2258 184 2296 212
rect 2324 184 2362 212
rect 2390 184 2428 212
rect 2456 184 2494 212
rect 2522 184 2560 212
rect 2588 184 2626 212
rect 2654 184 2692 212
rect 2720 184 2758 212
rect 2786 184 2824 212
rect 2852 184 2890 212
rect 2918 184 2956 212
rect 2984 184 3022 212
rect 3050 184 3088 212
rect 3116 184 3154 212
rect 3182 184 3220 212
rect 3248 184 3286 212
rect 3314 184 3352 212
rect 3380 184 3418 212
rect 3446 184 3484 212
rect 3512 184 3550 212
rect 3578 184 3616 212
rect 3644 184 3682 212
rect 3710 184 3748 212
rect 3776 184 3814 212
rect 3842 184 3880 212
rect 3908 184 3946 212
rect 3974 184 4012 212
rect 4040 184 4078 212
rect 4106 184 4144 212
rect 4172 184 4210 212
rect 4238 184 4276 212
rect 4304 184 4342 212
rect 4370 184 4408 212
rect 4436 184 4474 212
rect 4502 184 4540 212
rect 4568 184 4573 212
rect -4573 146 4573 184
rect -4573 118 -4568 146
rect -4540 118 -4502 146
rect -4474 118 -4436 146
rect -4408 118 -4370 146
rect -4342 118 -4304 146
rect -4276 118 -4238 146
rect -4210 118 -4172 146
rect -4144 118 -4106 146
rect -4078 118 -4040 146
rect -4012 118 -3974 146
rect -3946 118 -3908 146
rect -3880 118 -3842 146
rect -3814 118 -3776 146
rect -3748 118 -3710 146
rect -3682 118 -3644 146
rect -3616 118 -3578 146
rect -3550 118 -3512 146
rect -3484 118 -3446 146
rect -3418 118 -3380 146
rect -3352 118 -3314 146
rect -3286 118 -3248 146
rect -3220 118 -3182 146
rect -3154 118 -3116 146
rect -3088 118 -3050 146
rect -3022 118 -2984 146
rect -2956 118 -2918 146
rect -2890 118 -2852 146
rect -2824 118 -2786 146
rect -2758 118 -2720 146
rect -2692 118 -2654 146
rect -2626 118 -2588 146
rect -2560 118 -2522 146
rect -2494 118 -2456 146
rect -2428 118 -2390 146
rect -2362 118 -2324 146
rect -2296 118 -2258 146
rect -2230 118 -2192 146
rect -2164 118 -2126 146
rect -2098 118 -2060 146
rect -2032 118 -1994 146
rect -1966 118 -1928 146
rect -1900 118 -1862 146
rect -1834 118 -1796 146
rect -1768 118 -1730 146
rect -1702 118 -1664 146
rect -1636 118 -1598 146
rect -1570 118 -1532 146
rect -1504 118 -1466 146
rect -1438 118 -1400 146
rect -1372 118 -1334 146
rect -1306 118 -1268 146
rect -1240 118 -1202 146
rect -1174 118 -1136 146
rect -1108 118 -1070 146
rect -1042 118 -1004 146
rect -976 118 -938 146
rect -910 118 -872 146
rect -844 118 -806 146
rect -778 118 -740 146
rect -712 118 -674 146
rect -646 118 -608 146
rect -580 118 -542 146
rect -514 118 -476 146
rect -448 118 -410 146
rect -382 118 -344 146
rect -316 118 -278 146
rect -250 118 -212 146
rect -184 118 -146 146
rect -118 118 -80 146
rect -52 118 -14 146
rect 14 118 52 146
rect 80 118 118 146
rect 146 118 184 146
rect 212 118 250 146
rect 278 118 316 146
rect 344 118 382 146
rect 410 118 448 146
rect 476 118 514 146
rect 542 118 580 146
rect 608 118 646 146
rect 674 118 712 146
rect 740 118 778 146
rect 806 118 844 146
rect 872 118 910 146
rect 938 118 976 146
rect 1004 118 1042 146
rect 1070 118 1108 146
rect 1136 118 1174 146
rect 1202 118 1240 146
rect 1268 118 1306 146
rect 1334 118 1372 146
rect 1400 118 1438 146
rect 1466 118 1504 146
rect 1532 118 1570 146
rect 1598 118 1636 146
rect 1664 118 1702 146
rect 1730 118 1768 146
rect 1796 118 1834 146
rect 1862 118 1900 146
rect 1928 118 1966 146
rect 1994 118 2032 146
rect 2060 118 2098 146
rect 2126 118 2164 146
rect 2192 118 2230 146
rect 2258 118 2296 146
rect 2324 118 2362 146
rect 2390 118 2428 146
rect 2456 118 2494 146
rect 2522 118 2560 146
rect 2588 118 2626 146
rect 2654 118 2692 146
rect 2720 118 2758 146
rect 2786 118 2824 146
rect 2852 118 2890 146
rect 2918 118 2956 146
rect 2984 118 3022 146
rect 3050 118 3088 146
rect 3116 118 3154 146
rect 3182 118 3220 146
rect 3248 118 3286 146
rect 3314 118 3352 146
rect 3380 118 3418 146
rect 3446 118 3484 146
rect 3512 118 3550 146
rect 3578 118 3616 146
rect 3644 118 3682 146
rect 3710 118 3748 146
rect 3776 118 3814 146
rect 3842 118 3880 146
rect 3908 118 3946 146
rect 3974 118 4012 146
rect 4040 118 4078 146
rect 4106 118 4144 146
rect 4172 118 4210 146
rect 4238 118 4276 146
rect 4304 118 4342 146
rect 4370 118 4408 146
rect 4436 118 4474 146
rect 4502 118 4540 146
rect 4568 118 4573 146
rect -4573 80 4573 118
rect -4573 52 -4568 80
rect -4540 52 -4502 80
rect -4474 52 -4436 80
rect -4408 52 -4370 80
rect -4342 52 -4304 80
rect -4276 52 -4238 80
rect -4210 52 -4172 80
rect -4144 52 -4106 80
rect -4078 52 -4040 80
rect -4012 52 -3974 80
rect -3946 52 -3908 80
rect -3880 52 -3842 80
rect -3814 52 -3776 80
rect -3748 52 -3710 80
rect -3682 52 -3644 80
rect -3616 52 -3578 80
rect -3550 52 -3512 80
rect -3484 52 -3446 80
rect -3418 52 -3380 80
rect -3352 52 -3314 80
rect -3286 52 -3248 80
rect -3220 52 -3182 80
rect -3154 52 -3116 80
rect -3088 52 -3050 80
rect -3022 52 -2984 80
rect -2956 52 -2918 80
rect -2890 52 -2852 80
rect -2824 52 -2786 80
rect -2758 52 -2720 80
rect -2692 52 -2654 80
rect -2626 52 -2588 80
rect -2560 52 -2522 80
rect -2494 52 -2456 80
rect -2428 52 -2390 80
rect -2362 52 -2324 80
rect -2296 52 -2258 80
rect -2230 52 -2192 80
rect -2164 52 -2126 80
rect -2098 52 -2060 80
rect -2032 52 -1994 80
rect -1966 52 -1928 80
rect -1900 52 -1862 80
rect -1834 52 -1796 80
rect -1768 52 -1730 80
rect -1702 52 -1664 80
rect -1636 52 -1598 80
rect -1570 52 -1532 80
rect -1504 52 -1466 80
rect -1438 52 -1400 80
rect -1372 52 -1334 80
rect -1306 52 -1268 80
rect -1240 52 -1202 80
rect -1174 52 -1136 80
rect -1108 52 -1070 80
rect -1042 52 -1004 80
rect -976 52 -938 80
rect -910 52 -872 80
rect -844 52 -806 80
rect -778 52 -740 80
rect -712 52 -674 80
rect -646 52 -608 80
rect -580 52 -542 80
rect -514 52 -476 80
rect -448 52 -410 80
rect -382 52 -344 80
rect -316 52 -278 80
rect -250 52 -212 80
rect -184 52 -146 80
rect -118 52 -80 80
rect -52 52 -14 80
rect 14 52 52 80
rect 80 52 118 80
rect 146 52 184 80
rect 212 52 250 80
rect 278 52 316 80
rect 344 52 382 80
rect 410 52 448 80
rect 476 52 514 80
rect 542 52 580 80
rect 608 52 646 80
rect 674 52 712 80
rect 740 52 778 80
rect 806 52 844 80
rect 872 52 910 80
rect 938 52 976 80
rect 1004 52 1042 80
rect 1070 52 1108 80
rect 1136 52 1174 80
rect 1202 52 1240 80
rect 1268 52 1306 80
rect 1334 52 1372 80
rect 1400 52 1438 80
rect 1466 52 1504 80
rect 1532 52 1570 80
rect 1598 52 1636 80
rect 1664 52 1702 80
rect 1730 52 1768 80
rect 1796 52 1834 80
rect 1862 52 1900 80
rect 1928 52 1966 80
rect 1994 52 2032 80
rect 2060 52 2098 80
rect 2126 52 2164 80
rect 2192 52 2230 80
rect 2258 52 2296 80
rect 2324 52 2362 80
rect 2390 52 2428 80
rect 2456 52 2494 80
rect 2522 52 2560 80
rect 2588 52 2626 80
rect 2654 52 2692 80
rect 2720 52 2758 80
rect 2786 52 2824 80
rect 2852 52 2890 80
rect 2918 52 2956 80
rect 2984 52 3022 80
rect 3050 52 3088 80
rect 3116 52 3154 80
rect 3182 52 3220 80
rect 3248 52 3286 80
rect 3314 52 3352 80
rect 3380 52 3418 80
rect 3446 52 3484 80
rect 3512 52 3550 80
rect 3578 52 3616 80
rect 3644 52 3682 80
rect 3710 52 3748 80
rect 3776 52 3814 80
rect 3842 52 3880 80
rect 3908 52 3946 80
rect 3974 52 4012 80
rect 4040 52 4078 80
rect 4106 52 4144 80
rect 4172 52 4210 80
rect 4238 52 4276 80
rect 4304 52 4342 80
rect 4370 52 4408 80
rect 4436 52 4474 80
rect 4502 52 4540 80
rect 4568 52 4573 80
rect -4573 14 4573 52
rect -4573 -14 -4568 14
rect -4540 -14 -4502 14
rect -4474 -14 -4436 14
rect -4408 -14 -4370 14
rect -4342 -14 -4304 14
rect -4276 -14 -4238 14
rect -4210 -14 -4172 14
rect -4144 -14 -4106 14
rect -4078 -14 -4040 14
rect -4012 -14 -3974 14
rect -3946 -14 -3908 14
rect -3880 -14 -3842 14
rect -3814 -14 -3776 14
rect -3748 -14 -3710 14
rect -3682 -14 -3644 14
rect -3616 -14 -3578 14
rect -3550 -14 -3512 14
rect -3484 -14 -3446 14
rect -3418 -14 -3380 14
rect -3352 -14 -3314 14
rect -3286 -14 -3248 14
rect -3220 -14 -3182 14
rect -3154 -14 -3116 14
rect -3088 -14 -3050 14
rect -3022 -14 -2984 14
rect -2956 -14 -2918 14
rect -2890 -14 -2852 14
rect -2824 -14 -2786 14
rect -2758 -14 -2720 14
rect -2692 -14 -2654 14
rect -2626 -14 -2588 14
rect -2560 -14 -2522 14
rect -2494 -14 -2456 14
rect -2428 -14 -2390 14
rect -2362 -14 -2324 14
rect -2296 -14 -2258 14
rect -2230 -14 -2192 14
rect -2164 -14 -2126 14
rect -2098 -14 -2060 14
rect -2032 -14 -1994 14
rect -1966 -14 -1928 14
rect -1900 -14 -1862 14
rect -1834 -14 -1796 14
rect -1768 -14 -1730 14
rect -1702 -14 -1664 14
rect -1636 -14 -1598 14
rect -1570 -14 -1532 14
rect -1504 -14 -1466 14
rect -1438 -14 -1400 14
rect -1372 -14 -1334 14
rect -1306 -14 -1268 14
rect -1240 -14 -1202 14
rect -1174 -14 -1136 14
rect -1108 -14 -1070 14
rect -1042 -14 -1004 14
rect -976 -14 -938 14
rect -910 -14 -872 14
rect -844 -14 -806 14
rect -778 -14 -740 14
rect -712 -14 -674 14
rect -646 -14 -608 14
rect -580 -14 -542 14
rect -514 -14 -476 14
rect -448 -14 -410 14
rect -382 -14 -344 14
rect -316 -14 -278 14
rect -250 -14 -212 14
rect -184 -14 -146 14
rect -118 -14 -80 14
rect -52 -14 -14 14
rect 14 -14 52 14
rect 80 -14 118 14
rect 146 -14 184 14
rect 212 -14 250 14
rect 278 -14 316 14
rect 344 -14 382 14
rect 410 -14 448 14
rect 476 -14 514 14
rect 542 -14 580 14
rect 608 -14 646 14
rect 674 -14 712 14
rect 740 -14 778 14
rect 806 -14 844 14
rect 872 -14 910 14
rect 938 -14 976 14
rect 1004 -14 1042 14
rect 1070 -14 1108 14
rect 1136 -14 1174 14
rect 1202 -14 1240 14
rect 1268 -14 1306 14
rect 1334 -14 1372 14
rect 1400 -14 1438 14
rect 1466 -14 1504 14
rect 1532 -14 1570 14
rect 1598 -14 1636 14
rect 1664 -14 1702 14
rect 1730 -14 1768 14
rect 1796 -14 1834 14
rect 1862 -14 1900 14
rect 1928 -14 1966 14
rect 1994 -14 2032 14
rect 2060 -14 2098 14
rect 2126 -14 2164 14
rect 2192 -14 2230 14
rect 2258 -14 2296 14
rect 2324 -14 2362 14
rect 2390 -14 2428 14
rect 2456 -14 2494 14
rect 2522 -14 2560 14
rect 2588 -14 2626 14
rect 2654 -14 2692 14
rect 2720 -14 2758 14
rect 2786 -14 2824 14
rect 2852 -14 2890 14
rect 2918 -14 2956 14
rect 2984 -14 3022 14
rect 3050 -14 3088 14
rect 3116 -14 3154 14
rect 3182 -14 3220 14
rect 3248 -14 3286 14
rect 3314 -14 3352 14
rect 3380 -14 3418 14
rect 3446 -14 3484 14
rect 3512 -14 3550 14
rect 3578 -14 3616 14
rect 3644 -14 3682 14
rect 3710 -14 3748 14
rect 3776 -14 3814 14
rect 3842 -14 3880 14
rect 3908 -14 3946 14
rect 3974 -14 4012 14
rect 4040 -14 4078 14
rect 4106 -14 4144 14
rect 4172 -14 4210 14
rect 4238 -14 4276 14
rect 4304 -14 4342 14
rect 4370 -14 4408 14
rect 4436 -14 4474 14
rect 4502 -14 4540 14
rect 4568 -14 4573 14
rect -4573 -52 4573 -14
rect -4573 -80 -4568 -52
rect -4540 -80 -4502 -52
rect -4474 -80 -4436 -52
rect -4408 -80 -4370 -52
rect -4342 -80 -4304 -52
rect -4276 -80 -4238 -52
rect -4210 -80 -4172 -52
rect -4144 -80 -4106 -52
rect -4078 -80 -4040 -52
rect -4012 -80 -3974 -52
rect -3946 -80 -3908 -52
rect -3880 -80 -3842 -52
rect -3814 -80 -3776 -52
rect -3748 -80 -3710 -52
rect -3682 -80 -3644 -52
rect -3616 -80 -3578 -52
rect -3550 -80 -3512 -52
rect -3484 -80 -3446 -52
rect -3418 -80 -3380 -52
rect -3352 -80 -3314 -52
rect -3286 -80 -3248 -52
rect -3220 -80 -3182 -52
rect -3154 -80 -3116 -52
rect -3088 -80 -3050 -52
rect -3022 -80 -2984 -52
rect -2956 -80 -2918 -52
rect -2890 -80 -2852 -52
rect -2824 -80 -2786 -52
rect -2758 -80 -2720 -52
rect -2692 -80 -2654 -52
rect -2626 -80 -2588 -52
rect -2560 -80 -2522 -52
rect -2494 -80 -2456 -52
rect -2428 -80 -2390 -52
rect -2362 -80 -2324 -52
rect -2296 -80 -2258 -52
rect -2230 -80 -2192 -52
rect -2164 -80 -2126 -52
rect -2098 -80 -2060 -52
rect -2032 -80 -1994 -52
rect -1966 -80 -1928 -52
rect -1900 -80 -1862 -52
rect -1834 -80 -1796 -52
rect -1768 -80 -1730 -52
rect -1702 -80 -1664 -52
rect -1636 -80 -1598 -52
rect -1570 -80 -1532 -52
rect -1504 -80 -1466 -52
rect -1438 -80 -1400 -52
rect -1372 -80 -1334 -52
rect -1306 -80 -1268 -52
rect -1240 -80 -1202 -52
rect -1174 -80 -1136 -52
rect -1108 -80 -1070 -52
rect -1042 -80 -1004 -52
rect -976 -80 -938 -52
rect -910 -80 -872 -52
rect -844 -80 -806 -52
rect -778 -80 -740 -52
rect -712 -80 -674 -52
rect -646 -80 -608 -52
rect -580 -80 -542 -52
rect -514 -80 -476 -52
rect -448 -80 -410 -52
rect -382 -80 -344 -52
rect -316 -80 -278 -52
rect -250 -80 -212 -52
rect -184 -80 -146 -52
rect -118 -80 -80 -52
rect -52 -80 -14 -52
rect 14 -80 52 -52
rect 80 -80 118 -52
rect 146 -80 184 -52
rect 212 -80 250 -52
rect 278 -80 316 -52
rect 344 -80 382 -52
rect 410 -80 448 -52
rect 476 -80 514 -52
rect 542 -80 580 -52
rect 608 -80 646 -52
rect 674 -80 712 -52
rect 740 -80 778 -52
rect 806 -80 844 -52
rect 872 -80 910 -52
rect 938 -80 976 -52
rect 1004 -80 1042 -52
rect 1070 -80 1108 -52
rect 1136 -80 1174 -52
rect 1202 -80 1240 -52
rect 1268 -80 1306 -52
rect 1334 -80 1372 -52
rect 1400 -80 1438 -52
rect 1466 -80 1504 -52
rect 1532 -80 1570 -52
rect 1598 -80 1636 -52
rect 1664 -80 1702 -52
rect 1730 -80 1768 -52
rect 1796 -80 1834 -52
rect 1862 -80 1900 -52
rect 1928 -80 1966 -52
rect 1994 -80 2032 -52
rect 2060 -80 2098 -52
rect 2126 -80 2164 -52
rect 2192 -80 2230 -52
rect 2258 -80 2296 -52
rect 2324 -80 2362 -52
rect 2390 -80 2428 -52
rect 2456 -80 2494 -52
rect 2522 -80 2560 -52
rect 2588 -80 2626 -52
rect 2654 -80 2692 -52
rect 2720 -80 2758 -52
rect 2786 -80 2824 -52
rect 2852 -80 2890 -52
rect 2918 -80 2956 -52
rect 2984 -80 3022 -52
rect 3050 -80 3088 -52
rect 3116 -80 3154 -52
rect 3182 -80 3220 -52
rect 3248 -80 3286 -52
rect 3314 -80 3352 -52
rect 3380 -80 3418 -52
rect 3446 -80 3484 -52
rect 3512 -80 3550 -52
rect 3578 -80 3616 -52
rect 3644 -80 3682 -52
rect 3710 -80 3748 -52
rect 3776 -80 3814 -52
rect 3842 -80 3880 -52
rect 3908 -80 3946 -52
rect 3974 -80 4012 -52
rect 4040 -80 4078 -52
rect 4106 -80 4144 -52
rect 4172 -80 4210 -52
rect 4238 -80 4276 -52
rect 4304 -80 4342 -52
rect 4370 -80 4408 -52
rect 4436 -80 4474 -52
rect 4502 -80 4540 -52
rect 4568 -80 4573 -52
rect -4573 -118 4573 -80
rect -4573 -146 -4568 -118
rect -4540 -146 -4502 -118
rect -4474 -146 -4436 -118
rect -4408 -146 -4370 -118
rect -4342 -146 -4304 -118
rect -4276 -146 -4238 -118
rect -4210 -146 -4172 -118
rect -4144 -146 -4106 -118
rect -4078 -146 -4040 -118
rect -4012 -146 -3974 -118
rect -3946 -146 -3908 -118
rect -3880 -146 -3842 -118
rect -3814 -146 -3776 -118
rect -3748 -146 -3710 -118
rect -3682 -146 -3644 -118
rect -3616 -146 -3578 -118
rect -3550 -146 -3512 -118
rect -3484 -146 -3446 -118
rect -3418 -146 -3380 -118
rect -3352 -146 -3314 -118
rect -3286 -146 -3248 -118
rect -3220 -146 -3182 -118
rect -3154 -146 -3116 -118
rect -3088 -146 -3050 -118
rect -3022 -146 -2984 -118
rect -2956 -146 -2918 -118
rect -2890 -146 -2852 -118
rect -2824 -146 -2786 -118
rect -2758 -146 -2720 -118
rect -2692 -146 -2654 -118
rect -2626 -146 -2588 -118
rect -2560 -146 -2522 -118
rect -2494 -146 -2456 -118
rect -2428 -146 -2390 -118
rect -2362 -146 -2324 -118
rect -2296 -146 -2258 -118
rect -2230 -146 -2192 -118
rect -2164 -146 -2126 -118
rect -2098 -146 -2060 -118
rect -2032 -146 -1994 -118
rect -1966 -146 -1928 -118
rect -1900 -146 -1862 -118
rect -1834 -146 -1796 -118
rect -1768 -146 -1730 -118
rect -1702 -146 -1664 -118
rect -1636 -146 -1598 -118
rect -1570 -146 -1532 -118
rect -1504 -146 -1466 -118
rect -1438 -146 -1400 -118
rect -1372 -146 -1334 -118
rect -1306 -146 -1268 -118
rect -1240 -146 -1202 -118
rect -1174 -146 -1136 -118
rect -1108 -146 -1070 -118
rect -1042 -146 -1004 -118
rect -976 -146 -938 -118
rect -910 -146 -872 -118
rect -844 -146 -806 -118
rect -778 -146 -740 -118
rect -712 -146 -674 -118
rect -646 -146 -608 -118
rect -580 -146 -542 -118
rect -514 -146 -476 -118
rect -448 -146 -410 -118
rect -382 -146 -344 -118
rect -316 -146 -278 -118
rect -250 -146 -212 -118
rect -184 -146 -146 -118
rect -118 -146 -80 -118
rect -52 -146 -14 -118
rect 14 -146 52 -118
rect 80 -146 118 -118
rect 146 -146 184 -118
rect 212 -146 250 -118
rect 278 -146 316 -118
rect 344 -146 382 -118
rect 410 -146 448 -118
rect 476 -146 514 -118
rect 542 -146 580 -118
rect 608 -146 646 -118
rect 674 -146 712 -118
rect 740 -146 778 -118
rect 806 -146 844 -118
rect 872 -146 910 -118
rect 938 -146 976 -118
rect 1004 -146 1042 -118
rect 1070 -146 1108 -118
rect 1136 -146 1174 -118
rect 1202 -146 1240 -118
rect 1268 -146 1306 -118
rect 1334 -146 1372 -118
rect 1400 -146 1438 -118
rect 1466 -146 1504 -118
rect 1532 -146 1570 -118
rect 1598 -146 1636 -118
rect 1664 -146 1702 -118
rect 1730 -146 1768 -118
rect 1796 -146 1834 -118
rect 1862 -146 1900 -118
rect 1928 -146 1966 -118
rect 1994 -146 2032 -118
rect 2060 -146 2098 -118
rect 2126 -146 2164 -118
rect 2192 -146 2230 -118
rect 2258 -146 2296 -118
rect 2324 -146 2362 -118
rect 2390 -146 2428 -118
rect 2456 -146 2494 -118
rect 2522 -146 2560 -118
rect 2588 -146 2626 -118
rect 2654 -146 2692 -118
rect 2720 -146 2758 -118
rect 2786 -146 2824 -118
rect 2852 -146 2890 -118
rect 2918 -146 2956 -118
rect 2984 -146 3022 -118
rect 3050 -146 3088 -118
rect 3116 -146 3154 -118
rect 3182 -146 3220 -118
rect 3248 -146 3286 -118
rect 3314 -146 3352 -118
rect 3380 -146 3418 -118
rect 3446 -146 3484 -118
rect 3512 -146 3550 -118
rect 3578 -146 3616 -118
rect 3644 -146 3682 -118
rect 3710 -146 3748 -118
rect 3776 -146 3814 -118
rect 3842 -146 3880 -118
rect 3908 -146 3946 -118
rect 3974 -146 4012 -118
rect 4040 -146 4078 -118
rect 4106 -146 4144 -118
rect 4172 -146 4210 -118
rect 4238 -146 4276 -118
rect 4304 -146 4342 -118
rect 4370 -146 4408 -118
rect 4436 -146 4474 -118
rect 4502 -146 4540 -118
rect 4568 -146 4573 -118
rect -4573 -184 4573 -146
rect -4573 -212 -4568 -184
rect -4540 -212 -4502 -184
rect -4474 -212 -4436 -184
rect -4408 -212 -4370 -184
rect -4342 -212 -4304 -184
rect -4276 -212 -4238 -184
rect -4210 -212 -4172 -184
rect -4144 -212 -4106 -184
rect -4078 -212 -4040 -184
rect -4012 -212 -3974 -184
rect -3946 -212 -3908 -184
rect -3880 -212 -3842 -184
rect -3814 -212 -3776 -184
rect -3748 -212 -3710 -184
rect -3682 -212 -3644 -184
rect -3616 -212 -3578 -184
rect -3550 -212 -3512 -184
rect -3484 -212 -3446 -184
rect -3418 -212 -3380 -184
rect -3352 -212 -3314 -184
rect -3286 -212 -3248 -184
rect -3220 -212 -3182 -184
rect -3154 -212 -3116 -184
rect -3088 -212 -3050 -184
rect -3022 -212 -2984 -184
rect -2956 -212 -2918 -184
rect -2890 -212 -2852 -184
rect -2824 -212 -2786 -184
rect -2758 -212 -2720 -184
rect -2692 -212 -2654 -184
rect -2626 -212 -2588 -184
rect -2560 -212 -2522 -184
rect -2494 -212 -2456 -184
rect -2428 -212 -2390 -184
rect -2362 -212 -2324 -184
rect -2296 -212 -2258 -184
rect -2230 -212 -2192 -184
rect -2164 -212 -2126 -184
rect -2098 -212 -2060 -184
rect -2032 -212 -1994 -184
rect -1966 -212 -1928 -184
rect -1900 -212 -1862 -184
rect -1834 -212 -1796 -184
rect -1768 -212 -1730 -184
rect -1702 -212 -1664 -184
rect -1636 -212 -1598 -184
rect -1570 -212 -1532 -184
rect -1504 -212 -1466 -184
rect -1438 -212 -1400 -184
rect -1372 -212 -1334 -184
rect -1306 -212 -1268 -184
rect -1240 -212 -1202 -184
rect -1174 -212 -1136 -184
rect -1108 -212 -1070 -184
rect -1042 -212 -1004 -184
rect -976 -212 -938 -184
rect -910 -212 -872 -184
rect -844 -212 -806 -184
rect -778 -212 -740 -184
rect -712 -212 -674 -184
rect -646 -212 -608 -184
rect -580 -212 -542 -184
rect -514 -212 -476 -184
rect -448 -212 -410 -184
rect -382 -212 -344 -184
rect -316 -212 -278 -184
rect -250 -212 -212 -184
rect -184 -212 -146 -184
rect -118 -212 -80 -184
rect -52 -212 -14 -184
rect 14 -212 52 -184
rect 80 -212 118 -184
rect 146 -212 184 -184
rect 212 -212 250 -184
rect 278 -212 316 -184
rect 344 -212 382 -184
rect 410 -212 448 -184
rect 476 -212 514 -184
rect 542 -212 580 -184
rect 608 -212 646 -184
rect 674 -212 712 -184
rect 740 -212 778 -184
rect 806 -212 844 -184
rect 872 -212 910 -184
rect 938 -212 976 -184
rect 1004 -212 1042 -184
rect 1070 -212 1108 -184
rect 1136 -212 1174 -184
rect 1202 -212 1240 -184
rect 1268 -212 1306 -184
rect 1334 -212 1372 -184
rect 1400 -212 1438 -184
rect 1466 -212 1504 -184
rect 1532 -212 1570 -184
rect 1598 -212 1636 -184
rect 1664 -212 1702 -184
rect 1730 -212 1768 -184
rect 1796 -212 1834 -184
rect 1862 -212 1900 -184
rect 1928 -212 1966 -184
rect 1994 -212 2032 -184
rect 2060 -212 2098 -184
rect 2126 -212 2164 -184
rect 2192 -212 2230 -184
rect 2258 -212 2296 -184
rect 2324 -212 2362 -184
rect 2390 -212 2428 -184
rect 2456 -212 2494 -184
rect 2522 -212 2560 -184
rect 2588 -212 2626 -184
rect 2654 -212 2692 -184
rect 2720 -212 2758 -184
rect 2786 -212 2824 -184
rect 2852 -212 2890 -184
rect 2918 -212 2956 -184
rect 2984 -212 3022 -184
rect 3050 -212 3088 -184
rect 3116 -212 3154 -184
rect 3182 -212 3220 -184
rect 3248 -212 3286 -184
rect 3314 -212 3352 -184
rect 3380 -212 3418 -184
rect 3446 -212 3484 -184
rect 3512 -212 3550 -184
rect 3578 -212 3616 -184
rect 3644 -212 3682 -184
rect 3710 -212 3748 -184
rect 3776 -212 3814 -184
rect 3842 -212 3880 -184
rect 3908 -212 3946 -184
rect 3974 -212 4012 -184
rect 4040 -212 4078 -184
rect 4106 -212 4144 -184
rect 4172 -212 4210 -184
rect 4238 -212 4276 -184
rect 4304 -212 4342 -184
rect 4370 -212 4408 -184
rect 4436 -212 4474 -184
rect 4502 -212 4540 -184
rect 4568 -212 4573 -184
rect -4573 -250 4573 -212
rect -4573 -278 -4568 -250
rect -4540 -278 -4502 -250
rect -4474 -278 -4436 -250
rect -4408 -278 -4370 -250
rect -4342 -278 -4304 -250
rect -4276 -278 -4238 -250
rect -4210 -278 -4172 -250
rect -4144 -278 -4106 -250
rect -4078 -278 -4040 -250
rect -4012 -278 -3974 -250
rect -3946 -278 -3908 -250
rect -3880 -278 -3842 -250
rect -3814 -278 -3776 -250
rect -3748 -278 -3710 -250
rect -3682 -278 -3644 -250
rect -3616 -278 -3578 -250
rect -3550 -278 -3512 -250
rect -3484 -278 -3446 -250
rect -3418 -278 -3380 -250
rect -3352 -278 -3314 -250
rect -3286 -278 -3248 -250
rect -3220 -278 -3182 -250
rect -3154 -278 -3116 -250
rect -3088 -278 -3050 -250
rect -3022 -278 -2984 -250
rect -2956 -278 -2918 -250
rect -2890 -278 -2852 -250
rect -2824 -278 -2786 -250
rect -2758 -278 -2720 -250
rect -2692 -278 -2654 -250
rect -2626 -278 -2588 -250
rect -2560 -278 -2522 -250
rect -2494 -278 -2456 -250
rect -2428 -278 -2390 -250
rect -2362 -278 -2324 -250
rect -2296 -278 -2258 -250
rect -2230 -278 -2192 -250
rect -2164 -278 -2126 -250
rect -2098 -278 -2060 -250
rect -2032 -278 -1994 -250
rect -1966 -278 -1928 -250
rect -1900 -278 -1862 -250
rect -1834 -278 -1796 -250
rect -1768 -278 -1730 -250
rect -1702 -278 -1664 -250
rect -1636 -278 -1598 -250
rect -1570 -278 -1532 -250
rect -1504 -278 -1466 -250
rect -1438 -278 -1400 -250
rect -1372 -278 -1334 -250
rect -1306 -278 -1268 -250
rect -1240 -278 -1202 -250
rect -1174 -278 -1136 -250
rect -1108 -278 -1070 -250
rect -1042 -278 -1004 -250
rect -976 -278 -938 -250
rect -910 -278 -872 -250
rect -844 -278 -806 -250
rect -778 -278 -740 -250
rect -712 -278 -674 -250
rect -646 -278 -608 -250
rect -580 -278 -542 -250
rect -514 -278 -476 -250
rect -448 -278 -410 -250
rect -382 -278 -344 -250
rect -316 -278 -278 -250
rect -250 -278 -212 -250
rect -184 -278 -146 -250
rect -118 -278 -80 -250
rect -52 -278 -14 -250
rect 14 -278 52 -250
rect 80 -278 118 -250
rect 146 -278 184 -250
rect 212 -278 250 -250
rect 278 -278 316 -250
rect 344 -278 382 -250
rect 410 -278 448 -250
rect 476 -278 514 -250
rect 542 -278 580 -250
rect 608 -278 646 -250
rect 674 -278 712 -250
rect 740 -278 778 -250
rect 806 -278 844 -250
rect 872 -278 910 -250
rect 938 -278 976 -250
rect 1004 -278 1042 -250
rect 1070 -278 1108 -250
rect 1136 -278 1174 -250
rect 1202 -278 1240 -250
rect 1268 -278 1306 -250
rect 1334 -278 1372 -250
rect 1400 -278 1438 -250
rect 1466 -278 1504 -250
rect 1532 -278 1570 -250
rect 1598 -278 1636 -250
rect 1664 -278 1702 -250
rect 1730 -278 1768 -250
rect 1796 -278 1834 -250
rect 1862 -278 1900 -250
rect 1928 -278 1966 -250
rect 1994 -278 2032 -250
rect 2060 -278 2098 -250
rect 2126 -278 2164 -250
rect 2192 -278 2230 -250
rect 2258 -278 2296 -250
rect 2324 -278 2362 -250
rect 2390 -278 2428 -250
rect 2456 -278 2494 -250
rect 2522 -278 2560 -250
rect 2588 -278 2626 -250
rect 2654 -278 2692 -250
rect 2720 -278 2758 -250
rect 2786 -278 2824 -250
rect 2852 -278 2890 -250
rect 2918 -278 2956 -250
rect 2984 -278 3022 -250
rect 3050 -278 3088 -250
rect 3116 -278 3154 -250
rect 3182 -278 3220 -250
rect 3248 -278 3286 -250
rect 3314 -278 3352 -250
rect 3380 -278 3418 -250
rect 3446 -278 3484 -250
rect 3512 -278 3550 -250
rect 3578 -278 3616 -250
rect 3644 -278 3682 -250
rect 3710 -278 3748 -250
rect 3776 -278 3814 -250
rect 3842 -278 3880 -250
rect 3908 -278 3946 -250
rect 3974 -278 4012 -250
rect 4040 -278 4078 -250
rect 4106 -278 4144 -250
rect 4172 -278 4210 -250
rect 4238 -278 4276 -250
rect 4304 -278 4342 -250
rect 4370 -278 4408 -250
rect 4436 -278 4474 -250
rect 4502 -278 4540 -250
rect 4568 -278 4573 -250
rect -4573 -316 4573 -278
rect -4573 -344 -4568 -316
rect -4540 -344 -4502 -316
rect -4474 -344 -4436 -316
rect -4408 -344 -4370 -316
rect -4342 -344 -4304 -316
rect -4276 -344 -4238 -316
rect -4210 -344 -4172 -316
rect -4144 -344 -4106 -316
rect -4078 -344 -4040 -316
rect -4012 -344 -3974 -316
rect -3946 -344 -3908 -316
rect -3880 -344 -3842 -316
rect -3814 -344 -3776 -316
rect -3748 -344 -3710 -316
rect -3682 -344 -3644 -316
rect -3616 -344 -3578 -316
rect -3550 -344 -3512 -316
rect -3484 -344 -3446 -316
rect -3418 -344 -3380 -316
rect -3352 -344 -3314 -316
rect -3286 -344 -3248 -316
rect -3220 -344 -3182 -316
rect -3154 -344 -3116 -316
rect -3088 -344 -3050 -316
rect -3022 -344 -2984 -316
rect -2956 -344 -2918 -316
rect -2890 -344 -2852 -316
rect -2824 -344 -2786 -316
rect -2758 -344 -2720 -316
rect -2692 -344 -2654 -316
rect -2626 -344 -2588 -316
rect -2560 -344 -2522 -316
rect -2494 -344 -2456 -316
rect -2428 -344 -2390 -316
rect -2362 -344 -2324 -316
rect -2296 -344 -2258 -316
rect -2230 -344 -2192 -316
rect -2164 -344 -2126 -316
rect -2098 -344 -2060 -316
rect -2032 -344 -1994 -316
rect -1966 -344 -1928 -316
rect -1900 -344 -1862 -316
rect -1834 -344 -1796 -316
rect -1768 -344 -1730 -316
rect -1702 -344 -1664 -316
rect -1636 -344 -1598 -316
rect -1570 -344 -1532 -316
rect -1504 -344 -1466 -316
rect -1438 -344 -1400 -316
rect -1372 -344 -1334 -316
rect -1306 -344 -1268 -316
rect -1240 -344 -1202 -316
rect -1174 -344 -1136 -316
rect -1108 -344 -1070 -316
rect -1042 -344 -1004 -316
rect -976 -344 -938 -316
rect -910 -344 -872 -316
rect -844 -344 -806 -316
rect -778 -344 -740 -316
rect -712 -344 -674 -316
rect -646 -344 -608 -316
rect -580 -344 -542 -316
rect -514 -344 -476 -316
rect -448 -344 -410 -316
rect -382 -344 -344 -316
rect -316 -344 -278 -316
rect -250 -344 -212 -316
rect -184 -344 -146 -316
rect -118 -344 -80 -316
rect -52 -344 -14 -316
rect 14 -344 52 -316
rect 80 -344 118 -316
rect 146 -344 184 -316
rect 212 -344 250 -316
rect 278 -344 316 -316
rect 344 -344 382 -316
rect 410 -344 448 -316
rect 476 -344 514 -316
rect 542 -344 580 -316
rect 608 -344 646 -316
rect 674 -344 712 -316
rect 740 -344 778 -316
rect 806 -344 844 -316
rect 872 -344 910 -316
rect 938 -344 976 -316
rect 1004 -344 1042 -316
rect 1070 -344 1108 -316
rect 1136 -344 1174 -316
rect 1202 -344 1240 -316
rect 1268 -344 1306 -316
rect 1334 -344 1372 -316
rect 1400 -344 1438 -316
rect 1466 -344 1504 -316
rect 1532 -344 1570 -316
rect 1598 -344 1636 -316
rect 1664 -344 1702 -316
rect 1730 -344 1768 -316
rect 1796 -344 1834 -316
rect 1862 -344 1900 -316
rect 1928 -344 1966 -316
rect 1994 -344 2032 -316
rect 2060 -344 2098 -316
rect 2126 -344 2164 -316
rect 2192 -344 2230 -316
rect 2258 -344 2296 -316
rect 2324 -344 2362 -316
rect 2390 -344 2428 -316
rect 2456 -344 2494 -316
rect 2522 -344 2560 -316
rect 2588 -344 2626 -316
rect 2654 -344 2692 -316
rect 2720 -344 2758 -316
rect 2786 -344 2824 -316
rect 2852 -344 2890 -316
rect 2918 -344 2956 -316
rect 2984 -344 3022 -316
rect 3050 -344 3088 -316
rect 3116 -344 3154 -316
rect 3182 -344 3220 -316
rect 3248 -344 3286 -316
rect 3314 -344 3352 -316
rect 3380 -344 3418 -316
rect 3446 -344 3484 -316
rect 3512 -344 3550 -316
rect 3578 -344 3616 -316
rect 3644 -344 3682 -316
rect 3710 -344 3748 -316
rect 3776 -344 3814 -316
rect 3842 -344 3880 -316
rect 3908 -344 3946 -316
rect 3974 -344 4012 -316
rect 4040 -344 4078 -316
rect 4106 -344 4144 -316
rect 4172 -344 4210 -316
rect 4238 -344 4276 -316
rect 4304 -344 4342 -316
rect 4370 -344 4408 -316
rect 4436 -344 4474 -316
rect 4502 -344 4540 -316
rect 4568 -344 4573 -316
rect -4573 -382 4573 -344
rect -4573 -410 -4568 -382
rect -4540 -410 -4502 -382
rect -4474 -410 -4436 -382
rect -4408 -410 -4370 -382
rect -4342 -410 -4304 -382
rect -4276 -410 -4238 -382
rect -4210 -410 -4172 -382
rect -4144 -410 -4106 -382
rect -4078 -410 -4040 -382
rect -4012 -410 -3974 -382
rect -3946 -410 -3908 -382
rect -3880 -410 -3842 -382
rect -3814 -410 -3776 -382
rect -3748 -410 -3710 -382
rect -3682 -410 -3644 -382
rect -3616 -410 -3578 -382
rect -3550 -410 -3512 -382
rect -3484 -410 -3446 -382
rect -3418 -410 -3380 -382
rect -3352 -410 -3314 -382
rect -3286 -410 -3248 -382
rect -3220 -410 -3182 -382
rect -3154 -410 -3116 -382
rect -3088 -410 -3050 -382
rect -3022 -410 -2984 -382
rect -2956 -410 -2918 -382
rect -2890 -410 -2852 -382
rect -2824 -410 -2786 -382
rect -2758 -410 -2720 -382
rect -2692 -410 -2654 -382
rect -2626 -410 -2588 -382
rect -2560 -410 -2522 -382
rect -2494 -410 -2456 -382
rect -2428 -410 -2390 -382
rect -2362 -410 -2324 -382
rect -2296 -410 -2258 -382
rect -2230 -410 -2192 -382
rect -2164 -410 -2126 -382
rect -2098 -410 -2060 -382
rect -2032 -410 -1994 -382
rect -1966 -410 -1928 -382
rect -1900 -410 -1862 -382
rect -1834 -410 -1796 -382
rect -1768 -410 -1730 -382
rect -1702 -410 -1664 -382
rect -1636 -410 -1598 -382
rect -1570 -410 -1532 -382
rect -1504 -410 -1466 -382
rect -1438 -410 -1400 -382
rect -1372 -410 -1334 -382
rect -1306 -410 -1268 -382
rect -1240 -410 -1202 -382
rect -1174 -410 -1136 -382
rect -1108 -410 -1070 -382
rect -1042 -410 -1004 -382
rect -976 -410 -938 -382
rect -910 -410 -872 -382
rect -844 -410 -806 -382
rect -778 -410 -740 -382
rect -712 -410 -674 -382
rect -646 -410 -608 -382
rect -580 -410 -542 -382
rect -514 -410 -476 -382
rect -448 -410 -410 -382
rect -382 -410 -344 -382
rect -316 -410 -278 -382
rect -250 -410 -212 -382
rect -184 -410 -146 -382
rect -118 -410 -80 -382
rect -52 -410 -14 -382
rect 14 -410 52 -382
rect 80 -410 118 -382
rect 146 -410 184 -382
rect 212 -410 250 -382
rect 278 -410 316 -382
rect 344 -410 382 -382
rect 410 -410 448 -382
rect 476 -410 514 -382
rect 542 -410 580 -382
rect 608 -410 646 -382
rect 674 -410 712 -382
rect 740 -410 778 -382
rect 806 -410 844 -382
rect 872 -410 910 -382
rect 938 -410 976 -382
rect 1004 -410 1042 -382
rect 1070 -410 1108 -382
rect 1136 -410 1174 -382
rect 1202 -410 1240 -382
rect 1268 -410 1306 -382
rect 1334 -410 1372 -382
rect 1400 -410 1438 -382
rect 1466 -410 1504 -382
rect 1532 -410 1570 -382
rect 1598 -410 1636 -382
rect 1664 -410 1702 -382
rect 1730 -410 1768 -382
rect 1796 -410 1834 -382
rect 1862 -410 1900 -382
rect 1928 -410 1966 -382
rect 1994 -410 2032 -382
rect 2060 -410 2098 -382
rect 2126 -410 2164 -382
rect 2192 -410 2230 -382
rect 2258 -410 2296 -382
rect 2324 -410 2362 -382
rect 2390 -410 2428 -382
rect 2456 -410 2494 -382
rect 2522 -410 2560 -382
rect 2588 -410 2626 -382
rect 2654 -410 2692 -382
rect 2720 -410 2758 -382
rect 2786 -410 2824 -382
rect 2852 -410 2890 -382
rect 2918 -410 2956 -382
rect 2984 -410 3022 -382
rect 3050 -410 3088 -382
rect 3116 -410 3154 -382
rect 3182 -410 3220 -382
rect 3248 -410 3286 -382
rect 3314 -410 3352 -382
rect 3380 -410 3418 -382
rect 3446 -410 3484 -382
rect 3512 -410 3550 -382
rect 3578 -410 3616 -382
rect 3644 -410 3682 -382
rect 3710 -410 3748 -382
rect 3776 -410 3814 -382
rect 3842 -410 3880 -382
rect 3908 -410 3946 -382
rect 3974 -410 4012 -382
rect 4040 -410 4078 -382
rect 4106 -410 4144 -382
rect 4172 -410 4210 -382
rect 4238 -410 4276 -382
rect 4304 -410 4342 -382
rect 4370 -410 4408 -382
rect 4436 -410 4474 -382
rect 4502 -410 4540 -382
rect 4568 -410 4573 -382
rect -4573 -448 4573 -410
rect -4573 -476 -4568 -448
rect -4540 -476 -4502 -448
rect -4474 -476 -4436 -448
rect -4408 -476 -4370 -448
rect -4342 -476 -4304 -448
rect -4276 -476 -4238 -448
rect -4210 -476 -4172 -448
rect -4144 -476 -4106 -448
rect -4078 -476 -4040 -448
rect -4012 -476 -3974 -448
rect -3946 -476 -3908 -448
rect -3880 -476 -3842 -448
rect -3814 -476 -3776 -448
rect -3748 -476 -3710 -448
rect -3682 -476 -3644 -448
rect -3616 -476 -3578 -448
rect -3550 -476 -3512 -448
rect -3484 -476 -3446 -448
rect -3418 -476 -3380 -448
rect -3352 -476 -3314 -448
rect -3286 -476 -3248 -448
rect -3220 -476 -3182 -448
rect -3154 -476 -3116 -448
rect -3088 -476 -3050 -448
rect -3022 -476 -2984 -448
rect -2956 -476 -2918 -448
rect -2890 -476 -2852 -448
rect -2824 -476 -2786 -448
rect -2758 -476 -2720 -448
rect -2692 -476 -2654 -448
rect -2626 -476 -2588 -448
rect -2560 -476 -2522 -448
rect -2494 -476 -2456 -448
rect -2428 -476 -2390 -448
rect -2362 -476 -2324 -448
rect -2296 -476 -2258 -448
rect -2230 -476 -2192 -448
rect -2164 -476 -2126 -448
rect -2098 -476 -2060 -448
rect -2032 -476 -1994 -448
rect -1966 -476 -1928 -448
rect -1900 -476 -1862 -448
rect -1834 -476 -1796 -448
rect -1768 -476 -1730 -448
rect -1702 -476 -1664 -448
rect -1636 -476 -1598 -448
rect -1570 -476 -1532 -448
rect -1504 -476 -1466 -448
rect -1438 -476 -1400 -448
rect -1372 -476 -1334 -448
rect -1306 -476 -1268 -448
rect -1240 -476 -1202 -448
rect -1174 -476 -1136 -448
rect -1108 -476 -1070 -448
rect -1042 -476 -1004 -448
rect -976 -476 -938 -448
rect -910 -476 -872 -448
rect -844 -476 -806 -448
rect -778 -476 -740 -448
rect -712 -476 -674 -448
rect -646 -476 -608 -448
rect -580 -476 -542 -448
rect -514 -476 -476 -448
rect -448 -476 -410 -448
rect -382 -476 -344 -448
rect -316 -476 -278 -448
rect -250 -476 -212 -448
rect -184 -476 -146 -448
rect -118 -476 -80 -448
rect -52 -476 -14 -448
rect 14 -476 52 -448
rect 80 -476 118 -448
rect 146 -476 184 -448
rect 212 -476 250 -448
rect 278 -476 316 -448
rect 344 -476 382 -448
rect 410 -476 448 -448
rect 476 -476 514 -448
rect 542 -476 580 -448
rect 608 -476 646 -448
rect 674 -476 712 -448
rect 740 -476 778 -448
rect 806 -476 844 -448
rect 872 -476 910 -448
rect 938 -476 976 -448
rect 1004 -476 1042 -448
rect 1070 -476 1108 -448
rect 1136 -476 1174 -448
rect 1202 -476 1240 -448
rect 1268 -476 1306 -448
rect 1334 -476 1372 -448
rect 1400 -476 1438 -448
rect 1466 -476 1504 -448
rect 1532 -476 1570 -448
rect 1598 -476 1636 -448
rect 1664 -476 1702 -448
rect 1730 -476 1768 -448
rect 1796 -476 1834 -448
rect 1862 -476 1900 -448
rect 1928 -476 1966 -448
rect 1994 -476 2032 -448
rect 2060 -476 2098 -448
rect 2126 -476 2164 -448
rect 2192 -476 2230 -448
rect 2258 -476 2296 -448
rect 2324 -476 2362 -448
rect 2390 -476 2428 -448
rect 2456 -476 2494 -448
rect 2522 -476 2560 -448
rect 2588 -476 2626 -448
rect 2654 -476 2692 -448
rect 2720 -476 2758 -448
rect 2786 -476 2824 -448
rect 2852 -476 2890 -448
rect 2918 -476 2956 -448
rect 2984 -476 3022 -448
rect 3050 -476 3088 -448
rect 3116 -476 3154 -448
rect 3182 -476 3220 -448
rect 3248 -476 3286 -448
rect 3314 -476 3352 -448
rect 3380 -476 3418 -448
rect 3446 -476 3484 -448
rect 3512 -476 3550 -448
rect 3578 -476 3616 -448
rect 3644 -476 3682 -448
rect 3710 -476 3748 -448
rect 3776 -476 3814 -448
rect 3842 -476 3880 -448
rect 3908 -476 3946 -448
rect 3974 -476 4012 -448
rect 4040 -476 4078 -448
rect 4106 -476 4144 -448
rect 4172 -476 4210 -448
rect 4238 -476 4276 -448
rect 4304 -476 4342 -448
rect 4370 -476 4408 -448
rect 4436 -476 4474 -448
rect 4502 -476 4540 -448
rect 4568 -476 4573 -448
rect -4573 -514 4573 -476
rect -4573 -542 -4568 -514
rect -4540 -542 -4502 -514
rect -4474 -542 -4436 -514
rect -4408 -542 -4370 -514
rect -4342 -542 -4304 -514
rect -4276 -542 -4238 -514
rect -4210 -542 -4172 -514
rect -4144 -542 -4106 -514
rect -4078 -542 -4040 -514
rect -4012 -542 -3974 -514
rect -3946 -542 -3908 -514
rect -3880 -542 -3842 -514
rect -3814 -542 -3776 -514
rect -3748 -542 -3710 -514
rect -3682 -542 -3644 -514
rect -3616 -542 -3578 -514
rect -3550 -542 -3512 -514
rect -3484 -542 -3446 -514
rect -3418 -542 -3380 -514
rect -3352 -542 -3314 -514
rect -3286 -542 -3248 -514
rect -3220 -542 -3182 -514
rect -3154 -542 -3116 -514
rect -3088 -542 -3050 -514
rect -3022 -542 -2984 -514
rect -2956 -542 -2918 -514
rect -2890 -542 -2852 -514
rect -2824 -542 -2786 -514
rect -2758 -542 -2720 -514
rect -2692 -542 -2654 -514
rect -2626 -542 -2588 -514
rect -2560 -542 -2522 -514
rect -2494 -542 -2456 -514
rect -2428 -542 -2390 -514
rect -2362 -542 -2324 -514
rect -2296 -542 -2258 -514
rect -2230 -542 -2192 -514
rect -2164 -542 -2126 -514
rect -2098 -542 -2060 -514
rect -2032 -542 -1994 -514
rect -1966 -542 -1928 -514
rect -1900 -542 -1862 -514
rect -1834 -542 -1796 -514
rect -1768 -542 -1730 -514
rect -1702 -542 -1664 -514
rect -1636 -542 -1598 -514
rect -1570 -542 -1532 -514
rect -1504 -542 -1466 -514
rect -1438 -542 -1400 -514
rect -1372 -542 -1334 -514
rect -1306 -542 -1268 -514
rect -1240 -542 -1202 -514
rect -1174 -542 -1136 -514
rect -1108 -542 -1070 -514
rect -1042 -542 -1004 -514
rect -976 -542 -938 -514
rect -910 -542 -872 -514
rect -844 -542 -806 -514
rect -778 -542 -740 -514
rect -712 -542 -674 -514
rect -646 -542 -608 -514
rect -580 -542 -542 -514
rect -514 -542 -476 -514
rect -448 -542 -410 -514
rect -382 -542 -344 -514
rect -316 -542 -278 -514
rect -250 -542 -212 -514
rect -184 -542 -146 -514
rect -118 -542 -80 -514
rect -52 -542 -14 -514
rect 14 -542 52 -514
rect 80 -542 118 -514
rect 146 -542 184 -514
rect 212 -542 250 -514
rect 278 -542 316 -514
rect 344 -542 382 -514
rect 410 -542 448 -514
rect 476 -542 514 -514
rect 542 -542 580 -514
rect 608 -542 646 -514
rect 674 -542 712 -514
rect 740 -542 778 -514
rect 806 -542 844 -514
rect 872 -542 910 -514
rect 938 -542 976 -514
rect 1004 -542 1042 -514
rect 1070 -542 1108 -514
rect 1136 -542 1174 -514
rect 1202 -542 1240 -514
rect 1268 -542 1306 -514
rect 1334 -542 1372 -514
rect 1400 -542 1438 -514
rect 1466 -542 1504 -514
rect 1532 -542 1570 -514
rect 1598 -542 1636 -514
rect 1664 -542 1702 -514
rect 1730 -542 1768 -514
rect 1796 -542 1834 -514
rect 1862 -542 1900 -514
rect 1928 -542 1966 -514
rect 1994 -542 2032 -514
rect 2060 -542 2098 -514
rect 2126 -542 2164 -514
rect 2192 -542 2230 -514
rect 2258 -542 2296 -514
rect 2324 -542 2362 -514
rect 2390 -542 2428 -514
rect 2456 -542 2494 -514
rect 2522 -542 2560 -514
rect 2588 -542 2626 -514
rect 2654 -542 2692 -514
rect 2720 -542 2758 -514
rect 2786 -542 2824 -514
rect 2852 -542 2890 -514
rect 2918 -542 2956 -514
rect 2984 -542 3022 -514
rect 3050 -542 3088 -514
rect 3116 -542 3154 -514
rect 3182 -542 3220 -514
rect 3248 -542 3286 -514
rect 3314 -542 3352 -514
rect 3380 -542 3418 -514
rect 3446 -542 3484 -514
rect 3512 -542 3550 -514
rect 3578 -542 3616 -514
rect 3644 -542 3682 -514
rect 3710 -542 3748 -514
rect 3776 -542 3814 -514
rect 3842 -542 3880 -514
rect 3908 -542 3946 -514
rect 3974 -542 4012 -514
rect 4040 -542 4078 -514
rect 4106 -542 4144 -514
rect 4172 -542 4210 -514
rect 4238 -542 4276 -514
rect 4304 -542 4342 -514
rect 4370 -542 4408 -514
rect 4436 -542 4474 -514
rect 4502 -542 4540 -514
rect 4568 -542 4573 -514
rect -4573 -580 4573 -542
rect -4573 -608 -4568 -580
rect -4540 -608 -4502 -580
rect -4474 -608 -4436 -580
rect -4408 -608 -4370 -580
rect -4342 -608 -4304 -580
rect -4276 -608 -4238 -580
rect -4210 -608 -4172 -580
rect -4144 -608 -4106 -580
rect -4078 -608 -4040 -580
rect -4012 -608 -3974 -580
rect -3946 -608 -3908 -580
rect -3880 -608 -3842 -580
rect -3814 -608 -3776 -580
rect -3748 -608 -3710 -580
rect -3682 -608 -3644 -580
rect -3616 -608 -3578 -580
rect -3550 -608 -3512 -580
rect -3484 -608 -3446 -580
rect -3418 -608 -3380 -580
rect -3352 -608 -3314 -580
rect -3286 -608 -3248 -580
rect -3220 -608 -3182 -580
rect -3154 -608 -3116 -580
rect -3088 -608 -3050 -580
rect -3022 -608 -2984 -580
rect -2956 -608 -2918 -580
rect -2890 -608 -2852 -580
rect -2824 -608 -2786 -580
rect -2758 -608 -2720 -580
rect -2692 -608 -2654 -580
rect -2626 -608 -2588 -580
rect -2560 -608 -2522 -580
rect -2494 -608 -2456 -580
rect -2428 -608 -2390 -580
rect -2362 -608 -2324 -580
rect -2296 -608 -2258 -580
rect -2230 -608 -2192 -580
rect -2164 -608 -2126 -580
rect -2098 -608 -2060 -580
rect -2032 -608 -1994 -580
rect -1966 -608 -1928 -580
rect -1900 -608 -1862 -580
rect -1834 -608 -1796 -580
rect -1768 -608 -1730 -580
rect -1702 -608 -1664 -580
rect -1636 -608 -1598 -580
rect -1570 -608 -1532 -580
rect -1504 -608 -1466 -580
rect -1438 -608 -1400 -580
rect -1372 -608 -1334 -580
rect -1306 -608 -1268 -580
rect -1240 -608 -1202 -580
rect -1174 -608 -1136 -580
rect -1108 -608 -1070 -580
rect -1042 -608 -1004 -580
rect -976 -608 -938 -580
rect -910 -608 -872 -580
rect -844 -608 -806 -580
rect -778 -608 -740 -580
rect -712 -608 -674 -580
rect -646 -608 -608 -580
rect -580 -608 -542 -580
rect -514 -608 -476 -580
rect -448 -608 -410 -580
rect -382 -608 -344 -580
rect -316 -608 -278 -580
rect -250 -608 -212 -580
rect -184 -608 -146 -580
rect -118 -608 -80 -580
rect -52 -608 -14 -580
rect 14 -608 52 -580
rect 80 -608 118 -580
rect 146 -608 184 -580
rect 212 -608 250 -580
rect 278 -608 316 -580
rect 344 -608 382 -580
rect 410 -608 448 -580
rect 476 -608 514 -580
rect 542 -608 580 -580
rect 608 -608 646 -580
rect 674 -608 712 -580
rect 740 -608 778 -580
rect 806 -608 844 -580
rect 872 -608 910 -580
rect 938 -608 976 -580
rect 1004 -608 1042 -580
rect 1070 -608 1108 -580
rect 1136 -608 1174 -580
rect 1202 -608 1240 -580
rect 1268 -608 1306 -580
rect 1334 -608 1372 -580
rect 1400 -608 1438 -580
rect 1466 -608 1504 -580
rect 1532 -608 1570 -580
rect 1598 -608 1636 -580
rect 1664 -608 1702 -580
rect 1730 -608 1768 -580
rect 1796 -608 1834 -580
rect 1862 -608 1900 -580
rect 1928 -608 1966 -580
rect 1994 -608 2032 -580
rect 2060 -608 2098 -580
rect 2126 -608 2164 -580
rect 2192 -608 2230 -580
rect 2258 -608 2296 -580
rect 2324 -608 2362 -580
rect 2390 -608 2428 -580
rect 2456 -608 2494 -580
rect 2522 -608 2560 -580
rect 2588 -608 2626 -580
rect 2654 -608 2692 -580
rect 2720 -608 2758 -580
rect 2786 -608 2824 -580
rect 2852 -608 2890 -580
rect 2918 -608 2956 -580
rect 2984 -608 3022 -580
rect 3050 -608 3088 -580
rect 3116 -608 3154 -580
rect 3182 -608 3220 -580
rect 3248 -608 3286 -580
rect 3314 -608 3352 -580
rect 3380 -608 3418 -580
rect 3446 -608 3484 -580
rect 3512 -608 3550 -580
rect 3578 -608 3616 -580
rect 3644 -608 3682 -580
rect 3710 -608 3748 -580
rect 3776 -608 3814 -580
rect 3842 -608 3880 -580
rect 3908 -608 3946 -580
rect 3974 -608 4012 -580
rect 4040 -608 4078 -580
rect 4106 -608 4144 -580
rect 4172 -608 4210 -580
rect 4238 -608 4276 -580
rect 4304 -608 4342 -580
rect 4370 -608 4408 -580
rect 4436 -608 4474 -580
rect 4502 -608 4540 -580
rect 4568 -608 4573 -580
rect -4573 -646 4573 -608
rect -4573 -674 -4568 -646
rect -4540 -674 -4502 -646
rect -4474 -674 -4436 -646
rect -4408 -674 -4370 -646
rect -4342 -674 -4304 -646
rect -4276 -674 -4238 -646
rect -4210 -674 -4172 -646
rect -4144 -674 -4106 -646
rect -4078 -674 -4040 -646
rect -4012 -674 -3974 -646
rect -3946 -674 -3908 -646
rect -3880 -674 -3842 -646
rect -3814 -674 -3776 -646
rect -3748 -674 -3710 -646
rect -3682 -674 -3644 -646
rect -3616 -674 -3578 -646
rect -3550 -674 -3512 -646
rect -3484 -674 -3446 -646
rect -3418 -674 -3380 -646
rect -3352 -674 -3314 -646
rect -3286 -674 -3248 -646
rect -3220 -674 -3182 -646
rect -3154 -674 -3116 -646
rect -3088 -674 -3050 -646
rect -3022 -674 -2984 -646
rect -2956 -674 -2918 -646
rect -2890 -674 -2852 -646
rect -2824 -674 -2786 -646
rect -2758 -674 -2720 -646
rect -2692 -674 -2654 -646
rect -2626 -674 -2588 -646
rect -2560 -674 -2522 -646
rect -2494 -674 -2456 -646
rect -2428 -674 -2390 -646
rect -2362 -674 -2324 -646
rect -2296 -674 -2258 -646
rect -2230 -674 -2192 -646
rect -2164 -674 -2126 -646
rect -2098 -674 -2060 -646
rect -2032 -674 -1994 -646
rect -1966 -674 -1928 -646
rect -1900 -674 -1862 -646
rect -1834 -674 -1796 -646
rect -1768 -674 -1730 -646
rect -1702 -674 -1664 -646
rect -1636 -674 -1598 -646
rect -1570 -674 -1532 -646
rect -1504 -674 -1466 -646
rect -1438 -674 -1400 -646
rect -1372 -674 -1334 -646
rect -1306 -674 -1268 -646
rect -1240 -674 -1202 -646
rect -1174 -674 -1136 -646
rect -1108 -674 -1070 -646
rect -1042 -674 -1004 -646
rect -976 -674 -938 -646
rect -910 -674 -872 -646
rect -844 -674 -806 -646
rect -778 -674 -740 -646
rect -712 -674 -674 -646
rect -646 -674 -608 -646
rect -580 -674 -542 -646
rect -514 -674 -476 -646
rect -448 -674 -410 -646
rect -382 -674 -344 -646
rect -316 -674 -278 -646
rect -250 -674 -212 -646
rect -184 -674 -146 -646
rect -118 -674 -80 -646
rect -52 -674 -14 -646
rect 14 -674 52 -646
rect 80 -674 118 -646
rect 146 -674 184 -646
rect 212 -674 250 -646
rect 278 -674 316 -646
rect 344 -674 382 -646
rect 410 -674 448 -646
rect 476 -674 514 -646
rect 542 -674 580 -646
rect 608 -674 646 -646
rect 674 -674 712 -646
rect 740 -674 778 -646
rect 806 -674 844 -646
rect 872 -674 910 -646
rect 938 -674 976 -646
rect 1004 -674 1042 -646
rect 1070 -674 1108 -646
rect 1136 -674 1174 -646
rect 1202 -674 1240 -646
rect 1268 -674 1306 -646
rect 1334 -674 1372 -646
rect 1400 -674 1438 -646
rect 1466 -674 1504 -646
rect 1532 -674 1570 -646
rect 1598 -674 1636 -646
rect 1664 -674 1702 -646
rect 1730 -674 1768 -646
rect 1796 -674 1834 -646
rect 1862 -674 1900 -646
rect 1928 -674 1966 -646
rect 1994 -674 2032 -646
rect 2060 -674 2098 -646
rect 2126 -674 2164 -646
rect 2192 -674 2230 -646
rect 2258 -674 2296 -646
rect 2324 -674 2362 -646
rect 2390 -674 2428 -646
rect 2456 -674 2494 -646
rect 2522 -674 2560 -646
rect 2588 -674 2626 -646
rect 2654 -674 2692 -646
rect 2720 -674 2758 -646
rect 2786 -674 2824 -646
rect 2852 -674 2890 -646
rect 2918 -674 2956 -646
rect 2984 -674 3022 -646
rect 3050 -674 3088 -646
rect 3116 -674 3154 -646
rect 3182 -674 3220 -646
rect 3248 -674 3286 -646
rect 3314 -674 3352 -646
rect 3380 -674 3418 -646
rect 3446 -674 3484 -646
rect 3512 -674 3550 -646
rect 3578 -674 3616 -646
rect 3644 -674 3682 -646
rect 3710 -674 3748 -646
rect 3776 -674 3814 -646
rect 3842 -674 3880 -646
rect 3908 -674 3946 -646
rect 3974 -674 4012 -646
rect 4040 -674 4078 -646
rect 4106 -674 4144 -646
rect 4172 -674 4210 -646
rect 4238 -674 4276 -646
rect 4304 -674 4342 -646
rect 4370 -674 4408 -646
rect 4436 -674 4474 -646
rect 4502 -674 4540 -646
rect 4568 -674 4573 -646
rect -4573 -712 4573 -674
rect -4573 -740 -4568 -712
rect -4540 -740 -4502 -712
rect -4474 -740 -4436 -712
rect -4408 -740 -4370 -712
rect -4342 -740 -4304 -712
rect -4276 -740 -4238 -712
rect -4210 -740 -4172 -712
rect -4144 -740 -4106 -712
rect -4078 -740 -4040 -712
rect -4012 -740 -3974 -712
rect -3946 -740 -3908 -712
rect -3880 -740 -3842 -712
rect -3814 -740 -3776 -712
rect -3748 -740 -3710 -712
rect -3682 -740 -3644 -712
rect -3616 -740 -3578 -712
rect -3550 -740 -3512 -712
rect -3484 -740 -3446 -712
rect -3418 -740 -3380 -712
rect -3352 -740 -3314 -712
rect -3286 -740 -3248 -712
rect -3220 -740 -3182 -712
rect -3154 -740 -3116 -712
rect -3088 -740 -3050 -712
rect -3022 -740 -2984 -712
rect -2956 -740 -2918 -712
rect -2890 -740 -2852 -712
rect -2824 -740 -2786 -712
rect -2758 -740 -2720 -712
rect -2692 -740 -2654 -712
rect -2626 -740 -2588 -712
rect -2560 -740 -2522 -712
rect -2494 -740 -2456 -712
rect -2428 -740 -2390 -712
rect -2362 -740 -2324 -712
rect -2296 -740 -2258 -712
rect -2230 -740 -2192 -712
rect -2164 -740 -2126 -712
rect -2098 -740 -2060 -712
rect -2032 -740 -1994 -712
rect -1966 -740 -1928 -712
rect -1900 -740 -1862 -712
rect -1834 -740 -1796 -712
rect -1768 -740 -1730 -712
rect -1702 -740 -1664 -712
rect -1636 -740 -1598 -712
rect -1570 -740 -1532 -712
rect -1504 -740 -1466 -712
rect -1438 -740 -1400 -712
rect -1372 -740 -1334 -712
rect -1306 -740 -1268 -712
rect -1240 -740 -1202 -712
rect -1174 -740 -1136 -712
rect -1108 -740 -1070 -712
rect -1042 -740 -1004 -712
rect -976 -740 -938 -712
rect -910 -740 -872 -712
rect -844 -740 -806 -712
rect -778 -740 -740 -712
rect -712 -740 -674 -712
rect -646 -740 -608 -712
rect -580 -740 -542 -712
rect -514 -740 -476 -712
rect -448 -740 -410 -712
rect -382 -740 -344 -712
rect -316 -740 -278 -712
rect -250 -740 -212 -712
rect -184 -740 -146 -712
rect -118 -740 -80 -712
rect -52 -740 -14 -712
rect 14 -740 52 -712
rect 80 -740 118 -712
rect 146 -740 184 -712
rect 212 -740 250 -712
rect 278 -740 316 -712
rect 344 -740 382 -712
rect 410 -740 448 -712
rect 476 -740 514 -712
rect 542 -740 580 -712
rect 608 -740 646 -712
rect 674 -740 712 -712
rect 740 -740 778 -712
rect 806 -740 844 -712
rect 872 -740 910 -712
rect 938 -740 976 -712
rect 1004 -740 1042 -712
rect 1070 -740 1108 -712
rect 1136 -740 1174 -712
rect 1202 -740 1240 -712
rect 1268 -740 1306 -712
rect 1334 -740 1372 -712
rect 1400 -740 1438 -712
rect 1466 -740 1504 -712
rect 1532 -740 1570 -712
rect 1598 -740 1636 -712
rect 1664 -740 1702 -712
rect 1730 -740 1768 -712
rect 1796 -740 1834 -712
rect 1862 -740 1900 -712
rect 1928 -740 1966 -712
rect 1994 -740 2032 -712
rect 2060 -740 2098 -712
rect 2126 -740 2164 -712
rect 2192 -740 2230 -712
rect 2258 -740 2296 -712
rect 2324 -740 2362 -712
rect 2390 -740 2428 -712
rect 2456 -740 2494 -712
rect 2522 -740 2560 -712
rect 2588 -740 2626 -712
rect 2654 -740 2692 -712
rect 2720 -740 2758 -712
rect 2786 -740 2824 -712
rect 2852 -740 2890 -712
rect 2918 -740 2956 -712
rect 2984 -740 3022 -712
rect 3050 -740 3088 -712
rect 3116 -740 3154 -712
rect 3182 -740 3220 -712
rect 3248 -740 3286 -712
rect 3314 -740 3352 -712
rect 3380 -740 3418 -712
rect 3446 -740 3484 -712
rect 3512 -740 3550 -712
rect 3578 -740 3616 -712
rect 3644 -740 3682 -712
rect 3710 -740 3748 -712
rect 3776 -740 3814 -712
rect 3842 -740 3880 -712
rect 3908 -740 3946 -712
rect 3974 -740 4012 -712
rect 4040 -740 4078 -712
rect 4106 -740 4144 -712
rect 4172 -740 4210 -712
rect 4238 -740 4276 -712
rect 4304 -740 4342 -712
rect 4370 -740 4408 -712
rect 4436 -740 4474 -712
rect 4502 -740 4540 -712
rect 4568 -740 4573 -712
rect -4573 -745 4573 -740
<< end >>
