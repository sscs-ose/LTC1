magic
tech gf180mcuC
magscale 1 10
timestamp 1694582263
<< nwell >>
rect -442 -398 442 398
<< pmos >>
rect -268 68 -212 268
rect -108 68 -52 268
rect 52 68 108 268
rect 212 68 268 268
rect -268 -268 -212 -68
rect -108 -268 -52 -68
rect 52 -268 108 -68
rect 212 -268 268 -68
<< pdiff >>
rect -356 255 -268 268
rect -356 81 -343 255
rect -297 81 -268 255
rect -356 68 -268 81
rect -212 255 -108 268
rect -212 81 -183 255
rect -137 81 -108 255
rect -212 68 -108 81
rect -52 255 52 268
rect -52 81 -23 255
rect 23 81 52 255
rect -52 68 52 81
rect 108 255 212 268
rect 108 81 137 255
rect 183 81 212 255
rect 108 68 212 81
rect 268 255 356 268
rect 268 81 297 255
rect 343 81 356 255
rect 268 68 356 81
rect -356 -81 -268 -68
rect -356 -255 -343 -81
rect -297 -255 -268 -81
rect -356 -268 -268 -255
rect -212 -81 -108 -68
rect -212 -255 -183 -81
rect -137 -255 -108 -81
rect -212 -268 -108 -255
rect -52 -81 52 -68
rect -52 -255 -23 -81
rect 23 -255 52 -81
rect -52 -268 52 -255
rect 108 -81 212 -68
rect 108 -255 137 -81
rect 183 -255 212 -81
rect 108 -268 212 -255
rect 268 -81 356 -68
rect 268 -255 297 -81
rect 343 -255 356 -81
rect 268 -268 356 -255
<< pdiffc >>
rect -343 81 -297 255
rect -183 81 -137 255
rect -23 81 23 255
rect 137 81 183 255
rect 297 81 343 255
rect -343 -255 -297 -81
rect -183 -255 -137 -81
rect -23 -255 23 -81
rect 137 -255 183 -81
rect 297 -255 343 -81
<< polysilicon >>
rect -268 268 -212 312
rect -108 268 -52 312
rect 52 268 108 312
rect 212 268 268 312
rect -268 24 -212 68
rect -108 24 -52 68
rect 52 24 108 68
rect 212 24 268 68
rect -268 -68 -212 -24
rect -108 -68 -52 -24
rect 52 -68 108 -24
rect 212 -68 268 -24
rect -268 -312 -212 -268
rect -108 -312 -52 -268
rect 52 -312 108 -268
rect 212 -312 268 -268
<< metal1 >>
rect -343 255 -297 266
rect -343 70 -297 81
rect -183 255 -137 266
rect -183 70 -137 81
rect -23 255 23 266
rect -23 70 23 81
rect 137 255 183 266
rect 137 70 183 81
rect 297 255 343 266
rect 297 70 343 81
rect -343 -81 -297 -70
rect -343 -266 -297 -255
rect -183 -81 -137 -70
rect -183 -266 -137 -255
rect -23 -81 23 -70
rect -23 -266 23 -255
rect 137 -81 183 -70
rect 137 -266 183 -255
rect 297 -81 343 -70
rect 297 -266 343 -255
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 1 l 0.280 m 2 nf 4 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
