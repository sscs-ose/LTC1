* NGSPICE file created from OR_2_In_Layout_flat.ext - technology: gf180mcuC

.subckt OR_2_Input_PEX VDD A B OUT VSS
X0 VDD A.t0 a_86_440# VDD.t3 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X1 a_86_440# B.t0 a_390_68# VDD.t6 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X2 VDD a_390_68# OUT.t1 VDD.t7 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X3 a_390_68# A.t1 VSS.t1 VSS.t0 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X4 a_86_440# A.t2 VDD.t2 VDD.t1 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X5 a_390_68# B.t1 a_86_440# VDD.t0 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X6 OUT a_390_68# VSS.t6 VSS.t5 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X7 VSS B.t2 a_390_68# VSS.t2 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
R0 A.n0 A.t0 36.5005
R1 A.n2 A.n1 18.2505
R2 A.n1 A.t1 16.0344
R3 A.n0 A.t2 15.6434
R4 A.n1 A.n0 8.73443
R5 A A.n2 8.0005
R6 A A.n2 8.0005
R7 VDD.n11 VDD.t6 82.9108
R8 VDD.n19 VDD.t3 77.8347
R9 VDD.n2 VDD.t7 75.7026
R10 VDD.n23 VDD.t1 33.8415
R11 VDD.n29 VDD.t0 13.5369
R12 VDD.n1 VDD.n0 4.88224
R13 VDD.n4 VDD.n3 3.1505
R14 VDD.n7 VDD.n6 3.1505
R15 VDD.n6 VDD.n5 3.1505
R16 VDD.n10 VDD.n9 3.1505
R17 VDD.n9 VDD.n8 3.1505
R18 VDD.n13 VDD.n12 3.1505
R19 VDD.n12 VDD.n11 3.1505
R20 VDD.n16 VDD.n15 3.1505
R21 VDD.n15 VDD.n14 3.1505
R22 VDD.n31 VDD.n30 3.1505
R23 VDD.n30 VDD.n29 3.1505
R24 VDD.n28 VDD.n27 3.1505
R25 VDD.n27 VDD.n26 3.1505
R26 VDD.n25 VDD.n24 3.1505
R27 VDD.n24 VDD.n23 3.1505
R28 VDD.n20 VDD.n19 3.1505
R29 VDD.n22 VDD.n18 3.06224
R30 VDD.n21 VDD.n20 1.87197
R31 VDD.n18 VDD.t2 1.8205
R32 VDD.n18 VDD.n17 1.8205
R33 VDD.n22 VDD.n21 0.593718
R34 VDD.n3 VDD.n2 0.150506
R35 VDD.n16 VDD.n13 0.0864821
R36 VDD.n7 VDD.n4 0.0760357
R37 VDD.n10 VDD.n7 0.0760357
R38 VDD.n13 VDD.n10 0.0760357
R39 VDD.n31 VDD.n28 0.0760357
R40 VDD.n28 VDD.n25 0.0760357
R41 VDD.n25 VDD.n22 0.0487143
R42 VDD VDD.n16 0.0382679
R43 VDD VDD.n31 0.0382679
R44 VDD.n4 VDD.n1 0.0302321
R45 B.n1 B.t2 63.6148
R46 B.n0 B.t0 36.5005
R47 B.t2 B.n0 32.0684
R48 B.n0 B.t1 15.6434
R49 B B.n1 8.0005
R50 B B.n1 8.0005
R51 OUT.n1 OUT.n0 6.93911
R52 OUT.n1 OUT.t1 4.80398
R53 OUT OUT.n1 0.327239
R54 VSS.n6 VSS.t2 277.728
R55 VSS.n2 VSS.t5 112.273
R56 VSS.n11 VSS.t0 112.273
R57 VSS.n10 VSS.t1 6.91182
R58 VSS.n5 VSS.n1 3.6318
R59 VSS.n1 VSS.t6 3.2765
R60 VSS.n1 VSS.n0 3.2765
R61 VSS.n10 VSS.n9 2.6005
R62 VSS.n3 VSS.n2 2.6005
R63 VSS.n8 VSS.n7 2.6005
R64 VSS.n7 VSS.n6 2.6005
R65 VSS.n16 VSS.n15 2.6005
R66 VSS.n15 VSS.n14 2.6005
R67 VSS.n13 VSS.n12 2.6005
R68 VSS.n12 VSS.n11 2.6005
R69 VSS.n4 VSS.n3 1.64943
R70 VSS.n5 VSS.n4 0.532617
R71 VSS.n16 VSS.n13 0.0760357
R72 VSS.n13 VSS.n10 0.0760357
R73 VSS VSS.n16 0.0446964
R74 VSS VSS.n8 0.0318393
R75 VSS.n8 VSS.n5 0.0270179
C0 A VDD 0.234f
C1 A B 0.0842f
C2 OUT VDD 0.177f
C3 OUT B 0.00407f
C4 a_86_440# a_390_68# 0.293f
C5 A a_86_440# 0.208f
C6 B VDD 0.204f
C7 OUT a_86_440# 0.121f
C8 A a_390_68# 0.0208f
C9 OUT a_390_68# 0.119f
C10 VDD a_86_440# 0.792f
C11 B a_86_440# 0.0369f
C12 VDD a_390_68# 0.182f
C13 B a_390_68# 0.104f
.ends

