magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2083 -2083 4701 4911
<< isosubstrate >>
rect 1385 -83 2701 2911
<< nwell >>
rect -83 1213 1045 2911
rect 1385 1213 2701 2911
<< polysilicon >>
rect 286 914 426 1914
rect 530 914 670 1914
rect 1913 1213 2053 1314
rect 1697 1002 2053 1213
rect 1913 914 2053 1002
rect 2157 914 2297 1314
<< metal1 >>
rect 79 2749 165 2817
rect 196 1958 272 2787
rect 440 1794 516 2558
rect 684 1958 760 2787
rect 797 2749 883 2817
rect 1547 2749 1633 2817
rect 440 1718 760 1794
rect 684 1197 760 1718
rect 1823 1197 1899 2558
rect 2067 1358 2143 2787
rect 2453 2749 2539 2817
rect 684 1019 1773 1197
rect 1823 1019 2261 1197
rect 79 11 165 79
rect 196 42 272 870
rect 684 270 760 1019
rect 1823 270 1899 1019
rect 797 11 883 79
rect 1547 11 1633 79
rect 2067 39 2143 870
rect 2311 270 2387 2558
rect 2453 11 2539 79
use M1_NWELL_CDNS_40661953145223  M1_NWELL_CDNS_40661953145223_0
timestamp 1713338890
transform 1 0 45 0 1 2078
box -128 -833 128 833
use M1_NWELL_CDNS_40661953145223  M1_NWELL_CDNS_40661953145223_1
timestamp 1713338890
transform 1 0 917 0 1 2078
box -128 -833 128 833
use M1_NWELL_CDNS_40661953145223  M1_NWELL_CDNS_40661953145223_2
timestamp 1713338890
transform 1 0 1513 0 1 2078
box -128 -833 128 833
use M1_NWELL_CDNS_40661953145223  M1_NWELL_CDNS_40661953145223_3
timestamp 1713338890
transform 1 0 2573 0 1 2078
box -128 -833 128 833
use M1_NWELL_CDNS_40661953145225  M1_NWELL_CDNS_40661953145225_0
timestamp 1713338890
transform 1 0 2043 0 1 2783
box -504 -128 504 128
use M1_NWELL_CDNS_40661953145272  M1_NWELL_CDNS_40661953145272_0
timestamp 1713338890
transform 1 0 481 0 1 2783
box -410 -128 410 128
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_0
timestamp 1713338890
transform -1 0 600 0 1 1467
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_1
timestamp 1713338890
transform -1 0 356 0 1 1467
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_2
timestamp 1713338890
transform 1 0 1739 0 1 1108
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_3
timestamp 1713338890
transform 1 0 2219 0 1 1108
box -42 -89 42 89
use M1_PSUB_CDNS_69033583165609  M1_PSUB_CDNS_69033583165609_0
timestamp 1713338890
transform 1 0 45 0 -1 515
box -45 -515 45 515
use M1_PSUB_CDNS_69033583165609  M1_PSUB_CDNS_69033583165609_1
timestamp 1713338890
transform 1 0 2573 0 -1 515
box -45 -515 45 515
use M1_PSUB_CDNS_69033583165611  M1_PSUB_CDNS_69033583165611_0
timestamp 1713338890
transform 1 0 917 0 -1 468
box -45 -468 45 468
use M1_PSUB_CDNS_69033583165611  M1_PSUB_CDNS_69033583165611_1
timestamp 1713338890
transform 1 0 1513 0 -1 468
box -45 -468 45 468
use M1_PSUB_CDNS_69033583165612  M1_PSUB_CDNS_69033583165612_0
timestamp 1713338890
transform 1 0 2043 0 -1 45
box -421 -45 421 45
use M1_PSUB_CDNS_69033583165694  M1_PSUB_CDNS_69033583165694_0
timestamp 1713338890
transform 1 0 481 0 -1 45
box -327 -45 327 45
use nmos_6p0_CDNS_4066195314511  nmos_6p0_CDNS_4066195314511_0
timestamp 1713338890
transform 1 0 286 0 1 270
box -88 -44 228 644
use nmos_6p0_CDNS_4066195314511  nmos_6p0_CDNS_4066195314511_1
timestamp 1713338890
transform 1 0 530 0 1 270
box -88 -44 228 644
use nmos_6p0_CDNS_4066195314511  nmos_6p0_CDNS_4066195314511_2
timestamp 1713338890
transform 1 0 1913 0 1 270
box -88 -44 228 644
use nmos_6p0_CDNS_4066195314511  nmos_6p0_CDNS_4066195314511_3
timestamp 1713338890
transform 1 0 2157 0 1 270
box -88 -44 228 644
use pmos_6p0_CDNS_4066195314512  pmos_6p0_CDNS_4066195314512_0
timestamp 1713338890
transform 1 0 286 0 1 1958
box -208 -120 348 720
use pmos_6p0_CDNS_4066195314512  pmos_6p0_CDNS_4066195314512_1
timestamp 1713338890
transform -1 0 670 0 1 1958
box -208 -120 348 720
use pmos_6p0_CDNS_4066195314513  pmos_6p0_CDNS_4066195314513_0
timestamp 1713338890
transform 1 0 1913 0 1 1358
box -208 -120 348 1320
use pmos_6p0_CDNS_4066195314513  pmos_6p0_CDNS_4066195314513_1
timestamp 1713338890
transform 1 0 2157 0 1 1358
box -208 -120 348 1320
<< labels >>
rlabel metal1 s 92 2788 92 2788 4 VDD
port 1 nsew
rlabel metal1 s 349 1468 349 1468 4 OE
port 2 nsew
rlabel metal1 s 2254 2788 2254 2788 4 DVDD
port 3 nsew
rlabel metal1 s 2245 45 2245 45 4 DVSS
port 4 nsew
rlabel metal1 s 604 1468 604 1468 4 A
port 5 nsew
rlabel metal1 s 2349 1100 2349 1100 4 AB
port 6 nsew
rlabel metal1 s 263 45 263 45 4 VSS
port 7 nsew
<< end >>
