magic
tech gf180mcuC
magscale 1 10
timestamp 1699111554
<< nwell >>
rect -3024 -2040 3024 2040
<< nsubdiff >>
rect -3000 2003 3000 2016
rect -3000 1957 -2884 2003
rect 2884 1957 3000 2003
rect -3000 1944 3000 1957
rect -3000 1900 -2928 1944
rect -3000 -1900 -2987 1900
rect -2941 -1900 -2928 1900
rect 2928 1900 3000 1944
rect -3000 -1944 -2928 -1900
rect 2928 -1900 2941 1900
rect 2987 -1900 3000 1900
rect 2928 -1944 3000 -1900
rect -3000 -1957 3000 -1944
rect -3000 -2003 -2884 -1957
rect 2884 -2003 3000 -1957
rect -3000 -2016 3000 -2003
<< nsubdiffcont >>
rect -2884 1957 2884 2003
rect -2987 -1900 -2941 1900
rect 2941 -1900 2987 1900
rect -2884 -2003 2884 -1957
<< polysilicon >>
rect -2840 1843 -2440 1856
rect -2840 1797 -2827 1843
rect -2453 1797 -2440 1843
rect -2840 1754 -2440 1797
rect -2840 111 -2440 154
rect -2840 65 -2827 111
rect -2453 65 -2440 111
rect -2840 52 -2440 65
rect -2360 1843 -1960 1856
rect -2360 1797 -2347 1843
rect -1973 1797 -1960 1843
rect -2360 1754 -1960 1797
rect -2360 111 -1960 154
rect -2360 65 -2347 111
rect -1973 65 -1960 111
rect -2360 52 -1960 65
rect -1880 1843 -1480 1856
rect -1880 1797 -1867 1843
rect -1493 1797 -1480 1843
rect -1880 1754 -1480 1797
rect -1880 111 -1480 154
rect -1880 65 -1867 111
rect -1493 65 -1480 111
rect -1880 52 -1480 65
rect -1400 1843 -1000 1856
rect -1400 1797 -1387 1843
rect -1013 1797 -1000 1843
rect -1400 1754 -1000 1797
rect -1400 111 -1000 154
rect -1400 65 -1387 111
rect -1013 65 -1000 111
rect -1400 52 -1000 65
rect -920 1843 -520 1856
rect -920 1797 -907 1843
rect -533 1797 -520 1843
rect -920 1754 -520 1797
rect -920 111 -520 154
rect -920 65 -907 111
rect -533 65 -520 111
rect -920 52 -520 65
rect -440 1843 -40 1856
rect -440 1797 -427 1843
rect -53 1797 -40 1843
rect -440 1754 -40 1797
rect -440 111 -40 154
rect -440 65 -427 111
rect -53 65 -40 111
rect -440 52 -40 65
rect 40 1843 440 1856
rect 40 1797 53 1843
rect 427 1797 440 1843
rect 40 1754 440 1797
rect 40 111 440 154
rect 40 65 53 111
rect 427 65 440 111
rect 40 52 440 65
rect 520 1843 920 1856
rect 520 1797 533 1843
rect 907 1797 920 1843
rect 520 1754 920 1797
rect 520 111 920 154
rect 520 65 533 111
rect 907 65 920 111
rect 520 52 920 65
rect 1000 1843 1400 1856
rect 1000 1797 1013 1843
rect 1387 1797 1400 1843
rect 1000 1754 1400 1797
rect 1000 111 1400 154
rect 1000 65 1013 111
rect 1387 65 1400 111
rect 1000 52 1400 65
rect 1480 1843 1880 1856
rect 1480 1797 1493 1843
rect 1867 1797 1880 1843
rect 1480 1754 1880 1797
rect 1480 111 1880 154
rect 1480 65 1493 111
rect 1867 65 1880 111
rect 1480 52 1880 65
rect 1960 1843 2360 1856
rect 1960 1797 1973 1843
rect 2347 1797 2360 1843
rect 1960 1754 2360 1797
rect 1960 111 2360 154
rect 1960 65 1973 111
rect 2347 65 2360 111
rect 1960 52 2360 65
rect 2440 1843 2840 1856
rect 2440 1797 2453 1843
rect 2827 1797 2840 1843
rect 2440 1754 2840 1797
rect 2440 111 2840 154
rect 2440 65 2453 111
rect 2827 65 2840 111
rect 2440 52 2840 65
rect -2840 -65 -2440 -52
rect -2840 -111 -2827 -65
rect -2453 -111 -2440 -65
rect -2840 -154 -2440 -111
rect -2840 -1797 -2440 -1754
rect -2840 -1843 -2827 -1797
rect -2453 -1843 -2440 -1797
rect -2840 -1856 -2440 -1843
rect -2360 -65 -1960 -52
rect -2360 -111 -2347 -65
rect -1973 -111 -1960 -65
rect -2360 -154 -1960 -111
rect -2360 -1797 -1960 -1754
rect -2360 -1843 -2347 -1797
rect -1973 -1843 -1960 -1797
rect -2360 -1856 -1960 -1843
rect -1880 -65 -1480 -52
rect -1880 -111 -1867 -65
rect -1493 -111 -1480 -65
rect -1880 -154 -1480 -111
rect -1880 -1797 -1480 -1754
rect -1880 -1843 -1867 -1797
rect -1493 -1843 -1480 -1797
rect -1880 -1856 -1480 -1843
rect -1400 -65 -1000 -52
rect -1400 -111 -1387 -65
rect -1013 -111 -1000 -65
rect -1400 -154 -1000 -111
rect -1400 -1797 -1000 -1754
rect -1400 -1843 -1387 -1797
rect -1013 -1843 -1000 -1797
rect -1400 -1856 -1000 -1843
rect -920 -65 -520 -52
rect -920 -111 -907 -65
rect -533 -111 -520 -65
rect -920 -154 -520 -111
rect -920 -1797 -520 -1754
rect -920 -1843 -907 -1797
rect -533 -1843 -520 -1797
rect -920 -1856 -520 -1843
rect -440 -65 -40 -52
rect -440 -111 -427 -65
rect -53 -111 -40 -65
rect -440 -154 -40 -111
rect -440 -1797 -40 -1754
rect -440 -1843 -427 -1797
rect -53 -1843 -40 -1797
rect -440 -1856 -40 -1843
rect 40 -65 440 -52
rect 40 -111 53 -65
rect 427 -111 440 -65
rect 40 -154 440 -111
rect 40 -1797 440 -1754
rect 40 -1843 53 -1797
rect 427 -1843 440 -1797
rect 40 -1856 440 -1843
rect 520 -65 920 -52
rect 520 -111 533 -65
rect 907 -111 920 -65
rect 520 -154 920 -111
rect 520 -1797 920 -1754
rect 520 -1843 533 -1797
rect 907 -1843 920 -1797
rect 520 -1856 920 -1843
rect 1000 -65 1400 -52
rect 1000 -111 1013 -65
rect 1387 -111 1400 -65
rect 1000 -154 1400 -111
rect 1000 -1797 1400 -1754
rect 1000 -1843 1013 -1797
rect 1387 -1843 1400 -1797
rect 1000 -1856 1400 -1843
rect 1480 -65 1880 -52
rect 1480 -111 1493 -65
rect 1867 -111 1880 -65
rect 1480 -154 1880 -111
rect 1480 -1797 1880 -1754
rect 1480 -1843 1493 -1797
rect 1867 -1843 1880 -1797
rect 1480 -1856 1880 -1843
rect 1960 -65 2360 -52
rect 1960 -111 1973 -65
rect 2347 -111 2360 -65
rect 1960 -154 2360 -111
rect 1960 -1797 2360 -1754
rect 1960 -1843 1973 -1797
rect 2347 -1843 2360 -1797
rect 1960 -1856 2360 -1843
rect 2440 -65 2840 -52
rect 2440 -111 2453 -65
rect 2827 -111 2840 -65
rect 2440 -154 2840 -111
rect 2440 -1797 2840 -1754
rect 2440 -1843 2453 -1797
rect 2827 -1843 2840 -1797
rect 2440 -1856 2840 -1843
<< polycontact >>
rect -2827 1797 -2453 1843
rect -2827 65 -2453 111
rect -2347 1797 -1973 1843
rect -2347 65 -1973 111
rect -1867 1797 -1493 1843
rect -1867 65 -1493 111
rect -1387 1797 -1013 1843
rect -1387 65 -1013 111
rect -907 1797 -533 1843
rect -907 65 -533 111
rect -427 1797 -53 1843
rect -427 65 -53 111
rect 53 1797 427 1843
rect 53 65 427 111
rect 533 1797 907 1843
rect 533 65 907 111
rect 1013 1797 1387 1843
rect 1013 65 1387 111
rect 1493 1797 1867 1843
rect 1493 65 1867 111
rect 1973 1797 2347 1843
rect 1973 65 2347 111
rect 2453 1797 2827 1843
rect 2453 65 2827 111
rect -2827 -111 -2453 -65
rect -2827 -1843 -2453 -1797
rect -2347 -111 -1973 -65
rect -2347 -1843 -1973 -1797
rect -1867 -111 -1493 -65
rect -1867 -1843 -1493 -1797
rect -1387 -111 -1013 -65
rect -1387 -1843 -1013 -1797
rect -907 -111 -533 -65
rect -907 -1843 -533 -1797
rect -427 -111 -53 -65
rect -427 -1843 -53 -1797
rect 53 -111 427 -65
rect 53 -1843 427 -1797
rect 533 -111 907 -65
rect 533 -1843 907 -1797
rect 1013 -111 1387 -65
rect 1013 -1843 1387 -1797
rect 1493 -111 1867 -65
rect 1493 -1843 1867 -1797
rect 1973 -111 2347 -65
rect 1973 -1843 2347 -1797
rect 2453 -111 2827 -65
rect 2453 -1843 2827 -1797
<< ppolyres >>
rect -2840 154 -2440 1754
rect -2360 154 -1960 1754
rect -1880 154 -1480 1754
rect -1400 154 -1000 1754
rect -920 154 -520 1754
rect -440 154 -40 1754
rect 40 154 440 1754
rect 520 154 920 1754
rect 1000 154 1400 1754
rect 1480 154 1880 1754
rect 1960 154 2360 1754
rect 2440 154 2840 1754
rect -2840 -1754 -2440 -154
rect -2360 -1754 -1960 -154
rect -1880 -1754 -1480 -154
rect -1400 -1754 -1000 -154
rect -920 -1754 -520 -154
rect -440 -1754 -40 -154
rect 40 -1754 440 -154
rect 520 -1754 920 -154
rect 1000 -1754 1400 -154
rect 1480 -1754 1880 -154
rect 1960 -1754 2360 -154
rect 2440 -1754 2840 -154
<< metal1 >>
rect -2987 1957 -2884 2003
rect 2884 1957 2987 2003
rect -2987 1900 -2941 1957
rect 2941 1900 2987 1957
rect -2838 1797 -2827 1843
rect -2453 1797 -2442 1843
rect -2358 1797 -2347 1843
rect -1973 1797 -1962 1843
rect -1878 1797 -1867 1843
rect -1493 1797 -1482 1843
rect -1398 1797 -1387 1843
rect -1013 1797 -1002 1843
rect -918 1797 -907 1843
rect -533 1797 -522 1843
rect -438 1797 -427 1843
rect -53 1797 -42 1843
rect 42 1797 53 1843
rect 427 1797 438 1843
rect 522 1797 533 1843
rect 907 1797 918 1843
rect 1002 1797 1013 1843
rect 1387 1797 1398 1843
rect 1482 1797 1493 1843
rect 1867 1797 1878 1843
rect 1962 1797 1973 1843
rect 2347 1797 2358 1843
rect 2442 1797 2453 1843
rect 2827 1797 2838 1843
rect -2838 65 -2827 111
rect -2453 65 -2442 111
rect -2358 65 -2347 111
rect -1973 65 -1962 111
rect -1878 65 -1867 111
rect -1493 65 -1482 111
rect -1398 65 -1387 111
rect -1013 65 -1002 111
rect -918 65 -907 111
rect -533 65 -522 111
rect -438 65 -427 111
rect -53 65 -42 111
rect 42 65 53 111
rect 427 65 438 111
rect 522 65 533 111
rect 907 65 918 111
rect 1002 65 1013 111
rect 1387 65 1398 111
rect 1482 65 1493 111
rect 1867 65 1878 111
rect 1962 65 1973 111
rect 2347 65 2358 111
rect 2442 65 2453 111
rect 2827 65 2838 111
rect -2838 -111 -2827 -65
rect -2453 -111 -2442 -65
rect -2358 -111 -2347 -65
rect -1973 -111 -1962 -65
rect -1878 -111 -1867 -65
rect -1493 -111 -1482 -65
rect -1398 -111 -1387 -65
rect -1013 -111 -1002 -65
rect -918 -111 -907 -65
rect -533 -111 -522 -65
rect -438 -111 -427 -65
rect -53 -111 -42 -65
rect 42 -111 53 -65
rect 427 -111 438 -65
rect 522 -111 533 -65
rect 907 -111 918 -65
rect 1002 -111 1013 -65
rect 1387 -111 1398 -65
rect 1482 -111 1493 -65
rect 1867 -111 1878 -65
rect 1962 -111 1973 -65
rect 2347 -111 2358 -65
rect 2442 -111 2453 -65
rect 2827 -111 2838 -65
rect -2838 -1843 -2827 -1797
rect -2453 -1843 -2442 -1797
rect -2358 -1843 -2347 -1797
rect -1973 -1843 -1962 -1797
rect -1878 -1843 -1867 -1797
rect -1493 -1843 -1482 -1797
rect -1398 -1843 -1387 -1797
rect -1013 -1843 -1002 -1797
rect -918 -1843 -907 -1797
rect -533 -1843 -522 -1797
rect -438 -1843 -427 -1797
rect -53 -1843 -42 -1797
rect 42 -1843 53 -1797
rect 427 -1843 438 -1797
rect 522 -1843 533 -1797
rect 907 -1843 918 -1797
rect 1002 -1843 1013 -1797
rect 1387 -1843 1398 -1797
rect 1482 -1843 1493 -1797
rect 1867 -1843 1878 -1797
rect 1962 -1843 1973 -1797
rect 2347 -1843 2358 -1797
rect 2442 -1843 2453 -1797
rect 2827 -1843 2838 -1797
rect -2987 -1957 -2941 -1900
rect 2941 -1957 2987 -1900
rect -2987 -2003 -2884 -1957
rect 2884 -2003 2987 -1957
<< properties >>
string FIXED_BBOX -2964 -1980 2964 1980
string gencell ppolyf_u
string library gf180mcu
string parameters w 2.0 l 8.0 m 2 nx 12 wmin 0.80 lmin 1.00 rho 315 val 1.305k dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1
<< end >>
