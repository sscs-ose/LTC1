* NGSPICE file created from nmos_3p3_H9QVWA_flat.ext - technology: gf180mcuC

.subckt nmos_3p3_H9QVWA_flat B C OUT VDD VSS A
X0 OUT a_86_n207# VDD.t15 VDD.t14 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X1 VDD B.t0 a_86_n207# VDD.t20 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X2 VDD.t7 VDD.t5 VDD.t7 VDD.t6 pfet_03v3 ad=0 pd=0 as=89.8f ps=0.92u w=0.25u l=0.28u
X3 VDD C.t0 a_86_n207# VDD.t23 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X4 a_738_n196# B.t1 a_234_n196# VSS.t14 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X5 VSS C.t1 a_738_n196# VSS.t8 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X6 a_86_n207# B.t2 VDD.t17 VDD.t16 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X7 a_738_n196# C.t2 VSS.t7 VSS.t6 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X8 VDD a_86_n207# OUT.t0 VDD.t11 pfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X9 VSS C.t3 a_738_n196# VSS.t3 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X10 OUT a_86_n207# VSS.t2 VSS.t1 nfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X11 a_234_n196# A.t0 a_86_n207# VSS.t0 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X12 VDD A.t1 a_86_n207# VDD.t8 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X13 a_86_n207# A.t2 a_234_n196# VSS.t11 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X14 a_234_n196# B.t3 a_738_n196# VSS.t13 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X15 a_86_n207# C.t4 VDD.t19 VDD.t18 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X16 a_234_n196# A.t3 a_86_n207# VSS.t15 nfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
X17 a_738_n196# B.t4 a_234_n196# VSS.t12 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X18 a_86_n207# A.t4 VDD.t1 VDD.t0 pfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
X19 VDD.t4 VDD.t2 VDD.t4 VDD.t3 pfet_03v3 ad=0 pd=0 as=89.8f ps=0.92u w=0.25u l=0.28u
R0 VDD.n12 VDD.t14 96.0457
R1 VDD.n22 VDD.t23 84.7463
R2 VDD.n52 VDD.t3 73.4468
R3 VDD.n43 VDD.t16 62.1474
R4 VDD.n33 VDD.t0 53.828
R5 VDD.n39 VDD.t8 47.0815
R6 VDD.n49 VDD.t20 35.782
R7 VDD.n56 VDD.t18 24.4826
R8 VDD.n29 VDD.t2 18.4701
R9 VDD.n3 VDD.t5 18.4701
R10 VDD.n15 VDD.t6 13.1832
R11 VDD.n32 VDD.t1 9.36138
R12 VDD.n5 VDD.n4 9.36138
R13 VDD.n58 VDD.n57 8.72358
R14 VDD.n31 VDD.n30 6.3005
R15 VDD.n31 VDD.t17 6.3005
R16 VDD.n28 VDD.n27 6.3005
R17 VDD.n26 VDD.t4 6.3005
R18 VDD.n26 VDD.t19 6.3005
R19 VDD.n2 VDD.n1 6.3005
R20 VDD.n0 VDD.t7 6.3005
R21 VDD.n0 VDD.t15 6.3005
R22 VDD.n6 VDD.t11 4.86375
R23 VDD.n8 VDD.n7 3.1505
R24 VDD.n11 VDD.n10 3.1505
R25 VDD.n10 VDD.n9 3.1505
R26 VDD.n14 VDD.n13 3.1505
R27 VDD.n13 VDD.n12 3.1505
R28 VDD.n17 VDD.n16 3.1505
R29 VDD.n16 VDD.n15 3.1505
R30 VDD.n21 VDD.n20 3.1505
R31 VDD.n20 VDD.n19 3.1505
R32 VDD.n24 VDD.n23 3.1505
R33 VDD.n23 VDD.n22 3.1505
R34 VDD.n57 VDD.n25 3.1505
R35 VDD.n57 VDD.n56 3.1505
R36 VDD.n61 VDD.n60 3.1505
R37 VDD.n60 VDD.n59 3.1505
R38 VDD.n54 VDD.n53 3.1505
R39 VDD.n53 VDD.n52 3.1505
R40 VDD.n51 VDD.n50 3.1505
R41 VDD.n50 VDD.n49 3.1505
R42 VDD.n48 VDD.n47 3.1505
R43 VDD.n47 VDD.n46 3.1505
R44 VDD.n45 VDD.n44 3.1505
R45 VDD.n44 VDD.n43 3.1505
R46 VDD.n41 VDD.n40 3.1505
R47 VDD.n40 VDD.n39 3.1505
R48 VDD.n38 VDD.n37 3.1505
R49 VDD.n37 VDD.n36 3.1505
R50 VDD.n35 VDD.n34 3.1505
R51 VDD.n42 VDD.n31 3.06138
R52 VDD.n29 VDD.n28 2.86655
R53 VDD.n29 VDD.n26 2.86655
R54 VDD.n3 VDD.n2 2.86655
R55 VDD.n3 VDD.n0 2.86655
R56 VDD.n55 VDD.n29 0.172674
R57 VDD.n18 VDD.n3 0.172674
R58 VDD.n60 VDD.n58 0.162038
R59 VDD.n7 VDD.n6 0.127116
R60 VDD.n34 VDD.n33 0.126872
R61 VDD.n11 VDD.n8 0.0975588
R62 VDD.n14 VDD.n11 0.0975588
R63 VDD.n17 VDD.n14 0.0975588
R64 VDD.n24 VDD.n21 0.0975588
R65 VDD.n25 VDD.n24 0.0975588
R66 VDD.n54 VDD.n51 0.0975588
R67 VDD.n51 VDD.n48 0.0975588
R68 VDD.n48 VDD.n45 0.0975588
R69 VDD.n41 VDD.n38 0.0975588
R70 VDD.n38 VDD.n35 0.0975588
R71 VDD VDD.n25 0.0957941
R72 VDD.n21 VDD.n18 0.0913824
R73 VDD.n8 VDD.n5 0.0737353
R74 VDD.n61 VDD.n55 0.0631471
R75 VDD.n42 VDD.n41 0.0525588
R76 VDD.n35 VDD.n32 0.0507941
R77 VDD.n45 VDD.n42 0.0455
R78 VDD.n55 VDD.n54 0.0349118
R79 VDD.n18 VDD.n17 0.00667647
R80 VDD VDD.n61 0.00226471
R81 OUT OUT.n2 8.97809
R82 OUT.n1 OUT.n0 6.3005
R83 OUT.n1 OUT.t0 6.3005
R84 OUT OUT.n1 3.24041
R85 B B.t2 89.0293
R86 B.n0 B.t1 35.4088
R87 B.t2 B.n2 34.0527
R88 B.n1 B.n0 25.7624
R89 B.n2 B.n1 22.2916
R90 B.n2 B.t0 11.3416
R91 B.n1 B.t4 9.64693
R92 B.n0 B.t3 3.25943
R93 C.t0 C.t4 45.3938
R94 C.t3 C.t0 43.2791
R95 C.n0 C.t1 35.6691
R96 C.n1 C.n0 25.6316
R97 C C.n1 21.1146
R98 C.n1 C.t3 10.038
R99 C.n0 C.t2 3.25943
R100 VSS.n10 VSS.t8 294.385
R101 VSS.n19 VSS.t3 259.058
R102 VSS.n44 VSS.t13 223.732
R103 VSS.n32 VSS.t0 188.406
R104 VSS.n28 VSS.t15 157.202
R105 VSS.n29 VSS.t11 153.081
R106 VSS.n38 VSS.t12 117.754
R107 VSS.n22 VSS.t14 82.428
R108 VSS.n13 VSS.t6 47.1019
R109 VSS.n5 VSS.t1 14.3592
R110 VSS.n45 VSS.n43 10.3113
R111 VSS.n1 VSS.n0 5.6705
R112 VSS.n1 VSS.t2 5.6705
R113 VSS.n3 VSS.n2 5.6705
R114 VSS.n3 VSS.t7 5.6705
R115 VSS.n4 VSS.n3 3.92833
R116 VSS.n4 VSS.n1 3.27094
R117 VSS.n9 VSS.n8 2.6005
R118 VSS.n8 VSS.n7 2.6005
R119 VSS.n12 VSS.n11 2.6005
R120 VSS.n11 VSS.n10 2.6005
R121 VSS.n15 VSS.n14 2.6005
R122 VSS.n14 VSS.n13 2.6005
R123 VSS.n18 VSS.n17 2.6005
R124 VSS.n17 VSS.n16 2.6005
R125 VSS.n21 VSS.n20 2.6005
R126 VSS.n20 VSS.n19 2.6005
R127 VSS.n24 VSS.n23 2.6005
R128 VSS.n23 VSS.n22 2.6005
R129 VSS.n42 VSS.n25 2.6005
R130 VSS.n42 VSS.n41 2.6005
R131 VSS.n46 VSS.n45 2.6005
R132 VSS.n45 VSS.n44 2.6005
R133 VSS.n40 VSS.n39 2.6005
R134 VSS.n39 VSS.n38 2.6005
R135 VSS.n37 VSS.n36 2.6005
R136 VSS.n36 VSS.n35 2.6005
R137 VSS.n34 VSS.n33 2.6005
R138 VSS.n33 VSS.n32 2.6005
R139 VSS.n31 VSS.n30 2.6005
R140 VSS.n30 VSS.n29 2.6005
R141 VSS.n27 VSS.n26 2.6005
R142 VSS.n6 VSS.n5 2.23602
R143 VSS.n28 VSS.n27 1.77403
R144 VSS.n31 VSS.n28 0.482318
R145 VSS.n6 VSS.n4 0.32137
R146 VSS.n12 VSS.n9 0.0975588
R147 VSS.n15 VSS.n12 0.0975588
R148 VSS.n18 VSS.n15 0.0975588
R149 VSS.n21 VSS.n18 0.0975588
R150 VSS.n24 VSS.n21 0.0975588
R151 VSS.n25 VSS.n24 0.0975588
R152 VSS.n46 VSS.n40 0.0975588
R153 VSS.n40 VSS.n37 0.0975588
R154 VSS.n37 VSS.n34 0.0975588
R155 VSS.n34 VSS.n31 0.0975588
R156 VSS VSS.n46 0.0966765
R157 VSS.n43 VSS.n42 0.0950946
R158 VSS.n9 VSS.n6 0.0216765
R159 VSS VSS.n25 0.00138235
R160 A.n1 A.t0 33.6616
R161 A.n0 A.t1 33.5692
R162 A.n2 A.n1 22.7116
R163 A.n3 A.n2 16.8166
R164 A.n0 A.t4 11.4719
R165 A.n1 A.t2 10.9505
R166 A.n2 A.t3 10.9505
R167 A A.n3 6.68888
R168 A.n3 A.n0 4.04157
C0 B a_234_n196# 0.0545f
C1 B a_86_n207# 0.0592f
C2 a_234_n196# C 0.457f
C3 a_86_n207# C 0.111f
C4 a_86_n207# a_234_n196# 0.475f
C5 VDD a_738_n196# 0.00358f
C6 VDD OUT 0.181f
C7 B a_738_n196# 0.0349f
C8 B OUT 6.31e-20
C9 C a_738_n196# 0.502f
C10 C OUT 0.00142f
C11 VDD A 0.331f
C12 a_234_n196# a_738_n196# 0.32f
C13 a_86_n207# a_738_n196# 0.285f
C14 a_86_n207# OUT 0.0793f
C15 B A 0.111f
C16 C A 0.0302f
C17 a_234_n196# A 0.0352f
C18 a_86_n207# A 0.192f
C19 B VDD 0.748f
C20 VDD C 0.311f
C21 OUT a_738_n196# 0.0134f
C22 VDD a_234_n196# 0.00684f
C23 VDD a_86_n207# 1.07f
C24 B C 0.0273f
.ends

