magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2032 11097 3032 71968
<< metal5 >>
rect 0 63600 1000 65000
rect 0 62000 1000 63400
rect 0 50800 1000 52200
rect 0 49200 1000 50600
use GF_NI_BRK5_0  GF_NI_BRK5_0_0
timestamp 1713338890
transform 1 0 0 0 1 0
box -32 13097 1032 69968
use M5_M4_CDNS_69033583165696  M5_M4_CDNS_69033583165696_0
timestamp 1713338890
transform 1 0 498 0 1 49894
box -354 -602 354 602
use M5_M4_CDNS_69033583165696  M5_M4_CDNS_69033583165696_1
timestamp 1713338890
transform 1 0 506 0 1 64300
box -354 -602 354 602
<< labels >>
rlabel metal5 s 498 64258 498 64258 4 VSS
port 1 nsew
rlabel metal5 s 510 50023 510 50023 4 VSS
port 1 nsew
rlabel metal4 s 510 50023 510 50023 4 VSS
port 1 nsew
rlabel metal4 s 498 64258 498 64258 4 VSS
port 1 nsew
rlabel metal3 s 498 64258 498 64258 4 VSS
port 1 nsew
rlabel metal3 s 510 50023 510 50023 4 VSS
port 1 nsew
rlabel metal5 s 498 62718 498 62718 4 VDD
port 2 nsew
rlabel metal5 s 498 51518 498 51518 4 VDD
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 1000 70000
<< end >>
