magic
tech gf180mcuC
magscale 1 10
timestamp 1694691102
<< nwell >>
rect -89 903 10119 5761
<< nsubdiff >>
rect -39 5698 10069 5715
rect -39 5648 -22 5698
rect 24 5652 76 5698
rect 122 5652 174 5698
rect 220 5652 272 5698
rect 318 5652 370 5698
rect 416 5652 468 5698
rect 514 5652 566 5698
rect 612 5652 664 5698
rect 710 5652 762 5698
rect 808 5652 860 5698
rect 906 5652 958 5698
rect 1004 5652 1056 5698
rect 1102 5652 1154 5698
rect 1200 5652 1252 5698
rect 1298 5652 1350 5698
rect 1396 5652 1448 5698
rect 1494 5652 1546 5698
rect 1592 5652 1644 5698
rect 1690 5652 1742 5698
rect 1788 5652 1840 5698
rect 1886 5652 1938 5698
rect 1984 5652 2036 5698
rect 2082 5652 2134 5698
rect 2180 5652 2232 5698
rect 2278 5652 2330 5698
rect 2376 5652 2428 5698
rect 2474 5652 2526 5698
rect 2572 5652 2624 5698
rect 2670 5652 2722 5698
rect 2768 5652 2820 5698
rect 2866 5652 2918 5698
rect 2964 5652 3016 5698
rect 3062 5652 3114 5698
rect 3160 5652 3212 5698
rect 3258 5652 3310 5698
rect 3356 5652 3408 5698
rect 3454 5652 3506 5698
rect 3552 5652 3604 5698
rect 3650 5652 3702 5698
rect 3748 5652 3800 5698
rect 3846 5652 3898 5698
rect 3944 5652 3996 5698
rect 4042 5652 4094 5698
rect 4140 5652 4192 5698
rect 4238 5652 4290 5698
rect 4336 5652 4388 5698
rect 4434 5652 4486 5698
rect 4532 5652 4584 5698
rect 4630 5652 4682 5698
rect 4728 5652 4780 5698
rect 4826 5652 4878 5698
rect 4924 5652 4976 5698
rect 5022 5652 5074 5698
rect 5120 5652 5172 5698
rect 5218 5652 5270 5698
rect 5316 5652 5368 5698
rect 5414 5652 5466 5698
rect 5512 5652 5564 5698
rect 5610 5652 5662 5698
rect 5708 5652 5760 5698
rect 5806 5652 5858 5698
rect 5904 5652 5956 5698
rect 6002 5652 6054 5698
rect 6100 5652 6152 5698
rect 6198 5652 6250 5698
rect 6296 5652 6348 5698
rect 6394 5652 6446 5698
rect 6492 5652 6544 5698
rect 6590 5652 6642 5698
rect 6688 5652 6740 5698
rect 6786 5652 6838 5698
rect 6884 5652 6936 5698
rect 6982 5652 7034 5698
rect 7080 5652 7132 5698
rect 7178 5652 7230 5698
rect 7276 5652 7328 5698
rect 7374 5652 7426 5698
rect 7472 5652 7524 5698
rect 7570 5652 7622 5698
rect 7668 5652 7720 5698
rect 7766 5652 7818 5698
rect 7864 5652 7916 5698
rect 7962 5652 8014 5698
rect 8060 5652 8112 5698
rect 8158 5652 8210 5698
rect 8256 5652 8308 5698
rect 8354 5652 8406 5698
rect 8452 5652 8504 5698
rect 8550 5652 8602 5698
rect 8648 5652 8700 5698
rect 8746 5652 8798 5698
rect 8844 5652 8896 5698
rect 8942 5652 8994 5698
rect 9040 5652 9092 5698
rect 9138 5652 9190 5698
rect 9236 5652 9288 5698
rect 9334 5652 9386 5698
rect 9432 5652 9484 5698
rect 9530 5652 9582 5698
rect 9628 5652 9680 5698
rect 9726 5652 9778 5698
rect 9824 5652 9876 5698
rect 9922 5652 10006 5698
rect 24 5648 10006 5652
rect 10052 5648 10069 5698
rect -39 5635 10069 5648
rect -39 5596 41 5635
rect -39 5550 -22 5596
rect 24 5550 41 5596
rect 9989 5596 10069 5635
rect -39 5498 41 5550
rect -39 5452 -22 5498
rect 24 5452 41 5498
rect -39 5400 41 5452
rect -39 5354 -22 5400
rect 24 5354 41 5400
rect -39 5302 41 5354
rect -39 5256 -22 5302
rect 24 5256 41 5302
rect -39 5204 41 5256
rect -39 5158 -22 5204
rect 24 5158 41 5204
rect -39 5106 41 5158
rect -39 5060 -22 5106
rect 24 5060 41 5106
rect -39 5008 41 5060
rect -39 4962 -22 5008
rect 24 4962 41 5008
rect -39 4910 41 4962
rect -39 4864 -22 4910
rect 24 4864 41 4910
rect -39 4812 41 4864
rect -39 4766 -22 4812
rect 24 4766 41 4812
rect -39 4714 41 4766
rect -39 4668 -22 4714
rect 24 4668 41 4714
rect -39 4616 41 4668
rect -39 4570 -22 4616
rect 24 4570 41 4616
rect -39 4518 41 4570
rect -39 4472 -22 4518
rect 24 4472 41 4518
rect -39 4420 41 4472
rect -39 4374 -22 4420
rect 24 4374 41 4420
rect -39 4322 41 4374
rect -39 4276 -22 4322
rect 24 4276 41 4322
rect -39 4224 41 4276
rect -39 4178 -22 4224
rect 24 4178 41 4224
rect -39 4126 41 4178
rect -39 4080 -22 4126
rect 24 4080 41 4126
rect -39 4028 41 4080
rect -39 3982 -22 4028
rect 24 3982 41 4028
rect -39 3930 41 3982
rect -39 3884 -22 3930
rect 24 3884 41 3930
rect -39 3832 41 3884
rect -39 3786 -22 3832
rect 24 3786 41 3832
rect -39 3734 41 3786
rect -39 3688 -22 3734
rect 24 3688 41 3734
rect -39 3636 41 3688
rect -39 3590 -22 3636
rect 24 3590 41 3636
rect -39 3538 41 3590
rect 135 5507 9895 5579
rect 135 4927 207 5507
rect 9823 4927 9895 5507
rect 135 4855 9895 4927
rect 135 4275 207 4855
rect 9823 4275 9895 4855
rect 135 4203 9895 4275
rect 135 3623 207 4203
rect 9823 3623 9895 4203
rect 135 3551 9895 3623
rect 9989 5550 10006 5596
rect 10052 5550 10069 5596
rect 9989 5498 10069 5550
rect 9989 5452 10006 5498
rect 10052 5452 10069 5498
rect 9989 5400 10069 5452
rect 9989 5354 10006 5400
rect 10052 5354 10069 5400
rect 9989 5302 10069 5354
rect 9989 5256 10006 5302
rect 10052 5256 10069 5302
rect 9989 5204 10069 5256
rect 9989 5158 10006 5204
rect 10052 5158 10069 5204
rect 9989 5106 10069 5158
rect 9989 5060 10006 5106
rect 10052 5060 10069 5106
rect 9989 5008 10069 5060
rect 9989 4962 10006 5008
rect 10052 4962 10069 5008
rect 9989 4910 10069 4962
rect 9989 4864 10006 4910
rect 10052 4864 10069 4910
rect 9989 4812 10069 4864
rect 9989 4766 10006 4812
rect 10052 4766 10069 4812
rect 9989 4714 10069 4766
rect 9989 4668 10006 4714
rect 10052 4668 10069 4714
rect 9989 4616 10069 4668
rect 9989 4570 10006 4616
rect 10052 4570 10069 4616
rect 9989 4518 10069 4570
rect 9989 4472 10006 4518
rect 10052 4472 10069 4518
rect 9989 4420 10069 4472
rect 9989 4374 10006 4420
rect 10052 4374 10069 4420
rect 9989 4322 10069 4374
rect 9989 4276 10006 4322
rect 10052 4276 10069 4322
rect 9989 4224 10069 4276
rect 9989 4178 10006 4224
rect 10052 4178 10069 4224
rect 9989 4126 10069 4178
rect 9989 4080 10006 4126
rect 10052 4080 10069 4126
rect 9989 4028 10069 4080
rect 9989 3982 10006 4028
rect 10052 3982 10069 4028
rect 9989 3930 10069 3982
rect 9989 3884 10006 3930
rect 10052 3884 10069 3930
rect 9989 3832 10069 3884
rect 9989 3786 10006 3832
rect 10052 3786 10069 3832
rect 9989 3734 10069 3786
rect 9989 3688 10006 3734
rect 10052 3688 10069 3734
rect 9989 3636 10069 3688
rect 9989 3590 10006 3636
rect 10052 3590 10069 3636
rect -39 3492 -22 3538
rect 24 3492 41 3538
rect -39 3457 41 3492
rect 9989 3538 10069 3590
rect 9989 3492 10006 3538
rect 10052 3492 10069 3538
rect 9989 3457 10069 3492
rect -39 3440 10069 3457
rect -39 3394 -22 3440
rect 24 3394 76 3440
rect 122 3394 174 3440
rect 220 3394 272 3440
rect 318 3394 370 3440
rect 416 3394 468 3440
rect 514 3394 566 3440
rect 612 3394 664 3440
rect 710 3394 762 3440
rect 808 3394 860 3440
rect 906 3394 958 3440
rect 1004 3394 1056 3440
rect 1102 3394 1154 3440
rect 1200 3394 1252 3440
rect 1298 3394 1350 3440
rect 1396 3394 1448 3440
rect 1494 3394 1546 3440
rect 1592 3394 1644 3440
rect 1690 3394 1742 3440
rect 1788 3394 1840 3440
rect 1886 3394 1938 3440
rect 1984 3394 2036 3440
rect 2082 3394 2134 3440
rect 2180 3394 2232 3440
rect 2278 3394 2330 3440
rect 2376 3394 2428 3440
rect 2474 3394 2526 3440
rect 2572 3394 2624 3440
rect 2670 3394 2722 3440
rect 2768 3394 2820 3440
rect 2866 3394 2918 3440
rect 2964 3394 3016 3440
rect 3062 3394 3114 3440
rect 3160 3394 3212 3440
rect 3258 3394 3310 3440
rect 3356 3394 3408 3440
rect 3454 3394 3506 3440
rect 3552 3394 3604 3440
rect 3650 3394 3702 3440
rect 3748 3394 3800 3440
rect 3846 3394 3898 3440
rect 3944 3394 3996 3440
rect 4042 3394 4094 3440
rect 4140 3394 4192 3440
rect 4238 3394 4290 3440
rect 4336 3394 4388 3440
rect 4434 3394 4486 3440
rect 4532 3394 4584 3440
rect 4630 3394 4682 3440
rect 4728 3394 4780 3440
rect 4826 3394 4878 3440
rect 4924 3394 4976 3440
rect 5022 3394 5074 3440
rect 5120 3394 5172 3440
rect 5218 3394 5270 3440
rect 5316 3394 5368 3440
rect 5414 3394 5466 3440
rect 5512 3394 5564 3440
rect 5610 3394 5662 3440
rect 5708 3394 5760 3440
rect 5806 3394 5858 3440
rect 5904 3394 5956 3440
rect 6002 3394 6054 3440
rect 6100 3394 6152 3440
rect 6198 3394 6250 3440
rect 6296 3394 6348 3440
rect 6394 3394 6446 3440
rect 6492 3394 6544 3440
rect 6590 3394 6642 3440
rect 6688 3394 6740 3440
rect 6786 3394 6838 3440
rect 6884 3394 6936 3440
rect 6982 3394 7034 3440
rect 7080 3394 7132 3440
rect 7178 3394 7230 3440
rect 7276 3394 7328 3440
rect 7374 3394 7426 3440
rect 7472 3394 7524 3440
rect 7570 3394 7622 3440
rect 7668 3394 7720 3440
rect 7766 3394 7818 3440
rect 7864 3394 7916 3440
rect 7962 3394 8014 3440
rect 8060 3394 8112 3440
rect 8158 3394 8210 3440
rect 8256 3394 8308 3440
rect 8354 3394 8406 3440
rect 8452 3394 8504 3440
rect 8550 3394 8602 3440
rect 8648 3394 8700 3440
rect 8746 3394 8798 3440
rect 8844 3394 8896 3440
rect 8942 3394 8994 3440
rect 9040 3394 9092 3440
rect 9138 3394 9190 3440
rect 9236 3394 9288 3440
rect 9334 3394 9386 3440
rect 9432 3394 9484 3440
rect 9530 3394 9582 3440
rect 9628 3394 9680 3440
rect 9726 3394 9778 3440
rect 9824 3394 9876 3440
rect 9922 3394 10006 3440
rect 10052 3394 10069 3440
rect -39 3377 10069 3394
rect -39 3269 10069 3286
rect -39 3219 -22 3269
rect 24 3223 76 3269
rect 122 3223 174 3269
rect 220 3223 272 3269
rect 318 3223 370 3269
rect 416 3223 468 3269
rect 514 3223 566 3269
rect 612 3223 664 3269
rect 710 3223 762 3269
rect 808 3223 860 3269
rect 906 3223 958 3269
rect 1004 3223 1056 3269
rect 1102 3223 1154 3269
rect 1200 3223 1252 3269
rect 1298 3223 1350 3269
rect 1396 3223 1448 3269
rect 1494 3223 1546 3269
rect 1592 3223 1644 3269
rect 1690 3223 1742 3269
rect 1788 3223 1840 3269
rect 1886 3223 1938 3269
rect 1984 3223 2036 3269
rect 2082 3223 2134 3269
rect 2180 3223 2232 3269
rect 2278 3223 2330 3269
rect 2376 3223 2428 3269
rect 2474 3223 2526 3269
rect 2572 3223 2624 3269
rect 2670 3223 2722 3269
rect 2768 3223 2820 3269
rect 2866 3223 2918 3269
rect 2964 3223 3016 3269
rect 3062 3223 3114 3269
rect 3160 3223 3212 3269
rect 3258 3223 3310 3269
rect 3356 3223 3408 3269
rect 3454 3223 3506 3269
rect 3552 3223 3604 3269
rect 3650 3223 3702 3269
rect 3748 3223 3800 3269
rect 3846 3223 3898 3269
rect 3944 3223 3996 3269
rect 4042 3223 4094 3269
rect 4140 3223 4192 3269
rect 4238 3223 4290 3269
rect 4336 3223 4388 3269
rect 4434 3223 4486 3269
rect 4532 3223 4584 3269
rect 4630 3223 4682 3269
rect 4728 3223 4780 3269
rect 4826 3223 4878 3269
rect 4924 3223 4976 3269
rect 5022 3223 5074 3269
rect 5120 3223 5172 3269
rect 5218 3223 5270 3269
rect 5316 3223 5368 3269
rect 5414 3223 5466 3269
rect 5512 3223 5564 3269
rect 5610 3223 5662 3269
rect 5708 3223 5760 3269
rect 5806 3223 5858 3269
rect 5904 3223 5956 3269
rect 6002 3223 6054 3269
rect 6100 3223 6152 3269
rect 6198 3223 6250 3269
rect 6296 3223 6348 3269
rect 6394 3223 6446 3269
rect 6492 3223 6544 3269
rect 6590 3223 6642 3269
rect 6688 3223 6740 3269
rect 6786 3223 6838 3269
rect 6884 3223 6936 3269
rect 6982 3223 7034 3269
rect 7080 3223 7132 3269
rect 7178 3223 7230 3269
rect 7276 3223 7328 3269
rect 7374 3223 7426 3269
rect 7472 3223 7524 3269
rect 7570 3223 7622 3269
rect 7668 3223 7720 3269
rect 7766 3223 7818 3269
rect 7864 3223 7916 3269
rect 7962 3223 8014 3269
rect 8060 3223 8112 3269
rect 8158 3223 8210 3269
rect 8256 3223 8308 3269
rect 8354 3223 8406 3269
rect 8452 3223 8504 3269
rect 8550 3223 8602 3269
rect 8648 3223 8700 3269
rect 8746 3223 8798 3269
rect 8844 3223 8896 3269
rect 8942 3223 8994 3269
rect 9040 3223 9092 3269
rect 9138 3223 9190 3269
rect 9236 3223 9288 3269
rect 9334 3223 9386 3269
rect 9432 3223 9484 3269
rect 9530 3223 9582 3269
rect 9628 3223 9680 3269
rect 9726 3223 9778 3269
rect 9824 3223 9876 3269
rect 9922 3223 10006 3269
rect 24 3219 10006 3223
rect 10052 3219 10069 3269
rect -39 3206 10069 3219
rect -39 3167 41 3206
rect -39 3121 -22 3167
rect 24 3121 41 3167
rect 9989 3167 10069 3206
rect -39 3069 41 3121
rect -39 3023 -22 3069
rect 24 3023 41 3069
rect -39 2971 41 3023
rect -39 2925 -22 2971
rect 24 2925 41 2971
rect -39 2873 41 2925
rect -39 2827 -22 2873
rect 24 2827 41 2873
rect -39 2775 41 2827
rect -39 2729 -22 2775
rect 24 2729 41 2775
rect -39 2677 41 2729
rect -39 2631 -22 2677
rect 24 2631 41 2677
rect -39 2579 41 2631
rect -39 2533 -22 2579
rect 24 2533 41 2579
rect -39 2481 41 2533
rect -39 2435 -22 2481
rect 24 2435 41 2481
rect -39 2383 41 2435
rect -39 2337 -22 2383
rect 24 2337 41 2383
rect -39 2285 41 2337
rect -39 2239 -22 2285
rect 24 2239 41 2285
rect -39 2187 41 2239
rect -39 2141 -22 2187
rect 24 2141 41 2187
rect -39 2089 41 2141
rect -39 2043 -22 2089
rect 24 2043 41 2089
rect -39 1991 41 2043
rect -39 1945 -22 1991
rect 24 1945 41 1991
rect -39 1893 41 1945
rect -39 1847 -22 1893
rect 24 1847 41 1893
rect -39 1795 41 1847
rect -39 1749 -22 1795
rect 24 1749 41 1795
rect -39 1697 41 1749
rect -39 1651 -22 1697
rect 24 1651 41 1697
rect -39 1599 41 1651
rect -39 1553 -22 1599
rect 24 1553 41 1599
rect -39 1501 41 1553
rect -39 1455 -22 1501
rect 24 1455 41 1501
rect -39 1403 41 1455
rect -39 1357 -22 1403
rect 24 1357 41 1403
rect -39 1305 41 1357
rect -39 1259 -22 1305
rect 24 1259 41 1305
rect -39 1207 41 1259
rect -39 1161 -22 1207
rect 24 1161 41 1207
rect -39 1109 41 1161
rect 135 3078 9895 3150
rect 135 2498 207 3078
rect 9823 2498 9895 3078
rect 135 2426 9895 2498
rect 135 1846 207 2426
rect 9823 1846 9895 2426
rect 135 1774 9895 1846
rect 135 1194 207 1774
rect 9823 1194 9895 1774
rect 135 1122 9895 1194
rect 9989 3121 10006 3167
rect 10052 3121 10069 3167
rect 9989 3069 10069 3121
rect 9989 3023 10006 3069
rect 10052 3023 10069 3069
rect 9989 2971 10069 3023
rect 9989 2925 10006 2971
rect 10052 2925 10069 2971
rect 9989 2873 10069 2925
rect 9989 2827 10006 2873
rect 10052 2827 10069 2873
rect 9989 2775 10069 2827
rect 9989 2729 10006 2775
rect 10052 2729 10069 2775
rect 9989 2677 10069 2729
rect 9989 2631 10006 2677
rect 10052 2631 10069 2677
rect 9989 2579 10069 2631
rect 9989 2533 10006 2579
rect 10052 2533 10069 2579
rect 9989 2481 10069 2533
rect 9989 2435 10006 2481
rect 10052 2435 10069 2481
rect 9989 2383 10069 2435
rect 9989 2337 10006 2383
rect 10052 2337 10069 2383
rect 9989 2285 10069 2337
rect 9989 2239 10006 2285
rect 10052 2239 10069 2285
rect 9989 2187 10069 2239
rect 9989 2141 10006 2187
rect 10052 2141 10069 2187
rect 9989 2089 10069 2141
rect 9989 2043 10006 2089
rect 10052 2043 10069 2089
rect 9989 1991 10069 2043
rect 9989 1945 10006 1991
rect 10052 1945 10069 1991
rect 9989 1893 10069 1945
rect 9989 1847 10006 1893
rect 10052 1847 10069 1893
rect 9989 1795 10069 1847
rect 9989 1749 10006 1795
rect 10052 1749 10069 1795
rect 9989 1697 10069 1749
rect 9989 1651 10006 1697
rect 10052 1651 10069 1697
rect 9989 1599 10069 1651
rect 9989 1553 10006 1599
rect 10052 1553 10069 1599
rect 9989 1501 10069 1553
rect 9989 1455 10006 1501
rect 10052 1455 10069 1501
rect 9989 1403 10069 1455
rect 9989 1357 10006 1403
rect 10052 1357 10069 1403
rect 9989 1305 10069 1357
rect 9989 1259 10006 1305
rect 10052 1259 10069 1305
rect 9989 1207 10069 1259
rect 9989 1161 10006 1207
rect 10052 1161 10069 1207
rect -39 1063 -22 1109
rect 24 1063 41 1109
rect -39 1028 41 1063
rect 9989 1109 10069 1161
rect 9989 1063 10006 1109
rect 10052 1063 10069 1109
rect 9989 1028 10069 1063
rect -39 1011 10069 1028
rect -39 965 -22 1011
rect 24 965 76 1011
rect 122 965 174 1011
rect 220 965 272 1011
rect 318 965 370 1011
rect 416 965 468 1011
rect 514 965 566 1011
rect 612 965 664 1011
rect 710 965 762 1011
rect 808 965 860 1011
rect 906 965 958 1011
rect 1004 965 1056 1011
rect 1102 965 1154 1011
rect 1200 965 1252 1011
rect 1298 965 1350 1011
rect 1396 965 1448 1011
rect 1494 965 1546 1011
rect 1592 965 1644 1011
rect 1690 965 1742 1011
rect 1788 965 1840 1011
rect 1886 965 1938 1011
rect 1984 965 2036 1011
rect 2082 965 2134 1011
rect 2180 965 2232 1011
rect 2278 965 2330 1011
rect 2376 965 2428 1011
rect 2474 965 2526 1011
rect 2572 965 2624 1011
rect 2670 965 2722 1011
rect 2768 965 2820 1011
rect 2866 965 2918 1011
rect 2964 965 3016 1011
rect 3062 965 3114 1011
rect 3160 965 3212 1011
rect 3258 965 3310 1011
rect 3356 965 3408 1011
rect 3454 965 3506 1011
rect 3552 965 3604 1011
rect 3650 965 3702 1011
rect 3748 965 3800 1011
rect 3846 965 3898 1011
rect 3944 965 3996 1011
rect 4042 965 4094 1011
rect 4140 965 4192 1011
rect 4238 965 4290 1011
rect 4336 965 4388 1011
rect 4434 965 4486 1011
rect 4532 965 4584 1011
rect 4630 965 4682 1011
rect 4728 965 4780 1011
rect 4826 965 4878 1011
rect 4924 965 4976 1011
rect 5022 965 5074 1011
rect 5120 965 5172 1011
rect 5218 965 5270 1011
rect 5316 965 5368 1011
rect 5414 965 5466 1011
rect 5512 965 5564 1011
rect 5610 965 5662 1011
rect 5708 965 5760 1011
rect 5806 965 5858 1011
rect 5904 965 5956 1011
rect 6002 965 6054 1011
rect 6100 965 6152 1011
rect 6198 965 6250 1011
rect 6296 965 6348 1011
rect 6394 965 6446 1011
rect 6492 965 6544 1011
rect 6590 965 6642 1011
rect 6688 965 6740 1011
rect 6786 965 6838 1011
rect 6884 965 6936 1011
rect 6982 965 7034 1011
rect 7080 965 7132 1011
rect 7178 965 7230 1011
rect 7276 965 7328 1011
rect 7374 965 7426 1011
rect 7472 965 7524 1011
rect 7570 965 7622 1011
rect 7668 965 7720 1011
rect 7766 965 7818 1011
rect 7864 965 7916 1011
rect 7962 965 8014 1011
rect 8060 965 8112 1011
rect 8158 965 8210 1011
rect 8256 965 8308 1011
rect 8354 965 8406 1011
rect 8452 965 8504 1011
rect 8550 965 8602 1011
rect 8648 965 8700 1011
rect 8746 965 8798 1011
rect 8844 965 8896 1011
rect 8942 965 8994 1011
rect 9040 965 9092 1011
rect 9138 965 9190 1011
rect 9236 965 9288 1011
rect 9334 965 9386 1011
rect 9432 965 9484 1011
rect 9530 965 9582 1011
rect 9628 965 9680 1011
rect 9726 965 9778 1011
rect 9824 965 9876 1011
rect 9922 965 10006 1011
rect 10052 965 10069 1011
rect -39 948 10069 965
<< nsubdiffcont >>
rect -22 5648 24 5698
rect 76 5652 122 5698
rect 174 5652 220 5698
rect 272 5652 318 5698
rect 370 5652 416 5698
rect 468 5652 514 5698
rect 566 5652 612 5698
rect 664 5652 710 5698
rect 762 5652 808 5698
rect 860 5652 906 5698
rect 958 5652 1004 5698
rect 1056 5652 1102 5698
rect 1154 5652 1200 5698
rect 1252 5652 1298 5698
rect 1350 5652 1396 5698
rect 1448 5652 1494 5698
rect 1546 5652 1592 5698
rect 1644 5652 1690 5698
rect 1742 5652 1788 5698
rect 1840 5652 1886 5698
rect 1938 5652 1984 5698
rect 2036 5652 2082 5698
rect 2134 5652 2180 5698
rect 2232 5652 2278 5698
rect 2330 5652 2376 5698
rect 2428 5652 2474 5698
rect 2526 5652 2572 5698
rect 2624 5652 2670 5698
rect 2722 5652 2768 5698
rect 2820 5652 2866 5698
rect 2918 5652 2964 5698
rect 3016 5652 3062 5698
rect 3114 5652 3160 5698
rect 3212 5652 3258 5698
rect 3310 5652 3356 5698
rect 3408 5652 3454 5698
rect 3506 5652 3552 5698
rect 3604 5652 3650 5698
rect 3702 5652 3748 5698
rect 3800 5652 3846 5698
rect 3898 5652 3944 5698
rect 3996 5652 4042 5698
rect 4094 5652 4140 5698
rect 4192 5652 4238 5698
rect 4290 5652 4336 5698
rect 4388 5652 4434 5698
rect 4486 5652 4532 5698
rect 4584 5652 4630 5698
rect 4682 5652 4728 5698
rect 4780 5652 4826 5698
rect 4878 5652 4924 5698
rect 4976 5652 5022 5698
rect 5074 5652 5120 5698
rect 5172 5652 5218 5698
rect 5270 5652 5316 5698
rect 5368 5652 5414 5698
rect 5466 5652 5512 5698
rect 5564 5652 5610 5698
rect 5662 5652 5708 5698
rect 5760 5652 5806 5698
rect 5858 5652 5904 5698
rect 5956 5652 6002 5698
rect 6054 5652 6100 5698
rect 6152 5652 6198 5698
rect 6250 5652 6296 5698
rect 6348 5652 6394 5698
rect 6446 5652 6492 5698
rect 6544 5652 6590 5698
rect 6642 5652 6688 5698
rect 6740 5652 6786 5698
rect 6838 5652 6884 5698
rect 6936 5652 6982 5698
rect 7034 5652 7080 5698
rect 7132 5652 7178 5698
rect 7230 5652 7276 5698
rect 7328 5652 7374 5698
rect 7426 5652 7472 5698
rect 7524 5652 7570 5698
rect 7622 5652 7668 5698
rect 7720 5652 7766 5698
rect 7818 5652 7864 5698
rect 7916 5652 7962 5698
rect 8014 5652 8060 5698
rect 8112 5652 8158 5698
rect 8210 5652 8256 5698
rect 8308 5652 8354 5698
rect 8406 5652 8452 5698
rect 8504 5652 8550 5698
rect 8602 5652 8648 5698
rect 8700 5652 8746 5698
rect 8798 5652 8844 5698
rect 8896 5652 8942 5698
rect 8994 5652 9040 5698
rect 9092 5652 9138 5698
rect 9190 5652 9236 5698
rect 9288 5652 9334 5698
rect 9386 5652 9432 5698
rect 9484 5652 9530 5698
rect 9582 5652 9628 5698
rect 9680 5652 9726 5698
rect 9778 5652 9824 5698
rect 9876 5652 9922 5698
rect 10006 5648 10052 5698
rect -22 5550 24 5596
rect -22 5452 24 5498
rect -22 5354 24 5400
rect -22 5256 24 5302
rect -22 5158 24 5204
rect -22 5060 24 5106
rect -22 4962 24 5008
rect -22 4864 24 4910
rect -22 4766 24 4812
rect -22 4668 24 4714
rect -22 4570 24 4616
rect -22 4472 24 4518
rect -22 4374 24 4420
rect -22 4276 24 4322
rect -22 4178 24 4224
rect -22 4080 24 4126
rect -22 3982 24 4028
rect -22 3884 24 3930
rect -22 3786 24 3832
rect -22 3688 24 3734
rect -22 3590 24 3636
rect 10006 5550 10052 5596
rect 10006 5452 10052 5498
rect 10006 5354 10052 5400
rect 10006 5256 10052 5302
rect 10006 5158 10052 5204
rect 10006 5060 10052 5106
rect 10006 4962 10052 5008
rect 10006 4864 10052 4910
rect 10006 4766 10052 4812
rect 10006 4668 10052 4714
rect 10006 4570 10052 4616
rect 10006 4472 10052 4518
rect 10006 4374 10052 4420
rect 10006 4276 10052 4322
rect 10006 4178 10052 4224
rect 10006 4080 10052 4126
rect 10006 3982 10052 4028
rect 10006 3884 10052 3930
rect 10006 3786 10052 3832
rect 10006 3688 10052 3734
rect 10006 3590 10052 3636
rect -22 3492 24 3538
rect 10006 3492 10052 3538
rect -22 3394 24 3440
rect 76 3394 122 3440
rect 174 3394 220 3440
rect 272 3394 318 3440
rect 370 3394 416 3440
rect 468 3394 514 3440
rect 566 3394 612 3440
rect 664 3394 710 3440
rect 762 3394 808 3440
rect 860 3394 906 3440
rect 958 3394 1004 3440
rect 1056 3394 1102 3440
rect 1154 3394 1200 3440
rect 1252 3394 1298 3440
rect 1350 3394 1396 3440
rect 1448 3394 1494 3440
rect 1546 3394 1592 3440
rect 1644 3394 1690 3440
rect 1742 3394 1788 3440
rect 1840 3394 1886 3440
rect 1938 3394 1984 3440
rect 2036 3394 2082 3440
rect 2134 3394 2180 3440
rect 2232 3394 2278 3440
rect 2330 3394 2376 3440
rect 2428 3394 2474 3440
rect 2526 3394 2572 3440
rect 2624 3394 2670 3440
rect 2722 3394 2768 3440
rect 2820 3394 2866 3440
rect 2918 3394 2964 3440
rect 3016 3394 3062 3440
rect 3114 3394 3160 3440
rect 3212 3394 3258 3440
rect 3310 3394 3356 3440
rect 3408 3394 3454 3440
rect 3506 3394 3552 3440
rect 3604 3394 3650 3440
rect 3702 3394 3748 3440
rect 3800 3394 3846 3440
rect 3898 3394 3944 3440
rect 3996 3394 4042 3440
rect 4094 3394 4140 3440
rect 4192 3394 4238 3440
rect 4290 3394 4336 3440
rect 4388 3394 4434 3440
rect 4486 3394 4532 3440
rect 4584 3394 4630 3440
rect 4682 3394 4728 3440
rect 4780 3394 4826 3440
rect 4878 3394 4924 3440
rect 4976 3394 5022 3440
rect 5074 3394 5120 3440
rect 5172 3394 5218 3440
rect 5270 3394 5316 3440
rect 5368 3394 5414 3440
rect 5466 3394 5512 3440
rect 5564 3394 5610 3440
rect 5662 3394 5708 3440
rect 5760 3394 5806 3440
rect 5858 3394 5904 3440
rect 5956 3394 6002 3440
rect 6054 3394 6100 3440
rect 6152 3394 6198 3440
rect 6250 3394 6296 3440
rect 6348 3394 6394 3440
rect 6446 3394 6492 3440
rect 6544 3394 6590 3440
rect 6642 3394 6688 3440
rect 6740 3394 6786 3440
rect 6838 3394 6884 3440
rect 6936 3394 6982 3440
rect 7034 3394 7080 3440
rect 7132 3394 7178 3440
rect 7230 3394 7276 3440
rect 7328 3394 7374 3440
rect 7426 3394 7472 3440
rect 7524 3394 7570 3440
rect 7622 3394 7668 3440
rect 7720 3394 7766 3440
rect 7818 3394 7864 3440
rect 7916 3394 7962 3440
rect 8014 3394 8060 3440
rect 8112 3394 8158 3440
rect 8210 3394 8256 3440
rect 8308 3394 8354 3440
rect 8406 3394 8452 3440
rect 8504 3394 8550 3440
rect 8602 3394 8648 3440
rect 8700 3394 8746 3440
rect 8798 3394 8844 3440
rect 8896 3394 8942 3440
rect 8994 3394 9040 3440
rect 9092 3394 9138 3440
rect 9190 3394 9236 3440
rect 9288 3394 9334 3440
rect 9386 3394 9432 3440
rect 9484 3394 9530 3440
rect 9582 3394 9628 3440
rect 9680 3394 9726 3440
rect 9778 3394 9824 3440
rect 9876 3394 9922 3440
rect 10006 3394 10052 3440
rect -22 3219 24 3269
rect 76 3223 122 3269
rect 174 3223 220 3269
rect 272 3223 318 3269
rect 370 3223 416 3269
rect 468 3223 514 3269
rect 566 3223 612 3269
rect 664 3223 710 3269
rect 762 3223 808 3269
rect 860 3223 906 3269
rect 958 3223 1004 3269
rect 1056 3223 1102 3269
rect 1154 3223 1200 3269
rect 1252 3223 1298 3269
rect 1350 3223 1396 3269
rect 1448 3223 1494 3269
rect 1546 3223 1592 3269
rect 1644 3223 1690 3269
rect 1742 3223 1788 3269
rect 1840 3223 1886 3269
rect 1938 3223 1984 3269
rect 2036 3223 2082 3269
rect 2134 3223 2180 3269
rect 2232 3223 2278 3269
rect 2330 3223 2376 3269
rect 2428 3223 2474 3269
rect 2526 3223 2572 3269
rect 2624 3223 2670 3269
rect 2722 3223 2768 3269
rect 2820 3223 2866 3269
rect 2918 3223 2964 3269
rect 3016 3223 3062 3269
rect 3114 3223 3160 3269
rect 3212 3223 3258 3269
rect 3310 3223 3356 3269
rect 3408 3223 3454 3269
rect 3506 3223 3552 3269
rect 3604 3223 3650 3269
rect 3702 3223 3748 3269
rect 3800 3223 3846 3269
rect 3898 3223 3944 3269
rect 3996 3223 4042 3269
rect 4094 3223 4140 3269
rect 4192 3223 4238 3269
rect 4290 3223 4336 3269
rect 4388 3223 4434 3269
rect 4486 3223 4532 3269
rect 4584 3223 4630 3269
rect 4682 3223 4728 3269
rect 4780 3223 4826 3269
rect 4878 3223 4924 3269
rect 4976 3223 5022 3269
rect 5074 3223 5120 3269
rect 5172 3223 5218 3269
rect 5270 3223 5316 3269
rect 5368 3223 5414 3269
rect 5466 3223 5512 3269
rect 5564 3223 5610 3269
rect 5662 3223 5708 3269
rect 5760 3223 5806 3269
rect 5858 3223 5904 3269
rect 5956 3223 6002 3269
rect 6054 3223 6100 3269
rect 6152 3223 6198 3269
rect 6250 3223 6296 3269
rect 6348 3223 6394 3269
rect 6446 3223 6492 3269
rect 6544 3223 6590 3269
rect 6642 3223 6688 3269
rect 6740 3223 6786 3269
rect 6838 3223 6884 3269
rect 6936 3223 6982 3269
rect 7034 3223 7080 3269
rect 7132 3223 7178 3269
rect 7230 3223 7276 3269
rect 7328 3223 7374 3269
rect 7426 3223 7472 3269
rect 7524 3223 7570 3269
rect 7622 3223 7668 3269
rect 7720 3223 7766 3269
rect 7818 3223 7864 3269
rect 7916 3223 7962 3269
rect 8014 3223 8060 3269
rect 8112 3223 8158 3269
rect 8210 3223 8256 3269
rect 8308 3223 8354 3269
rect 8406 3223 8452 3269
rect 8504 3223 8550 3269
rect 8602 3223 8648 3269
rect 8700 3223 8746 3269
rect 8798 3223 8844 3269
rect 8896 3223 8942 3269
rect 8994 3223 9040 3269
rect 9092 3223 9138 3269
rect 9190 3223 9236 3269
rect 9288 3223 9334 3269
rect 9386 3223 9432 3269
rect 9484 3223 9530 3269
rect 9582 3223 9628 3269
rect 9680 3223 9726 3269
rect 9778 3223 9824 3269
rect 9876 3223 9922 3269
rect 10006 3219 10052 3269
rect -22 3121 24 3167
rect -22 3023 24 3069
rect -22 2925 24 2971
rect -22 2827 24 2873
rect -22 2729 24 2775
rect -22 2631 24 2677
rect -22 2533 24 2579
rect -22 2435 24 2481
rect -22 2337 24 2383
rect -22 2239 24 2285
rect -22 2141 24 2187
rect -22 2043 24 2089
rect -22 1945 24 1991
rect -22 1847 24 1893
rect -22 1749 24 1795
rect -22 1651 24 1697
rect -22 1553 24 1599
rect -22 1455 24 1501
rect -22 1357 24 1403
rect -22 1259 24 1305
rect -22 1161 24 1207
rect 10006 3121 10052 3167
rect 10006 3023 10052 3069
rect 10006 2925 10052 2971
rect 10006 2827 10052 2873
rect 10006 2729 10052 2775
rect 10006 2631 10052 2677
rect 10006 2533 10052 2579
rect 10006 2435 10052 2481
rect 10006 2337 10052 2383
rect 10006 2239 10052 2285
rect 10006 2141 10052 2187
rect 10006 2043 10052 2089
rect 10006 1945 10052 1991
rect 10006 1847 10052 1893
rect 10006 1749 10052 1795
rect 10006 1651 10052 1697
rect 10006 1553 10052 1599
rect 10006 1455 10052 1501
rect 10006 1357 10052 1403
rect 10006 1259 10052 1305
rect 10006 1161 10052 1207
rect -22 1063 24 1109
rect 10006 1063 10052 1109
rect -22 965 24 1011
rect 76 965 122 1011
rect 174 965 220 1011
rect 272 965 318 1011
rect 370 965 416 1011
rect 468 965 514 1011
rect 566 965 612 1011
rect 664 965 710 1011
rect 762 965 808 1011
rect 860 965 906 1011
rect 958 965 1004 1011
rect 1056 965 1102 1011
rect 1154 965 1200 1011
rect 1252 965 1298 1011
rect 1350 965 1396 1011
rect 1448 965 1494 1011
rect 1546 965 1592 1011
rect 1644 965 1690 1011
rect 1742 965 1788 1011
rect 1840 965 1886 1011
rect 1938 965 1984 1011
rect 2036 965 2082 1011
rect 2134 965 2180 1011
rect 2232 965 2278 1011
rect 2330 965 2376 1011
rect 2428 965 2474 1011
rect 2526 965 2572 1011
rect 2624 965 2670 1011
rect 2722 965 2768 1011
rect 2820 965 2866 1011
rect 2918 965 2964 1011
rect 3016 965 3062 1011
rect 3114 965 3160 1011
rect 3212 965 3258 1011
rect 3310 965 3356 1011
rect 3408 965 3454 1011
rect 3506 965 3552 1011
rect 3604 965 3650 1011
rect 3702 965 3748 1011
rect 3800 965 3846 1011
rect 3898 965 3944 1011
rect 3996 965 4042 1011
rect 4094 965 4140 1011
rect 4192 965 4238 1011
rect 4290 965 4336 1011
rect 4388 965 4434 1011
rect 4486 965 4532 1011
rect 4584 965 4630 1011
rect 4682 965 4728 1011
rect 4780 965 4826 1011
rect 4878 965 4924 1011
rect 4976 965 5022 1011
rect 5074 965 5120 1011
rect 5172 965 5218 1011
rect 5270 965 5316 1011
rect 5368 965 5414 1011
rect 5466 965 5512 1011
rect 5564 965 5610 1011
rect 5662 965 5708 1011
rect 5760 965 5806 1011
rect 5858 965 5904 1011
rect 5956 965 6002 1011
rect 6054 965 6100 1011
rect 6152 965 6198 1011
rect 6250 965 6296 1011
rect 6348 965 6394 1011
rect 6446 965 6492 1011
rect 6544 965 6590 1011
rect 6642 965 6688 1011
rect 6740 965 6786 1011
rect 6838 965 6884 1011
rect 6936 965 6982 1011
rect 7034 965 7080 1011
rect 7132 965 7178 1011
rect 7230 965 7276 1011
rect 7328 965 7374 1011
rect 7426 965 7472 1011
rect 7524 965 7570 1011
rect 7622 965 7668 1011
rect 7720 965 7766 1011
rect 7818 965 7864 1011
rect 7916 965 7962 1011
rect 8014 965 8060 1011
rect 8112 965 8158 1011
rect 8210 965 8256 1011
rect 8308 965 8354 1011
rect 8406 965 8452 1011
rect 8504 965 8550 1011
rect 8602 965 8648 1011
rect 8700 965 8746 1011
rect 8798 965 8844 1011
rect 8896 965 8942 1011
rect 8994 965 9040 1011
rect 9092 965 9138 1011
rect 9190 965 9236 1011
rect 9288 965 9334 1011
rect 9386 965 9432 1011
rect 9484 965 9530 1011
rect 9582 965 9628 1011
rect 9680 965 9726 1011
rect 9778 965 9824 1011
rect 9876 965 9922 1011
rect 10006 965 10052 1011
<< polysilicon >>
rect 295 5406 495 5419
rect 295 5360 308 5406
rect 482 5360 495 5406
rect 295 5317 495 5360
rect 295 5074 495 5117
rect 295 5028 308 5074
rect 482 5028 495 5074
rect 295 5015 495 5028
rect 575 5406 775 5419
rect 575 5360 588 5406
rect 762 5360 775 5406
rect 575 5317 775 5360
rect 575 5074 775 5117
rect 575 5028 588 5074
rect 762 5028 775 5074
rect 575 5015 775 5028
rect 855 5406 1055 5419
rect 855 5360 868 5406
rect 1042 5360 1055 5406
rect 855 5317 1055 5360
rect 855 5074 1055 5117
rect 855 5028 868 5074
rect 1042 5028 1055 5074
rect 855 5015 1055 5028
rect 1135 5406 1335 5419
rect 1135 5360 1148 5406
rect 1322 5360 1335 5406
rect 1135 5317 1335 5360
rect 1135 5074 1335 5117
rect 1135 5028 1148 5074
rect 1322 5028 1335 5074
rect 1135 5015 1335 5028
rect 1415 5406 1615 5419
rect 1415 5360 1428 5406
rect 1602 5360 1615 5406
rect 1415 5317 1615 5360
rect 1415 5074 1615 5117
rect 1415 5028 1428 5074
rect 1602 5028 1615 5074
rect 1415 5015 1615 5028
rect 1695 5406 1895 5419
rect 1695 5360 1708 5406
rect 1882 5360 1895 5406
rect 1695 5317 1895 5360
rect 1695 5074 1895 5117
rect 1695 5028 1708 5074
rect 1882 5028 1895 5074
rect 1695 5015 1895 5028
rect 1975 5406 2175 5419
rect 1975 5360 1988 5406
rect 2162 5360 2175 5406
rect 1975 5317 2175 5360
rect 1975 5074 2175 5117
rect 1975 5028 1988 5074
rect 2162 5028 2175 5074
rect 1975 5015 2175 5028
rect 2255 5406 2455 5419
rect 2255 5360 2268 5406
rect 2442 5360 2455 5406
rect 2255 5317 2455 5360
rect 2255 5074 2455 5117
rect 2255 5028 2268 5074
rect 2442 5028 2455 5074
rect 2255 5015 2455 5028
rect 2535 5406 2735 5419
rect 2535 5360 2548 5406
rect 2722 5360 2735 5406
rect 2535 5317 2735 5360
rect 2535 5074 2735 5117
rect 2535 5028 2548 5074
rect 2722 5028 2735 5074
rect 2535 5015 2735 5028
rect 2815 5406 3015 5419
rect 2815 5360 2828 5406
rect 3002 5360 3015 5406
rect 2815 5317 3015 5360
rect 2815 5074 3015 5117
rect 2815 5028 2828 5074
rect 3002 5028 3015 5074
rect 2815 5015 3015 5028
rect 3095 5406 3295 5419
rect 3095 5360 3108 5406
rect 3282 5360 3295 5406
rect 3095 5317 3295 5360
rect 3095 5074 3295 5117
rect 3095 5028 3108 5074
rect 3282 5028 3295 5074
rect 3095 5015 3295 5028
rect 3375 5406 3575 5419
rect 3375 5360 3388 5406
rect 3562 5360 3575 5406
rect 3375 5317 3575 5360
rect 3375 5074 3575 5117
rect 3375 5028 3388 5074
rect 3562 5028 3575 5074
rect 3375 5015 3575 5028
rect 3655 5406 3855 5419
rect 3655 5360 3668 5406
rect 3842 5360 3855 5406
rect 3655 5317 3855 5360
rect 3655 5074 3855 5117
rect 3655 5028 3668 5074
rect 3842 5028 3855 5074
rect 3655 5015 3855 5028
rect 3935 5406 4135 5419
rect 3935 5360 3948 5406
rect 4122 5360 4135 5406
rect 3935 5317 4135 5360
rect 3935 5074 4135 5117
rect 3935 5028 3948 5074
rect 4122 5028 4135 5074
rect 3935 5015 4135 5028
rect 4215 5406 4415 5419
rect 4215 5360 4228 5406
rect 4402 5360 4415 5406
rect 4215 5317 4415 5360
rect 4215 5074 4415 5117
rect 4215 5028 4228 5074
rect 4402 5028 4415 5074
rect 4215 5015 4415 5028
rect 4495 5406 4695 5419
rect 4495 5360 4508 5406
rect 4682 5360 4695 5406
rect 4495 5317 4695 5360
rect 4495 5074 4695 5117
rect 4495 5028 4508 5074
rect 4682 5028 4695 5074
rect 4495 5015 4695 5028
rect 4775 5406 4975 5419
rect 4775 5360 4788 5406
rect 4962 5360 4975 5406
rect 4775 5317 4975 5360
rect 4775 5074 4975 5117
rect 4775 5028 4788 5074
rect 4962 5028 4975 5074
rect 4775 5015 4975 5028
rect 5055 5406 5255 5419
rect 5055 5360 5068 5406
rect 5242 5360 5255 5406
rect 5055 5317 5255 5360
rect 5055 5074 5255 5117
rect 5055 5028 5068 5074
rect 5242 5028 5255 5074
rect 5055 5015 5255 5028
rect 5335 5406 5535 5419
rect 5335 5360 5348 5406
rect 5522 5360 5535 5406
rect 5335 5317 5535 5360
rect 5335 5074 5535 5117
rect 5335 5028 5348 5074
rect 5522 5028 5535 5074
rect 5335 5015 5535 5028
rect 5615 5406 5815 5419
rect 5615 5360 5628 5406
rect 5802 5360 5815 5406
rect 5615 5317 5815 5360
rect 5615 5074 5815 5117
rect 5615 5028 5628 5074
rect 5802 5028 5815 5074
rect 5615 5015 5815 5028
rect 5895 5406 6095 5419
rect 5895 5360 5908 5406
rect 6082 5360 6095 5406
rect 5895 5317 6095 5360
rect 5895 5074 6095 5117
rect 5895 5028 5908 5074
rect 6082 5028 6095 5074
rect 5895 5015 6095 5028
rect 6175 5406 6375 5419
rect 6175 5360 6188 5406
rect 6362 5360 6375 5406
rect 6175 5317 6375 5360
rect 6175 5074 6375 5117
rect 6175 5028 6188 5074
rect 6362 5028 6375 5074
rect 6175 5015 6375 5028
rect 6455 5406 6655 5419
rect 6455 5360 6468 5406
rect 6642 5360 6655 5406
rect 6455 5317 6655 5360
rect 6455 5074 6655 5117
rect 6455 5028 6468 5074
rect 6642 5028 6655 5074
rect 6455 5015 6655 5028
rect 6735 5406 6935 5419
rect 6735 5360 6748 5406
rect 6922 5360 6935 5406
rect 6735 5317 6935 5360
rect 6735 5074 6935 5117
rect 6735 5028 6748 5074
rect 6922 5028 6935 5074
rect 6735 5015 6935 5028
rect 7015 5406 7215 5419
rect 7015 5360 7028 5406
rect 7202 5360 7215 5406
rect 7015 5317 7215 5360
rect 7015 5074 7215 5117
rect 7015 5028 7028 5074
rect 7202 5028 7215 5074
rect 7015 5015 7215 5028
rect 7295 5406 7495 5419
rect 7295 5360 7308 5406
rect 7482 5360 7495 5406
rect 7295 5317 7495 5360
rect 7295 5074 7495 5117
rect 7295 5028 7308 5074
rect 7482 5028 7495 5074
rect 7295 5015 7495 5028
rect 7575 5406 7775 5419
rect 7575 5360 7588 5406
rect 7762 5360 7775 5406
rect 7575 5317 7775 5360
rect 7575 5074 7775 5117
rect 7575 5028 7588 5074
rect 7762 5028 7775 5074
rect 7575 5015 7775 5028
rect 7855 5406 8055 5419
rect 7855 5360 7868 5406
rect 8042 5360 8055 5406
rect 7855 5317 8055 5360
rect 7855 5074 8055 5117
rect 7855 5028 7868 5074
rect 8042 5028 8055 5074
rect 7855 5015 8055 5028
rect 8135 5406 8335 5419
rect 8135 5360 8148 5406
rect 8322 5360 8335 5406
rect 8135 5317 8335 5360
rect 8135 5074 8335 5117
rect 8135 5028 8148 5074
rect 8322 5028 8335 5074
rect 8135 5015 8335 5028
rect 8415 5406 8615 5419
rect 8415 5360 8428 5406
rect 8602 5360 8615 5406
rect 8415 5317 8615 5360
rect 8415 5074 8615 5117
rect 8415 5028 8428 5074
rect 8602 5028 8615 5074
rect 8415 5015 8615 5028
rect 8695 5406 8895 5419
rect 8695 5360 8708 5406
rect 8882 5360 8895 5406
rect 8695 5317 8895 5360
rect 8695 5074 8895 5117
rect 8695 5028 8708 5074
rect 8882 5028 8895 5074
rect 8695 5015 8895 5028
rect 8975 5406 9175 5419
rect 8975 5360 8988 5406
rect 9162 5360 9175 5406
rect 8975 5317 9175 5360
rect 8975 5074 9175 5117
rect 8975 5028 8988 5074
rect 9162 5028 9175 5074
rect 8975 5015 9175 5028
rect 9255 5406 9455 5419
rect 9255 5360 9268 5406
rect 9442 5360 9455 5406
rect 9255 5317 9455 5360
rect 9255 5074 9455 5117
rect 9255 5028 9268 5074
rect 9442 5028 9455 5074
rect 9255 5015 9455 5028
rect 9535 5406 9735 5419
rect 9535 5360 9548 5406
rect 9722 5360 9735 5406
rect 9535 5317 9735 5360
rect 9535 5074 9735 5117
rect 9535 5028 9548 5074
rect 9722 5028 9735 5074
rect 9535 5015 9735 5028
rect 295 4754 495 4767
rect 295 4708 308 4754
rect 482 4708 495 4754
rect 295 4665 495 4708
rect 295 4422 495 4465
rect 295 4376 308 4422
rect 482 4376 495 4422
rect 295 4363 495 4376
rect 575 4754 775 4767
rect 575 4708 588 4754
rect 762 4708 775 4754
rect 575 4665 775 4708
rect 575 4422 775 4465
rect 575 4376 588 4422
rect 762 4376 775 4422
rect 575 4363 775 4376
rect 855 4754 1055 4767
rect 855 4708 868 4754
rect 1042 4708 1055 4754
rect 855 4665 1055 4708
rect 855 4422 1055 4465
rect 855 4376 868 4422
rect 1042 4376 1055 4422
rect 855 4363 1055 4376
rect 1135 4754 1335 4767
rect 1135 4708 1148 4754
rect 1322 4708 1335 4754
rect 1135 4665 1335 4708
rect 1135 4422 1335 4465
rect 1135 4376 1148 4422
rect 1322 4376 1335 4422
rect 1135 4363 1335 4376
rect 1415 4754 1615 4767
rect 1415 4708 1428 4754
rect 1602 4708 1615 4754
rect 1415 4665 1615 4708
rect 1415 4422 1615 4465
rect 1415 4376 1428 4422
rect 1602 4376 1615 4422
rect 1415 4363 1615 4376
rect 1695 4754 1895 4767
rect 1695 4708 1708 4754
rect 1882 4708 1895 4754
rect 1695 4665 1895 4708
rect 1695 4422 1895 4465
rect 1695 4376 1708 4422
rect 1882 4376 1895 4422
rect 1695 4363 1895 4376
rect 1975 4754 2175 4767
rect 1975 4708 1988 4754
rect 2162 4708 2175 4754
rect 1975 4665 2175 4708
rect 1975 4422 2175 4465
rect 1975 4376 1988 4422
rect 2162 4376 2175 4422
rect 1975 4363 2175 4376
rect 2255 4754 2455 4767
rect 2255 4708 2268 4754
rect 2442 4708 2455 4754
rect 2255 4665 2455 4708
rect 2255 4422 2455 4465
rect 2255 4376 2268 4422
rect 2442 4376 2455 4422
rect 2255 4363 2455 4376
rect 2535 4754 2735 4767
rect 2535 4708 2548 4754
rect 2722 4708 2735 4754
rect 2535 4665 2735 4708
rect 2535 4422 2735 4465
rect 2535 4376 2548 4422
rect 2722 4376 2735 4422
rect 2535 4363 2735 4376
rect 2815 4754 3015 4767
rect 2815 4708 2828 4754
rect 3002 4708 3015 4754
rect 2815 4665 3015 4708
rect 2815 4422 3015 4465
rect 2815 4376 2828 4422
rect 3002 4376 3015 4422
rect 2815 4363 3015 4376
rect 3095 4754 3295 4767
rect 3095 4708 3108 4754
rect 3282 4708 3295 4754
rect 3095 4665 3295 4708
rect 3095 4422 3295 4465
rect 3095 4376 3108 4422
rect 3282 4376 3295 4422
rect 3095 4363 3295 4376
rect 3375 4754 3575 4767
rect 3375 4708 3388 4754
rect 3562 4708 3575 4754
rect 3375 4665 3575 4708
rect 3375 4422 3575 4465
rect 3375 4376 3388 4422
rect 3562 4376 3575 4422
rect 3375 4363 3575 4376
rect 3655 4754 3855 4767
rect 3655 4708 3668 4754
rect 3842 4708 3855 4754
rect 3655 4665 3855 4708
rect 3655 4422 3855 4465
rect 3655 4376 3668 4422
rect 3842 4376 3855 4422
rect 3655 4363 3855 4376
rect 3935 4754 4135 4767
rect 3935 4708 3948 4754
rect 4122 4708 4135 4754
rect 3935 4665 4135 4708
rect 3935 4422 4135 4465
rect 3935 4376 3948 4422
rect 4122 4376 4135 4422
rect 3935 4363 4135 4376
rect 4215 4754 4415 4767
rect 4215 4708 4228 4754
rect 4402 4708 4415 4754
rect 4215 4665 4415 4708
rect 4215 4422 4415 4465
rect 4215 4376 4228 4422
rect 4402 4376 4415 4422
rect 4215 4363 4415 4376
rect 4495 4754 4695 4767
rect 4495 4708 4508 4754
rect 4682 4708 4695 4754
rect 4495 4665 4695 4708
rect 4495 4422 4695 4465
rect 4495 4376 4508 4422
rect 4682 4376 4695 4422
rect 4495 4363 4695 4376
rect 4775 4754 4975 4767
rect 4775 4708 4788 4754
rect 4962 4708 4975 4754
rect 4775 4665 4975 4708
rect 4775 4422 4975 4465
rect 4775 4376 4788 4422
rect 4962 4376 4975 4422
rect 4775 4363 4975 4376
rect 5055 4754 5255 4767
rect 5055 4708 5068 4754
rect 5242 4708 5255 4754
rect 5055 4665 5255 4708
rect 5055 4422 5255 4465
rect 5055 4376 5068 4422
rect 5242 4376 5255 4422
rect 5055 4363 5255 4376
rect 5335 4754 5535 4767
rect 5335 4708 5348 4754
rect 5522 4708 5535 4754
rect 5335 4665 5535 4708
rect 5335 4422 5535 4465
rect 5335 4376 5348 4422
rect 5522 4376 5535 4422
rect 5335 4363 5535 4376
rect 5615 4754 5815 4767
rect 5615 4708 5628 4754
rect 5802 4708 5815 4754
rect 5615 4665 5815 4708
rect 5615 4422 5815 4465
rect 5615 4376 5628 4422
rect 5802 4376 5815 4422
rect 5615 4363 5815 4376
rect 5895 4754 6095 4767
rect 5895 4708 5908 4754
rect 6082 4708 6095 4754
rect 5895 4665 6095 4708
rect 5895 4422 6095 4465
rect 5895 4376 5908 4422
rect 6082 4376 6095 4422
rect 5895 4363 6095 4376
rect 6175 4754 6375 4767
rect 6175 4708 6188 4754
rect 6362 4708 6375 4754
rect 6175 4665 6375 4708
rect 6175 4422 6375 4465
rect 6175 4376 6188 4422
rect 6362 4376 6375 4422
rect 6175 4363 6375 4376
rect 6455 4754 6655 4767
rect 6455 4708 6468 4754
rect 6642 4708 6655 4754
rect 6455 4665 6655 4708
rect 6455 4422 6655 4465
rect 6455 4376 6468 4422
rect 6642 4376 6655 4422
rect 6455 4363 6655 4376
rect 6735 4754 6935 4767
rect 6735 4708 6748 4754
rect 6922 4708 6935 4754
rect 6735 4665 6935 4708
rect 6735 4422 6935 4465
rect 6735 4376 6748 4422
rect 6922 4376 6935 4422
rect 6735 4363 6935 4376
rect 7015 4754 7215 4767
rect 7015 4708 7028 4754
rect 7202 4708 7215 4754
rect 7015 4665 7215 4708
rect 7015 4422 7215 4465
rect 7015 4376 7028 4422
rect 7202 4376 7215 4422
rect 7015 4363 7215 4376
rect 7295 4754 7495 4767
rect 7295 4708 7308 4754
rect 7482 4708 7495 4754
rect 7295 4665 7495 4708
rect 7295 4422 7495 4465
rect 7295 4376 7308 4422
rect 7482 4376 7495 4422
rect 7295 4363 7495 4376
rect 7575 4754 7775 4767
rect 7575 4708 7588 4754
rect 7762 4708 7775 4754
rect 7575 4665 7775 4708
rect 7575 4422 7775 4465
rect 7575 4376 7588 4422
rect 7762 4376 7775 4422
rect 7575 4363 7775 4376
rect 7855 4754 8055 4767
rect 7855 4708 7868 4754
rect 8042 4708 8055 4754
rect 7855 4665 8055 4708
rect 7855 4422 8055 4465
rect 7855 4376 7868 4422
rect 8042 4376 8055 4422
rect 7855 4363 8055 4376
rect 8135 4754 8335 4767
rect 8135 4708 8148 4754
rect 8322 4708 8335 4754
rect 8135 4665 8335 4708
rect 8135 4422 8335 4465
rect 8135 4376 8148 4422
rect 8322 4376 8335 4422
rect 8135 4363 8335 4376
rect 8415 4754 8615 4767
rect 8415 4708 8428 4754
rect 8602 4708 8615 4754
rect 8415 4665 8615 4708
rect 8415 4422 8615 4465
rect 8415 4376 8428 4422
rect 8602 4376 8615 4422
rect 8415 4363 8615 4376
rect 8695 4754 8895 4767
rect 8695 4708 8708 4754
rect 8882 4708 8895 4754
rect 8695 4665 8895 4708
rect 8695 4422 8895 4465
rect 8695 4376 8708 4422
rect 8882 4376 8895 4422
rect 8695 4363 8895 4376
rect 8975 4754 9175 4767
rect 8975 4708 8988 4754
rect 9162 4708 9175 4754
rect 8975 4665 9175 4708
rect 8975 4422 9175 4465
rect 8975 4376 8988 4422
rect 9162 4376 9175 4422
rect 8975 4363 9175 4376
rect 9255 4754 9455 4767
rect 9255 4708 9268 4754
rect 9442 4708 9455 4754
rect 9255 4665 9455 4708
rect 9255 4422 9455 4465
rect 9255 4376 9268 4422
rect 9442 4376 9455 4422
rect 9255 4363 9455 4376
rect 9535 4754 9735 4767
rect 9535 4708 9548 4754
rect 9722 4708 9735 4754
rect 9535 4665 9735 4708
rect 9535 4422 9735 4465
rect 9535 4376 9548 4422
rect 9722 4376 9735 4422
rect 9535 4363 9735 4376
rect 295 4102 495 4115
rect 295 4056 308 4102
rect 482 4056 495 4102
rect 295 4013 495 4056
rect 295 3770 495 3813
rect 295 3724 308 3770
rect 482 3724 495 3770
rect 295 3711 495 3724
rect 575 4102 775 4115
rect 575 4056 588 4102
rect 762 4056 775 4102
rect 575 4013 775 4056
rect 575 3770 775 3813
rect 575 3724 588 3770
rect 762 3724 775 3770
rect 575 3711 775 3724
rect 855 4102 1055 4115
rect 855 4056 868 4102
rect 1042 4056 1055 4102
rect 855 4013 1055 4056
rect 855 3770 1055 3813
rect 855 3724 868 3770
rect 1042 3724 1055 3770
rect 855 3711 1055 3724
rect 1135 4102 1335 4115
rect 1135 4056 1148 4102
rect 1322 4056 1335 4102
rect 1135 4013 1335 4056
rect 1135 3770 1335 3813
rect 1135 3724 1148 3770
rect 1322 3724 1335 3770
rect 1135 3711 1335 3724
rect 1415 4102 1615 4115
rect 1415 4056 1428 4102
rect 1602 4056 1615 4102
rect 1415 4013 1615 4056
rect 1415 3770 1615 3813
rect 1415 3724 1428 3770
rect 1602 3724 1615 3770
rect 1415 3711 1615 3724
rect 1695 4102 1895 4115
rect 1695 4056 1708 4102
rect 1882 4056 1895 4102
rect 1695 4013 1895 4056
rect 1695 3770 1895 3813
rect 1695 3724 1708 3770
rect 1882 3724 1895 3770
rect 1695 3711 1895 3724
rect 1975 4102 2175 4115
rect 1975 4056 1988 4102
rect 2162 4056 2175 4102
rect 1975 4013 2175 4056
rect 1975 3770 2175 3813
rect 1975 3724 1988 3770
rect 2162 3724 2175 3770
rect 1975 3711 2175 3724
rect 2255 4102 2455 4115
rect 2255 4056 2268 4102
rect 2442 4056 2455 4102
rect 2255 4013 2455 4056
rect 2255 3770 2455 3813
rect 2255 3724 2268 3770
rect 2442 3724 2455 3770
rect 2255 3711 2455 3724
rect 2535 4102 2735 4115
rect 2535 4056 2548 4102
rect 2722 4056 2735 4102
rect 2535 4013 2735 4056
rect 2535 3770 2735 3813
rect 2535 3724 2548 3770
rect 2722 3724 2735 3770
rect 2535 3711 2735 3724
rect 2815 4102 3015 4115
rect 2815 4056 2828 4102
rect 3002 4056 3015 4102
rect 2815 4013 3015 4056
rect 2815 3770 3015 3813
rect 2815 3724 2828 3770
rect 3002 3724 3015 3770
rect 2815 3711 3015 3724
rect 3095 4102 3295 4115
rect 3095 4056 3108 4102
rect 3282 4056 3295 4102
rect 3095 4013 3295 4056
rect 3095 3770 3295 3813
rect 3095 3724 3108 3770
rect 3282 3724 3295 3770
rect 3095 3711 3295 3724
rect 3375 4102 3575 4115
rect 3375 4056 3388 4102
rect 3562 4056 3575 4102
rect 3375 4013 3575 4056
rect 3375 3770 3575 3813
rect 3375 3724 3388 3770
rect 3562 3724 3575 3770
rect 3375 3711 3575 3724
rect 3655 4102 3855 4115
rect 3655 4056 3668 4102
rect 3842 4056 3855 4102
rect 3655 4013 3855 4056
rect 3655 3770 3855 3813
rect 3655 3724 3668 3770
rect 3842 3724 3855 3770
rect 3655 3711 3855 3724
rect 3935 4102 4135 4115
rect 3935 4056 3948 4102
rect 4122 4056 4135 4102
rect 3935 4013 4135 4056
rect 3935 3770 4135 3813
rect 3935 3724 3948 3770
rect 4122 3724 4135 3770
rect 3935 3711 4135 3724
rect 4215 4102 4415 4115
rect 4215 4056 4228 4102
rect 4402 4056 4415 4102
rect 4215 4013 4415 4056
rect 4215 3770 4415 3813
rect 4215 3724 4228 3770
rect 4402 3724 4415 3770
rect 4215 3711 4415 3724
rect 4495 4102 4695 4115
rect 4495 4056 4508 4102
rect 4682 4056 4695 4102
rect 4495 4013 4695 4056
rect 4495 3770 4695 3813
rect 4495 3724 4508 3770
rect 4682 3724 4695 3770
rect 4495 3711 4695 3724
rect 4775 4102 4975 4115
rect 4775 4056 4788 4102
rect 4962 4056 4975 4102
rect 4775 4013 4975 4056
rect 4775 3770 4975 3813
rect 4775 3724 4788 3770
rect 4962 3724 4975 3770
rect 4775 3711 4975 3724
rect 5055 4102 5255 4115
rect 5055 4056 5068 4102
rect 5242 4056 5255 4102
rect 5055 4013 5255 4056
rect 5055 3770 5255 3813
rect 5055 3724 5068 3770
rect 5242 3724 5255 3770
rect 5055 3711 5255 3724
rect 5335 4102 5535 4115
rect 5335 4056 5348 4102
rect 5522 4056 5535 4102
rect 5335 4013 5535 4056
rect 5335 3770 5535 3813
rect 5335 3724 5348 3770
rect 5522 3724 5535 3770
rect 5335 3711 5535 3724
rect 5615 4102 5815 4115
rect 5615 4056 5628 4102
rect 5802 4056 5815 4102
rect 5615 4013 5815 4056
rect 5615 3770 5815 3813
rect 5615 3724 5628 3770
rect 5802 3724 5815 3770
rect 5615 3711 5815 3724
rect 5895 4102 6095 4115
rect 5895 4056 5908 4102
rect 6082 4056 6095 4102
rect 5895 4013 6095 4056
rect 5895 3770 6095 3813
rect 5895 3724 5908 3770
rect 6082 3724 6095 3770
rect 5895 3711 6095 3724
rect 6175 4102 6375 4115
rect 6175 4056 6188 4102
rect 6362 4056 6375 4102
rect 6175 4013 6375 4056
rect 6175 3770 6375 3813
rect 6175 3724 6188 3770
rect 6362 3724 6375 3770
rect 6175 3711 6375 3724
rect 6455 4102 6655 4115
rect 6455 4056 6468 4102
rect 6642 4056 6655 4102
rect 6455 4013 6655 4056
rect 6455 3770 6655 3813
rect 6455 3724 6468 3770
rect 6642 3724 6655 3770
rect 6455 3711 6655 3724
rect 6735 4102 6935 4115
rect 6735 4056 6748 4102
rect 6922 4056 6935 4102
rect 6735 4013 6935 4056
rect 6735 3770 6935 3813
rect 6735 3724 6748 3770
rect 6922 3724 6935 3770
rect 6735 3711 6935 3724
rect 7015 4102 7215 4115
rect 7015 4056 7028 4102
rect 7202 4056 7215 4102
rect 7015 4013 7215 4056
rect 7015 3770 7215 3813
rect 7015 3724 7028 3770
rect 7202 3724 7215 3770
rect 7015 3711 7215 3724
rect 7295 4102 7495 4115
rect 7295 4056 7308 4102
rect 7482 4056 7495 4102
rect 7295 4013 7495 4056
rect 7295 3770 7495 3813
rect 7295 3724 7308 3770
rect 7482 3724 7495 3770
rect 7295 3711 7495 3724
rect 7575 4102 7775 4115
rect 7575 4056 7588 4102
rect 7762 4056 7775 4102
rect 7575 4013 7775 4056
rect 7575 3770 7775 3813
rect 7575 3724 7588 3770
rect 7762 3724 7775 3770
rect 7575 3711 7775 3724
rect 7855 4102 8055 4115
rect 7855 4056 7868 4102
rect 8042 4056 8055 4102
rect 7855 4013 8055 4056
rect 7855 3770 8055 3813
rect 7855 3724 7868 3770
rect 8042 3724 8055 3770
rect 7855 3711 8055 3724
rect 8135 4102 8335 4115
rect 8135 4056 8148 4102
rect 8322 4056 8335 4102
rect 8135 4013 8335 4056
rect 8135 3770 8335 3813
rect 8135 3724 8148 3770
rect 8322 3724 8335 3770
rect 8135 3711 8335 3724
rect 8415 4102 8615 4115
rect 8415 4056 8428 4102
rect 8602 4056 8615 4102
rect 8415 4013 8615 4056
rect 8415 3770 8615 3813
rect 8415 3724 8428 3770
rect 8602 3724 8615 3770
rect 8415 3711 8615 3724
rect 8695 4102 8895 4115
rect 8695 4056 8708 4102
rect 8882 4056 8895 4102
rect 8695 4013 8895 4056
rect 8695 3770 8895 3813
rect 8695 3724 8708 3770
rect 8882 3724 8895 3770
rect 8695 3711 8895 3724
rect 8975 4102 9175 4115
rect 8975 4056 8988 4102
rect 9162 4056 9175 4102
rect 8975 4013 9175 4056
rect 8975 3770 9175 3813
rect 8975 3724 8988 3770
rect 9162 3724 9175 3770
rect 8975 3711 9175 3724
rect 9255 4102 9455 4115
rect 9255 4056 9268 4102
rect 9442 4056 9455 4102
rect 9255 4013 9455 4056
rect 9255 3770 9455 3813
rect 9255 3724 9268 3770
rect 9442 3724 9455 3770
rect 9255 3711 9455 3724
rect 9535 4102 9735 4115
rect 9535 4056 9548 4102
rect 9722 4056 9735 4102
rect 9535 4013 9735 4056
rect 9535 3770 9735 3813
rect 9535 3724 9548 3770
rect 9722 3724 9735 3770
rect 9535 3711 9735 3724
rect 295 2977 495 2990
rect 295 2931 308 2977
rect 482 2931 495 2977
rect 295 2888 495 2931
rect 295 2645 495 2688
rect 295 2599 308 2645
rect 482 2599 495 2645
rect 295 2586 495 2599
rect 575 2977 775 2990
rect 575 2931 588 2977
rect 762 2931 775 2977
rect 575 2888 775 2931
rect 575 2645 775 2688
rect 575 2599 588 2645
rect 762 2599 775 2645
rect 575 2586 775 2599
rect 855 2977 1055 2990
rect 855 2931 868 2977
rect 1042 2931 1055 2977
rect 855 2888 1055 2931
rect 855 2645 1055 2688
rect 855 2599 868 2645
rect 1042 2599 1055 2645
rect 855 2586 1055 2599
rect 1135 2977 1335 2990
rect 1135 2931 1148 2977
rect 1322 2931 1335 2977
rect 1135 2888 1335 2931
rect 1135 2645 1335 2688
rect 1135 2599 1148 2645
rect 1322 2599 1335 2645
rect 1135 2586 1335 2599
rect 1415 2977 1615 2990
rect 1415 2931 1428 2977
rect 1602 2931 1615 2977
rect 1415 2888 1615 2931
rect 1415 2645 1615 2688
rect 1415 2599 1428 2645
rect 1602 2599 1615 2645
rect 1415 2586 1615 2599
rect 1695 2977 1895 2990
rect 1695 2931 1708 2977
rect 1882 2931 1895 2977
rect 1695 2888 1895 2931
rect 1695 2645 1895 2688
rect 1695 2599 1708 2645
rect 1882 2599 1895 2645
rect 1695 2586 1895 2599
rect 1975 2977 2175 2990
rect 1975 2931 1988 2977
rect 2162 2931 2175 2977
rect 1975 2888 2175 2931
rect 1975 2645 2175 2688
rect 1975 2599 1988 2645
rect 2162 2599 2175 2645
rect 1975 2586 2175 2599
rect 2255 2977 2455 2990
rect 2255 2931 2268 2977
rect 2442 2931 2455 2977
rect 2255 2888 2455 2931
rect 2255 2645 2455 2688
rect 2255 2599 2268 2645
rect 2442 2599 2455 2645
rect 2255 2586 2455 2599
rect 2535 2977 2735 2990
rect 2535 2931 2548 2977
rect 2722 2931 2735 2977
rect 2535 2888 2735 2931
rect 2535 2645 2735 2688
rect 2535 2599 2548 2645
rect 2722 2599 2735 2645
rect 2535 2586 2735 2599
rect 2815 2977 3015 2990
rect 2815 2931 2828 2977
rect 3002 2931 3015 2977
rect 2815 2888 3015 2931
rect 2815 2645 3015 2688
rect 2815 2599 2828 2645
rect 3002 2599 3015 2645
rect 2815 2586 3015 2599
rect 3095 2977 3295 2990
rect 3095 2931 3108 2977
rect 3282 2931 3295 2977
rect 3095 2888 3295 2931
rect 3095 2645 3295 2688
rect 3095 2599 3108 2645
rect 3282 2599 3295 2645
rect 3095 2586 3295 2599
rect 3375 2977 3575 2990
rect 3375 2931 3388 2977
rect 3562 2931 3575 2977
rect 3375 2888 3575 2931
rect 3375 2645 3575 2688
rect 3375 2599 3388 2645
rect 3562 2599 3575 2645
rect 3375 2586 3575 2599
rect 3655 2977 3855 2990
rect 3655 2931 3668 2977
rect 3842 2931 3855 2977
rect 3655 2888 3855 2931
rect 3655 2645 3855 2688
rect 3655 2599 3668 2645
rect 3842 2599 3855 2645
rect 3655 2586 3855 2599
rect 3935 2977 4135 2990
rect 3935 2931 3948 2977
rect 4122 2931 4135 2977
rect 3935 2888 4135 2931
rect 3935 2645 4135 2688
rect 3935 2599 3948 2645
rect 4122 2599 4135 2645
rect 3935 2586 4135 2599
rect 4215 2977 4415 2990
rect 4215 2931 4228 2977
rect 4402 2931 4415 2977
rect 4215 2888 4415 2931
rect 4215 2645 4415 2688
rect 4215 2599 4228 2645
rect 4402 2599 4415 2645
rect 4215 2586 4415 2599
rect 4495 2977 4695 2990
rect 4495 2931 4508 2977
rect 4682 2931 4695 2977
rect 4495 2888 4695 2931
rect 4495 2645 4695 2688
rect 4495 2599 4508 2645
rect 4682 2599 4695 2645
rect 4495 2586 4695 2599
rect 4775 2977 4975 2990
rect 4775 2931 4788 2977
rect 4962 2931 4975 2977
rect 4775 2888 4975 2931
rect 4775 2645 4975 2688
rect 4775 2599 4788 2645
rect 4962 2599 4975 2645
rect 4775 2586 4975 2599
rect 5055 2977 5255 2990
rect 5055 2931 5068 2977
rect 5242 2931 5255 2977
rect 5055 2888 5255 2931
rect 5055 2645 5255 2688
rect 5055 2599 5068 2645
rect 5242 2599 5255 2645
rect 5055 2586 5255 2599
rect 5335 2977 5535 2990
rect 5335 2931 5348 2977
rect 5522 2931 5535 2977
rect 5335 2888 5535 2931
rect 5335 2645 5535 2688
rect 5335 2599 5348 2645
rect 5522 2599 5535 2645
rect 5335 2586 5535 2599
rect 5615 2977 5815 2990
rect 5615 2931 5628 2977
rect 5802 2931 5815 2977
rect 5615 2888 5815 2931
rect 5615 2645 5815 2688
rect 5615 2599 5628 2645
rect 5802 2599 5815 2645
rect 5615 2586 5815 2599
rect 5895 2977 6095 2990
rect 5895 2931 5908 2977
rect 6082 2931 6095 2977
rect 5895 2888 6095 2931
rect 5895 2645 6095 2688
rect 5895 2599 5908 2645
rect 6082 2599 6095 2645
rect 5895 2586 6095 2599
rect 6175 2977 6375 2990
rect 6175 2931 6188 2977
rect 6362 2931 6375 2977
rect 6175 2888 6375 2931
rect 6175 2645 6375 2688
rect 6175 2599 6188 2645
rect 6362 2599 6375 2645
rect 6175 2586 6375 2599
rect 6455 2977 6655 2990
rect 6455 2931 6468 2977
rect 6642 2931 6655 2977
rect 6455 2888 6655 2931
rect 6455 2645 6655 2688
rect 6455 2599 6468 2645
rect 6642 2599 6655 2645
rect 6455 2586 6655 2599
rect 6735 2977 6935 2990
rect 6735 2931 6748 2977
rect 6922 2931 6935 2977
rect 6735 2888 6935 2931
rect 6735 2645 6935 2688
rect 6735 2599 6748 2645
rect 6922 2599 6935 2645
rect 6735 2586 6935 2599
rect 7015 2977 7215 2990
rect 7015 2931 7028 2977
rect 7202 2931 7215 2977
rect 7015 2888 7215 2931
rect 7015 2645 7215 2688
rect 7015 2599 7028 2645
rect 7202 2599 7215 2645
rect 7015 2586 7215 2599
rect 7295 2977 7495 2990
rect 7295 2931 7308 2977
rect 7482 2931 7495 2977
rect 7295 2888 7495 2931
rect 7295 2645 7495 2688
rect 7295 2599 7308 2645
rect 7482 2599 7495 2645
rect 7295 2586 7495 2599
rect 7575 2977 7775 2990
rect 7575 2931 7588 2977
rect 7762 2931 7775 2977
rect 7575 2888 7775 2931
rect 7575 2645 7775 2688
rect 7575 2599 7588 2645
rect 7762 2599 7775 2645
rect 7575 2586 7775 2599
rect 7855 2977 8055 2990
rect 7855 2931 7868 2977
rect 8042 2931 8055 2977
rect 7855 2888 8055 2931
rect 7855 2645 8055 2688
rect 7855 2599 7868 2645
rect 8042 2599 8055 2645
rect 7855 2586 8055 2599
rect 8135 2977 8335 2990
rect 8135 2931 8148 2977
rect 8322 2931 8335 2977
rect 8135 2888 8335 2931
rect 8135 2645 8335 2688
rect 8135 2599 8148 2645
rect 8322 2599 8335 2645
rect 8135 2586 8335 2599
rect 8415 2977 8615 2990
rect 8415 2931 8428 2977
rect 8602 2931 8615 2977
rect 8415 2888 8615 2931
rect 8415 2645 8615 2688
rect 8415 2599 8428 2645
rect 8602 2599 8615 2645
rect 8415 2586 8615 2599
rect 8695 2977 8895 2990
rect 8695 2931 8708 2977
rect 8882 2931 8895 2977
rect 8695 2888 8895 2931
rect 8695 2645 8895 2688
rect 8695 2599 8708 2645
rect 8882 2599 8895 2645
rect 8695 2586 8895 2599
rect 8975 2977 9175 2990
rect 8975 2931 8988 2977
rect 9162 2931 9175 2977
rect 8975 2888 9175 2931
rect 8975 2645 9175 2688
rect 8975 2599 8988 2645
rect 9162 2599 9175 2645
rect 8975 2586 9175 2599
rect 9255 2977 9455 2990
rect 9255 2931 9268 2977
rect 9442 2931 9455 2977
rect 9255 2888 9455 2931
rect 9255 2645 9455 2688
rect 9255 2599 9268 2645
rect 9442 2599 9455 2645
rect 9255 2586 9455 2599
rect 9535 2977 9735 2990
rect 9535 2931 9548 2977
rect 9722 2931 9735 2977
rect 9535 2888 9735 2931
rect 9535 2645 9735 2688
rect 9535 2599 9548 2645
rect 9722 2599 9735 2645
rect 9535 2586 9735 2599
rect 295 2325 495 2338
rect 295 2279 308 2325
rect 482 2279 495 2325
rect 295 2236 495 2279
rect 295 1993 495 2036
rect 295 1947 308 1993
rect 482 1947 495 1993
rect 295 1934 495 1947
rect 575 2325 775 2338
rect 575 2279 588 2325
rect 762 2279 775 2325
rect 575 2236 775 2279
rect 575 1993 775 2036
rect 575 1947 588 1993
rect 762 1947 775 1993
rect 575 1934 775 1947
rect 855 2325 1055 2338
rect 855 2279 868 2325
rect 1042 2279 1055 2325
rect 855 2236 1055 2279
rect 855 1993 1055 2036
rect 855 1947 868 1993
rect 1042 1947 1055 1993
rect 855 1934 1055 1947
rect 1135 2325 1335 2338
rect 1135 2279 1148 2325
rect 1322 2279 1335 2325
rect 1135 2236 1335 2279
rect 1135 1993 1335 2036
rect 1135 1947 1148 1993
rect 1322 1947 1335 1993
rect 1135 1934 1335 1947
rect 1415 2325 1615 2338
rect 1415 2279 1428 2325
rect 1602 2279 1615 2325
rect 1415 2236 1615 2279
rect 1415 1993 1615 2036
rect 1415 1947 1428 1993
rect 1602 1947 1615 1993
rect 1415 1934 1615 1947
rect 1695 2325 1895 2338
rect 1695 2279 1708 2325
rect 1882 2279 1895 2325
rect 1695 2236 1895 2279
rect 1695 1993 1895 2036
rect 1695 1947 1708 1993
rect 1882 1947 1895 1993
rect 1695 1934 1895 1947
rect 1975 2325 2175 2338
rect 1975 2279 1988 2325
rect 2162 2279 2175 2325
rect 1975 2236 2175 2279
rect 1975 1993 2175 2036
rect 1975 1947 1988 1993
rect 2162 1947 2175 1993
rect 1975 1934 2175 1947
rect 2255 2325 2455 2338
rect 2255 2279 2268 2325
rect 2442 2279 2455 2325
rect 2255 2236 2455 2279
rect 2255 1993 2455 2036
rect 2255 1947 2268 1993
rect 2442 1947 2455 1993
rect 2255 1934 2455 1947
rect 2535 2325 2735 2338
rect 2535 2279 2548 2325
rect 2722 2279 2735 2325
rect 2535 2236 2735 2279
rect 2535 1993 2735 2036
rect 2535 1947 2548 1993
rect 2722 1947 2735 1993
rect 2535 1934 2735 1947
rect 2815 2325 3015 2338
rect 2815 2279 2828 2325
rect 3002 2279 3015 2325
rect 2815 2236 3015 2279
rect 2815 1993 3015 2036
rect 2815 1947 2828 1993
rect 3002 1947 3015 1993
rect 2815 1934 3015 1947
rect 3095 2325 3295 2338
rect 3095 2279 3108 2325
rect 3282 2279 3295 2325
rect 3095 2236 3295 2279
rect 3095 1993 3295 2036
rect 3095 1947 3108 1993
rect 3282 1947 3295 1993
rect 3095 1934 3295 1947
rect 3375 2325 3575 2338
rect 3375 2279 3388 2325
rect 3562 2279 3575 2325
rect 3375 2236 3575 2279
rect 3375 1993 3575 2036
rect 3375 1947 3388 1993
rect 3562 1947 3575 1993
rect 3375 1934 3575 1947
rect 3655 2325 3855 2338
rect 3655 2279 3668 2325
rect 3842 2279 3855 2325
rect 3655 2236 3855 2279
rect 3655 1993 3855 2036
rect 3655 1947 3668 1993
rect 3842 1947 3855 1993
rect 3655 1934 3855 1947
rect 3935 2325 4135 2338
rect 3935 2279 3948 2325
rect 4122 2279 4135 2325
rect 3935 2236 4135 2279
rect 3935 1993 4135 2036
rect 3935 1947 3948 1993
rect 4122 1947 4135 1993
rect 3935 1934 4135 1947
rect 4215 2325 4415 2338
rect 4215 2279 4228 2325
rect 4402 2279 4415 2325
rect 4215 2236 4415 2279
rect 4215 1993 4415 2036
rect 4215 1947 4228 1993
rect 4402 1947 4415 1993
rect 4215 1934 4415 1947
rect 4495 2325 4695 2338
rect 4495 2279 4508 2325
rect 4682 2279 4695 2325
rect 4495 2236 4695 2279
rect 4495 1993 4695 2036
rect 4495 1947 4508 1993
rect 4682 1947 4695 1993
rect 4495 1934 4695 1947
rect 4775 2325 4975 2338
rect 4775 2279 4788 2325
rect 4962 2279 4975 2325
rect 4775 2236 4975 2279
rect 4775 1993 4975 2036
rect 4775 1947 4788 1993
rect 4962 1947 4975 1993
rect 4775 1934 4975 1947
rect 5055 2325 5255 2338
rect 5055 2279 5068 2325
rect 5242 2279 5255 2325
rect 5055 2236 5255 2279
rect 5055 1993 5255 2036
rect 5055 1947 5068 1993
rect 5242 1947 5255 1993
rect 5055 1934 5255 1947
rect 5335 2325 5535 2338
rect 5335 2279 5348 2325
rect 5522 2279 5535 2325
rect 5335 2236 5535 2279
rect 5335 1993 5535 2036
rect 5335 1947 5348 1993
rect 5522 1947 5535 1993
rect 5335 1934 5535 1947
rect 5615 2325 5815 2338
rect 5615 2279 5628 2325
rect 5802 2279 5815 2325
rect 5615 2236 5815 2279
rect 5615 1993 5815 2036
rect 5615 1947 5628 1993
rect 5802 1947 5815 1993
rect 5615 1934 5815 1947
rect 5895 2325 6095 2338
rect 5895 2279 5908 2325
rect 6082 2279 6095 2325
rect 5895 2236 6095 2279
rect 5895 1993 6095 2036
rect 5895 1947 5908 1993
rect 6082 1947 6095 1993
rect 5895 1934 6095 1947
rect 6175 2325 6375 2338
rect 6175 2279 6188 2325
rect 6362 2279 6375 2325
rect 6175 2236 6375 2279
rect 6175 1993 6375 2036
rect 6175 1947 6188 1993
rect 6362 1947 6375 1993
rect 6175 1934 6375 1947
rect 6455 2325 6655 2338
rect 6455 2279 6468 2325
rect 6642 2279 6655 2325
rect 6455 2236 6655 2279
rect 6455 1993 6655 2036
rect 6455 1947 6468 1993
rect 6642 1947 6655 1993
rect 6455 1934 6655 1947
rect 6735 2325 6935 2338
rect 6735 2279 6748 2325
rect 6922 2279 6935 2325
rect 6735 2236 6935 2279
rect 6735 1993 6935 2036
rect 6735 1947 6748 1993
rect 6922 1947 6935 1993
rect 6735 1934 6935 1947
rect 7015 2325 7215 2338
rect 7015 2279 7028 2325
rect 7202 2279 7215 2325
rect 7015 2236 7215 2279
rect 7015 1993 7215 2036
rect 7015 1947 7028 1993
rect 7202 1947 7215 1993
rect 7015 1934 7215 1947
rect 7295 2325 7495 2338
rect 7295 2279 7308 2325
rect 7482 2279 7495 2325
rect 7295 2236 7495 2279
rect 7295 1993 7495 2036
rect 7295 1947 7308 1993
rect 7482 1947 7495 1993
rect 7295 1934 7495 1947
rect 7575 2325 7775 2338
rect 7575 2279 7588 2325
rect 7762 2279 7775 2325
rect 7575 2236 7775 2279
rect 7575 1993 7775 2036
rect 7575 1947 7588 1993
rect 7762 1947 7775 1993
rect 7575 1934 7775 1947
rect 7855 2325 8055 2338
rect 7855 2279 7868 2325
rect 8042 2279 8055 2325
rect 7855 2236 8055 2279
rect 7855 1993 8055 2036
rect 7855 1947 7868 1993
rect 8042 1947 8055 1993
rect 7855 1934 8055 1947
rect 8135 2325 8335 2338
rect 8135 2279 8148 2325
rect 8322 2279 8335 2325
rect 8135 2236 8335 2279
rect 8135 1993 8335 2036
rect 8135 1947 8148 1993
rect 8322 1947 8335 1993
rect 8135 1934 8335 1947
rect 8415 2325 8615 2338
rect 8415 2279 8428 2325
rect 8602 2279 8615 2325
rect 8415 2236 8615 2279
rect 8415 1993 8615 2036
rect 8415 1947 8428 1993
rect 8602 1947 8615 1993
rect 8415 1934 8615 1947
rect 8695 2325 8895 2338
rect 8695 2279 8708 2325
rect 8882 2279 8895 2325
rect 8695 2236 8895 2279
rect 8695 1993 8895 2036
rect 8695 1947 8708 1993
rect 8882 1947 8895 1993
rect 8695 1934 8895 1947
rect 8975 2325 9175 2338
rect 8975 2279 8988 2325
rect 9162 2279 9175 2325
rect 8975 2236 9175 2279
rect 8975 1993 9175 2036
rect 8975 1947 8988 1993
rect 9162 1947 9175 1993
rect 8975 1934 9175 1947
rect 9255 2325 9455 2338
rect 9255 2279 9268 2325
rect 9442 2279 9455 2325
rect 9255 2236 9455 2279
rect 9255 1993 9455 2036
rect 9255 1947 9268 1993
rect 9442 1947 9455 1993
rect 9255 1934 9455 1947
rect 9535 2325 9735 2338
rect 9535 2279 9548 2325
rect 9722 2279 9735 2325
rect 9535 2236 9735 2279
rect 9535 1993 9735 2036
rect 9535 1947 9548 1993
rect 9722 1947 9735 1993
rect 9535 1934 9735 1947
rect 295 1673 495 1686
rect 295 1627 308 1673
rect 482 1627 495 1673
rect 295 1584 495 1627
rect 295 1341 495 1384
rect 295 1295 308 1341
rect 482 1295 495 1341
rect 295 1282 495 1295
rect 575 1673 775 1686
rect 575 1627 588 1673
rect 762 1627 775 1673
rect 575 1584 775 1627
rect 575 1341 775 1384
rect 575 1295 588 1341
rect 762 1295 775 1341
rect 575 1282 775 1295
rect 855 1673 1055 1686
rect 855 1627 868 1673
rect 1042 1627 1055 1673
rect 855 1584 1055 1627
rect 855 1341 1055 1384
rect 855 1295 868 1341
rect 1042 1295 1055 1341
rect 855 1282 1055 1295
rect 1135 1673 1335 1686
rect 1135 1627 1148 1673
rect 1322 1627 1335 1673
rect 1135 1584 1335 1627
rect 1135 1341 1335 1384
rect 1135 1295 1148 1341
rect 1322 1295 1335 1341
rect 1135 1282 1335 1295
rect 1415 1673 1615 1686
rect 1415 1627 1428 1673
rect 1602 1627 1615 1673
rect 1415 1584 1615 1627
rect 1415 1341 1615 1384
rect 1415 1295 1428 1341
rect 1602 1295 1615 1341
rect 1415 1282 1615 1295
rect 1695 1673 1895 1686
rect 1695 1627 1708 1673
rect 1882 1627 1895 1673
rect 1695 1584 1895 1627
rect 1695 1341 1895 1384
rect 1695 1295 1708 1341
rect 1882 1295 1895 1341
rect 1695 1282 1895 1295
rect 1975 1673 2175 1686
rect 1975 1627 1988 1673
rect 2162 1627 2175 1673
rect 1975 1584 2175 1627
rect 1975 1341 2175 1384
rect 1975 1295 1988 1341
rect 2162 1295 2175 1341
rect 1975 1282 2175 1295
rect 2255 1673 2455 1686
rect 2255 1627 2268 1673
rect 2442 1627 2455 1673
rect 2255 1584 2455 1627
rect 2255 1341 2455 1384
rect 2255 1295 2268 1341
rect 2442 1295 2455 1341
rect 2255 1282 2455 1295
rect 2535 1673 2735 1686
rect 2535 1627 2548 1673
rect 2722 1627 2735 1673
rect 2535 1584 2735 1627
rect 2535 1341 2735 1384
rect 2535 1295 2548 1341
rect 2722 1295 2735 1341
rect 2535 1282 2735 1295
rect 2815 1673 3015 1686
rect 2815 1627 2828 1673
rect 3002 1627 3015 1673
rect 2815 1584 3015 1627
rect 2815 1341 3015 1384
rect 2815 1295 2828 1341
rect 3002 1295 3015 1341
rect 2815 1282 3015 1295
rect 3095 1673 3295 1686
rect 3095 1627 3108 1673
rect 3282 1627 3295 1673
rect 3095 1584 3295 1627
rect 3095 1341 3295 1384
rect 3095 1295 3108 1341
rect 3282 1295 3295 1341
rect 3095 1282 3295 1295
rect 3375 1673 3575 1686
rect 3375 1627 3388 1673
rect 3562 1627 3575 1673
rect 3375 1584 3575 1627
rect 3375 1341 3575 1384
rect 3375 1295 3388 1341
rect 3562 1295 3575 1341
rect 3375 1282 3575 1295
rect 3655 1673 3855 1686
rect 3655 1627 3668 1673
rect 3842 1627 3855 1673
rect 3655 1584 3855 1627
rect 3655 1341 3855 1384
rect 3655 1295 3668 1341
rect 3842 1295 3855 1341
rect 3655 1282 3855 1295
rect 3935 1673 4135 1686
rect 3935 1627 3948 1673
rect 4122 1627 4135 1673
rect 3935 1584 4135 1627
rect 3935 1341 4135 1384
rect 3935 1295 3948 1341
rect 4122 1295 4135 1341
rect 3935 1282 4135 1295
rect 4215 1673 4415 1686
rect 4215 1627 4228 1673
rect 4402 1627 4415 1673
rect 4215 1584 4415 1627
rect 4215 1341 4415 1384
rect 4215 1295 4228 1341
rect 4402 1295 4415 1341
rect 4215 1282 4415 1295
rect 4495 1673 4695 1686
rect 4495 1627 4508 1673
rect 4682 1627 4695 1673
rect 4495 1584 4695 1627
rect 4495 1341 4695 1384
rect 4495 1295 4508 1341
rect 4682 1295 4695 1341
rect 4495 1282 4695 1295
rect 4775 1673 4975 1686
rect 4775 1627 4788 1673
rect 4962 1627 4975 1673
rect 4775 1584 4975 1627
rect 4775 1341 4975 1384
rect 4775 1295 4788 1341
rect 4962 1295 4975 1341
rect 4775 1282 4975 1295
rect 5055 1673 5255 1686
rect 5055 1627 5068 1673
rect 5242 1627 5255 1673
rect 5055 1584 5255 1627
rect 5055 1341 5255 1384
rect 5055 1295 5068 1341
rect 5242 1295 5255 1341
rect 5055 1282 5255 1295
rect 5335 1673 5535 1686
rect 5335 1627 5348 1673
rect 5522 1627 5535 1673
rect 5335 1584 5535 1627
rect 5335 1341 5535 1384
rect 5335 1295 5348 1341
rect 5522 1295 5535 1341
rect 5335 1282 5535 1295
rect 5615 1673 5815 1686
rect 5615 1627 5628 1673
rect 5802 1627 5815 1673
rect 5615 1584 5815 1627
rect 5615 1341 5815 1384
rect 5615 1295 5628 1341
rect 5802 1295 5815 1341
rect 5615 1282 5815 1295
rect 5895 1673 6095 1686
rect 5895 1627 5908 1673
rect 6082 1627 6095 1673
rect 5895 1584 6095 1627
rect 5895 1341 6095 1384
rect 5895 1295 5908 1341
rect 6082 1295 6095 1341
rect 5895 1282 6095 1295
rect 6175 1673 6375 1686
rect 6175 1627 6188 1673
rect 6362 1627 6375 1673
rect 6175 1584 6375 1627
rect 6175 1341 6375 1384
rect 6175 1295 6188 1341
rect 6362 1295 6375 1341
rect 6175 1282 6375 1295
rect 6455 1673 6655 1686
rect 6455 1627 6468 1673
rect 6642 1627 6655 1673
rect 6455 1584 6655 1627
rect 6455 1341 6655 1384
rect 6455 1295 6468 1341
rect 6642 1295 6655 1341
rect 6455 1282 6655 1295
rect 6735 1673 6935 1686
rect 6735 1627 6748 1673
rect 6922 1627 6935 1673
rect 6735 1584 6935 1627
rect 6735 1341 6935 1384
rect 6735 1295 6748 1341
rect 6922 1295 6935 1341
rect 6735 1282 6935 1295
rect 7015 1673 7215 1686
rect 7015 1627 7028 1673
rect 7202 1627 7215 1673
rect 7015 1584 7215 1627
rect 7015 1341 7215 1384
rect 7015 1295 7028 1341
rect 7202 1295 7215 1341
rect 7015 1282 7215 1295
rect 7295 1673 7495 1686
rect 7295 1627 7308 1673
rect 7482 1627 7495 1673
rect 7295 1584 7495 1627
rect 7295 1341 7495 1384
rect 7295 1295 7308 1341
rect 7482 1295 7495 1341
rect 7295 1282 7495 1295
rect 7575 1673 7775 1686
rect 7575 1627 7588 1673
rect 7762 1627 7775 1673
rect 7575 1584 7775 1627
rect 7575 1341 7775 1384
rect 7575 1295 7588 1341
rect 7762 1295 7775 1341
rect 7575 1282 7775 1295
rect 7855 1673 8055 1686
rect 7855 1627 7868 1673
rect 8042 1627 8055 1673
rect 7855 1584 8055 1627
rect 7855 1341 8055 1384
rect 7855 1295 7868 1341
rect 8042 1295 8055 1341
rect 7855 1282 8055 1295
rect 8135 1673 8335 1686
rect 8135 1627 8148 1673
rect 8322 1627 8335 1673
rect 8135 1584 8335 1627
rect 8135 1341 8335 1384
rect 8135 1295 8148 1341
rect 8322 1295 8335 1341
rect 8135 1282 8335 1295
rect 8415 1673 8615 1686
rect 8415 1627 8428 1673
rect 8602 1627 8615 1673
rect 8415 1584 8615 1627
rect 8415 1341 8615 1384
rect 8415 1295 8428 1341
rect 8602 1295 8615 1341
rect 8415 1282 8615 1295
rect 8695 1673 8895 1686
rect 8695 1627 8708 1673
rect 8882 1627 8895 1673
rect 8695 1584 8895 1627
rect 8695 1341 8895 1384
rect 8695 1295 8708 1341
rect 8882 1295 8895 1341
rect 8695 1282 8895 1295
rect 8975 1673 9175 1686
rect 8975 1627 8988 1673
rect 9162 1627 9175 1673
rect 8975 1584 9175 1627
rect 8975 1341 9175 1384
rect 8975 1295 8988 1341
rect 9162 1295 9175 1341
rect 8975 1282 9175 1295
rect 9255 1673 9455 1686
rect 9255 1627 9268 1673
rect 9442 1627 9455 1673
rect 9255 1584 9455 1627
rect 9255 1341 9455 1384
rect 9255 1295 9268 1341
rect 9442 1295 9455 1341
rect 9255 1282 9455 1295
rect 9535 1673 9735 1686
rect 9535 1627 9548 1673
rect 9722 1627 9735 1673
rect 9535 1584 9735 1627
rect 9535 1341 9735 1384
rect 9535 1295 9548 1341
rect 9722 1295 9735 1341
rect 9535 1282 9735 1295
<< polycontact >>
rect 308 5360 482 5406
rect 308 5028 482 5074
rect 588 5360 762 5406
rect 588 5028 762 5074
rect 868 5360 1042 5406
rect 868 5028 1042 5074
rect 1148 5360 1322 5406
rect 1148 5028 1322 5074
rect 1428 5360 1602 5406
rect 1428 5028 1602 5074
rect 1708 5360 1882 5406
rect 1708 5028 1882 5074
rect 1988 5360 2162 5406
rect 1988 5028 2162 5074
rect 2268 5360 2442 5406
rect 2268 5028 2442 5074
rect 2548 5360 2722 5406
rect 2548 5028 2722 5074
rect 2828 5360 3002 5406
rect 2828 5028 3002 5074
rect 3108 5360 3282 5406
rect 3108 5028 3282 5074
rect 3388 5360 3562 5406
rect 3388 5028 3562 5074
rect 3668 5360 3842 5406
rect 3668 5028 3842 5074
rect 3948 5360 4122 5406
rect 3948 5028 4122 5074
rect 4228 5360 4402 5406
rect 4228 5028 4402 5074
rect 4508 5360 4682 5406
rect 4508 5028 4682 5074
rect 4788 5360 4962 5406
rect 4788 5028 4962 5074
rect 5068 5360 5242 5406
rect 5068 5028 5242 5074
rect 5348 5360 5522 5406
rect 5348 5028 5522 5074
rect 5628 5360 5802 5406
rect 5628 5028 5802 5074
rect 5908 5360 6082 5406
rect 5908 5028 6082 5074
rect 6188 5360 6362 5406
rect 6188 5028 6362 5074
rect 6468 5360 6642 5406
rect 6468 5028 6642 5074
rect 6748 5360 6922 5406
rect 6748 5028 6922 5074
rect 7028 5360 7202 5406
rect 7028 5028 7202 5074
rect 7308 5360 7482 5406
rect 7308 5028 7482 5074
rect 7588 5360 7762 5406
rect 7588 5028 7762 5074
rect 7868 5360 8042 5406
rect 7868 5028 8042 5074
rect 8148 5360 8322 5406
rect 8148 5028 8322 5074
rect 8428 5360 8602 5406
rect 8428 5028 8602 5074
rect 8708 5360 8882 5406
rect 8708 5028 8882 5074
rect 8988 5360 9162 5406
rect 8988 5028 9162 5074
rect 9268 5360 9442 5406
rect 9268 5028 9442 5074
rect 9548 5360 9722 5406
rect 9548 5028 9722 5074
rect 308 4708 482 4754
rect 308 4376 482 4422
rect 588 4708 762 4754
rect 588 4376 762 4422
rect 868 4708 1042 4754
rect 868 4376 1042 4422
rect 1148 4708 1322 4754
rect 1148 4376 1322 4422
rect 1428 4708 1602 4754
rect 1428 4376 1602 4422
rect 1708 4708 1882 4754
rect 1708 4376 1882 4422
rect 1988 4708 2162 4754
rect 1988 4376 2162 4422
rect 2268 4708 2442 4754
rect 2268 4376 2442 4422
rect 2548 4708 2722 4754
rect 2548 4376 2722 4422
rect 2828 4708 3002 4754
rect 2828 4376 3002 4422
rect 3108 4708 3282 4754
rect 3108 4376 3282 4422
rect 3388 4708 3562 4754
rect 3388 4376 3562 4422
rect 3668 4708 3842 4754
rect 3668 4376 3842 4422
rect 3948 4708 4122 4754
rect 3948 4376 4122 4422
rect 4228 4708 4402 4754
rect 4228 4376 4402 4422
rect 4508 4708 4682 4754
rect 4508 4376 4682 4422
rect 4788 4708 4962 4754
rect 4788 4376 4962 4422
rect 5068 4708 5242 4754
rect 5068 4376 5242 4422
rect 5348 4708 5522 4754
rect 5348 4376 5522 4422
rect 5628 4708 5802 4754
rect 5628 4376 5802 4422
rect 5908 4708 6082 4754
rect 5908 4376 6082 4422
rect 6188 4708 6362 4754
rect 6188 4376 6362 4422
rect 6468 4708 6642 4754
rect 6468 4376 6642 4422
rect 6748 4708 6922 4754
rect 6748 4376 6922 4422
rect 7028 4708 7202 4754
rect 7028 4376 7202 4422
rect 7308 4708 7482 4754
rect 7308 4376 7482 4422
rect 7588 4708 7762 4754
rect 7588 4376 7762 4422
rect 7868 4708 8042 4754
rect 7868 4376 8042 4422
rect 8148 4708 8322 4754
rect 8148 4376 8322 4422
rect 8428 4708 8602 4754
rect 8428 4376 8602 4422
rect 8708 4708 8882 4754
rect 8708 4376 8882 4422
rect 8988 4708 9162 4754
rect 8988 4376 9162 4422
rect 9268 4708 9442 4754
rect 9268 4376 9442 4422
rect 9548 4708 9722 4754
rect 9548 4376 9722 4422
rect 308 4056 482 4102
rect 308 3724 482 3770
rect 588 4056 762 4102
rect 588 3724 762 3770
rect 868 4056 1042 4102
rect 868 3724 1042 3770
rect 1148 4056 1322 4102
rect 1148 3724 1322 3770
rect 1428 4056 1602 4102
rect 1428 3724 1602 3770
rect 1708 4056 1882 4102
rect 1708 3724 1882 3770
rect 1988 4056 2162 4102
rect 1988 3724 2162 3770
rect 2268 4056 2442 4102
rect 2268 3724 2442 3770
rect 2548 4056 2722 4102
rect 2548 3724 2722 3770
rect 2828 4056 3002 4102
rect 2828 3724 3002 3770
rect 3108 4056 3282 4102
rect 3108 3724 3282 3770
rect 3388 4056 3562 4102
rect 3388 3724 3562 3770
rect 3668 4056 3842 4102
rect 3668 3724 3842 3770
rect 3948 4056 4122 4102
rect 3948 3724 4122 3770
rect 4228 4056 4402 4102
rect 4228 3724 4402 3770
rect 4508 4056 4682 4102
rect 4508 3724 4682 3770
rect 4788 4056 4962 4102
rect 4788 3724 4962 3770
rect 5068 4056 5242 4102
rect 5068 3724 5242 3770
rect 5348 4056 5522 4102
rect 5348 3724 5522 3770
rect 5628 4056 5802 4102
rect 5628 3724 5802 3770
rect 5908 4056 6082 4102
rect 5908 3724 6082 3770
rect 6188 4056 6362 4102
rect 6188 3724 6362 3770
rect 6468 4056 6642 4102
rect 6468 3724 6642 3770
rect 6748 4056 6922 4102
rect 6748 3724 6922 3770
rect 7028 4056 7202 4102
rect 7028 3724 7202 3770
rect 7308 4056 7482 4102
rect 7308 3724 7482 3770
rect 7588 4056 7762 4102
rect 7588 3724 7762 3770
rect 7868 4056 8042 4102
rect 7868 3724 8042 3770
rect 8148 4056 8322 4102
rect 8148 3724 8322 3770
rect 8428 4056 8602 4102
rect 8428 3724 8602 3770
rect 8708 4056 8882 4102
rect 8708 3724 8882 3770
rect 8988 4056 9162 4102
rect 8988 3724 9162 3770
rect 9268 4056 9442 4102
rect 9268 3724 9442 3770
rect 9548 4056 9722 4102
rect 9548 3724 9722 3770
rect 308 2931 482 2977
rect 308 2599 482 2645
rect 588 2931 762 2977
rect 588 2599 762 2645
rect 868 2931 1042 2977
rect 868 2599 1042 2645
rect 1148 2931 1322 2977
rect 1148 2599 1322 2645
rect 1428 2931 1602 2977
rect 1428 2599 1602 2645
rect 1708 2931 1882 2977
rect 1708 2599 1882 2645
rect 1988 2931 2162 2977
rect 1988 2599 2162 2645
rect 2268 2931 2442 2977
rect 2268 2599 2442 2645
rect 2548 2931 2722 2977
rect 2548 2599 2722 2645
rect 2828 2931 3002 2977
rect 2828 2599 3002 2645
rect 3108 2931 3282 2977
rect 3108 2599 3282 2645
rect 3388 2931 3562 2977
rect 3388 2599 3562 2645
rect 3668 2931 3842 2977
rect 3668 2599 3842 2645
rect 3948 2931 4122 2977
rect 3948 2599 4122 2645
rect 4228 2931 4402 2977
rect 4228 2599 4402 2645
rect 4508 2931 4682 2977
rect 4508 2599 4682 2645
rect 4788 2931 4962 2977
rect 4788 2599 4962 2645
rect 5068 2931 5242 2977
rect 5068 2599 5242 2645
rect 5348 2931 5522 2977
rect 5348 2599 5522 2645
rect 5628 2931 5802 2977
rect 5628 2599 5802 2645
rect 5908 2931 6082 2977
rect 5908 2599 6082 2645
rect 6188 2931 6362 2977
rect 6188 2599 6362 2645
rect 6468 2931 6642 2977
rect 6468 2599 6642 2645
rect 6748 2931 6922 2977
rect 6748 2599 6922 2645
rect 7028 2931 7202 2977
rect 7028 2599 7202 2645
rect 7308 2931 7482 2977
rect 7308 2599 7482 2645
rect 7588 2931 7762 2977
rect 7588 2599 7762 2645
rect 7868 2931 8042 2977
rect 7868 2599 8042 2645
rect 8148 2931 8322 2977
rect 8148 2599 8322 2645
rect 8428 2931 8602 2977
rect 8428 2599 8602 2645
rect 8708 2931 8882 2977
rect 8708 2599 8882 2645
rect 8988 2931 9162 2977
rect 8988 2599 9162 2645
rect 9268 2931 9442 2977
rect 9268 2599 9442 2645
rect 9548 2931 9722 2977
rect 9548 2599 9722 2645
rect 308 2279 482 2325
rect 308 1947 482 1993
rect 588 2279 762 2325
rect 588 1947 762 1993
rect 868 2279 1042 2325
rect 868 1947 1042 1993
rect 1148 2279 1322 2325
rect 1148 1947 1322 1993
rect 1428 2279 1602 2325
rect 1428 1947 1602 1993
rect 1708 2279 1882 2325
rect 1708 1947 1882 1993
rect 1988 2279 2162 2325
rect 1988 1947 2162 1993
rect 2268 2279 2442 2325
rect 2268 1947 2442 1993
rect 2548 2279 2722 2325
rect 2548 1947 2722 1993
rect 2828 2279 3002 2325
rect 2828 1947 3002 1993
rect 3108 2279 3282 2325
rect 3108 1947 3282 1993
rect 3388 2279 3562 2325
rect 3388 1947 3562 1993
rect 3668 2279 3842 2325
rect 3668 1947 3842 1993
rect 3948 2279 4122 2325
rect 3948 1947 4122 1993
rect 4228 2279 4402 2325
rect 4228 1947 4402 1993
rect 4508 2279 4682 2325
rect 4508 1947 4682 1993
rect 4788 2279 4962 2325
rect 4788 1947 4962 1993
rect 5068 2279 5242 2325
rect 5068 1947 5242 1993
rect 5348 2279 5522 2325
rect 5348 1947 5522 1993
rect 5628 2279 5802 2325
rect 5628 1947 5802 1993
rect 5908 2279 6082 2325
rect 5908 1947 6082 1993
rect 6188 2279 6362 2325
rect 6188 1947 6362 1993
rect 6468 2279 6642 2325
rect 6468 1947 6642 1993
rect 6748 2279 6922 2325
rect 6748 1947 6922 1993
rect 7028 2279 7202 2325
rect 7028 1947 7202 1993
rect 7308 2279 7482 2325
rect 7308 1947 7482 1993
rect 7588 2279 7762 2325
rect 7588 1947 7762 1993
rect 7868 2279 8042 2325
rect 7868 1947 8042 1993
rect 8148 2279 8322 2325
rect 8148 1947 8322 1993
rect 8428 2279 8602 2325
rect 8428 1947 8602 1993
rect 8708 2279 8882 2325
rect 8708 1947 8882 1993
rect 8988 2279 9162 2325
rect 8988 1947 9162 1993
rect 9268 2279 9442 2325
rect 9268 1947 9442 1993
rect 9548 2279 9722 2325
rect 9548 1947 9722 1993
rect 308 1627 482 1673
rect 308 1295 482 1341
rect 588 1627 762 1673
rect 588 1295 762 1341
rect 868 1627 1042 1673
rect 868 1295 1042 1341
rect 1148 1627 1322 1673
rect 1148 1295 1322 1341
rect 1428 1627 1602 1673
rect 1428 1295 1602 1341
rect 1708 1627 1882 1673
rect 1708 1295 1882 1341
rect 1988 1627 2162 1673
rect 1988 1295 2162 1341
rect 2268 1627 2442 1673
rect 2268 1295 2442 1341
rect 2548 1627 2722 1673
rect 2548 1295 2722 1341
rect 2828 1627 3002 1673
rect 2828 1295 3002 1341
rect 3108 1627 3282 1673
rect 3108 1295 3282 1341
rect 3388 1627 3562 1673
rect 3388 1295 3562 1341
rect 3668 1627 3842 1673
rect 3668 1295 3842 1341
rect 3948 1627 4122 1673
rect 3948 1295 4122 1341
rect 4228 1627 4402 1673
rect 4228 1295 4402 1341
rect 4508 1627 4682 1673
rect 4508 1295 4682 1341
rect 4788 1627 4962 1673
rect 4788 1295 4962 1341
rect 5068 1627 5242 1673
rect 5068 1295 5242 1341
rect 5348 1627 5522 1673
rect 5348 1295 5522 1341
rect 5628 1627 5802 1673
rect 5628 1295 5802 1341
rect 5908 1627 6082 1673
rect 5908 1295 6082 1341
rect 6188 1627 6362 1673
rect 6188 1295 6362 1341
rect 6468 1627 6642 1673
rect 6468 1295 6642 1341
rect 6748 1627 6922 1673
rect 6748 1295 6922 1341
rect 7028 1627 7202 1673
rect 7028 1295 7202 1341
rect 7308 1627 7482 1673
rect 7308 1295 7482 1341
rect 7588 1627 7762 1673
rect 7588 1295 7762 1341
rect 7868 1627 8042 1673
rect 7868 1295 8042 1341
rect 8148 1627 8322 1673
rect 8148 1295 8322 1341
rect 8428 1627 8602 1673
rect 8428 1295 8602 1341
rect 8708 1627 8882 1673
rect 8708 1295 8882 1341
rect 8988 1627 9162 1673
rect 8988 1295 9162 1341
rect 9268 1627 9442 1673
rect 9268 1295 9442 1341
rect 9548 1627 9722 1673
rect 9548 1295 9722 1341
<< ppolyres >>
rect 295 5117 495 5317
rect 575 5117 775 5317
rect 855 5117 1055 5317
rect 1135 5117 1335 5317
rect 1415 5117 1615 5317
rect 1695 5117 1895 5317
rect 1975 5117 2175 5317
rect 2255 5117 2455 5317
rect 2535 5117 2735 5317
rect 2815 5117 3015 5317
rect 3095 5117 3295 5317
rect 3375 5117 3575 5317
rect 3655 5117 3855 5317
rect 3935 5117 4135 5317
rect 4215 5117 4415 5317
rect 4495 5117 4695 5317
rect 4775 5117 4975 5317
rect 5055 5117 5255 5317
rect 5335 5117 5535 5317
rect 5615 5117 5815 5317
rect 5895 5117 6095 5317
rect 6175 5117 6375 5317
rect 6455 5117 6655 5317
rect 6735 5117 6935 5317
rect 7015 5117 7215 5317
rect 7295 5117 7495 5317
rect 7575 5117 7775 5317
rect 7855 5117 8055 5317
rect 8135 5117 8335 5317
rect 8415 5117 8615 5317
rect 8695 5117 8895 5317
rect 8975 5117 9175 5317
rect 9255 5117 9455 5317
rect 9535 5117 9735 5317
rect 295 4465 495 4665
rect 575 4465 775 4665
rect 855 4465 1055 4665
rect 1135 4465 1335 4665
rect 1415 4465 1615 4665
rect 1695 4465 1895 4665
rect 1975 4465 2175 4665
rect 2255 4465 2455 4665
rect 2535 4465 2735 4665
rect 2815 4465 3015 4665
rect 3095 4465 3295 4665
rect 3375 4465 3575 4665
rect 3655 4465 3855 4665
rect 3935 4465 4135 4665
rect 4215 4465 4415 4665
rect 4495 4465 4695 4665
rect 4775 4465 4975 4665
rect 5055 4465 5255 4665
rect 5335 4465 5535 4665
rect 5615 4465 5815 4665
rect 5895 4465 6095 4665
rect 6175 4465 6375 4665
rect 6455 4465 6655 4665
rect 6735 4465 6935 4665
rect 7015 4465 7215 4665
rect 7295 4465 7495 4665
rect 7575 4465 7775 4665
rect 7855 4465 8055 4665
rect 8135 4465 8335 4665
rect 8415 4465 8615 4665
rect 8695 4465 8895 4665
rect 8975 4465 9175 4665
rect 9255 4465 9455 4665
rect 9535 4465 9735 4665
rect 295 3813 495 4013
rect 575 3813 775 4013
rect 855 3813 1055 4013
rect 1135 3813 1335 4013
rect 1415 3813 1615 4013
rect 1695 3813 1895 4013
rect 1975 3813 2175 4013
rect 2255 3813 2455 4013
rect 2535 3813 2735 4013
rect 2815 3813 3015 4013
rect 3095 3813 3295 4013
rect 3375 3813 3575 4013
rect 3655 3813 3855 4013
rect 3935 3813 4135 4013
rect 4215 3813 4415 4013
rect 4495 3813 4695 4013
rect 4775 3813 4975 4013
rect 5055 3813 5255 4013
rect 5335 3813 5535 4013
rect 5615 3813 5815 4013
rect 5895 3813 6095 4013
rect 6175 3813 6375 4013
rect 6455 3813 6655 4013
rect 6735 3813 6935 4013
rect 7015 3813 7215 4013
rect 7295 3813 7495 4013
rect 7575 3813 7775 4013
rect 7855 3813 8055 4013
rect 8135 3813 8335 4013
rect 8415 3813 8615 4013
rect 8695 3813 8895 4013
rect 8975 3813 9175 4013
rect 9255 3813 9455 4013
rect 9535 3813 9735 4013
rect 295 2688 495 2888
rect 575 2688 775 2888
rect 855 2688 1055 2888
rect 1135 2688 1335 2888
rect 1415 2688 1615 2888
rect 1695 2688 1895 2888
rect 1975 2688 2175 2888
rect 2255 2688 2455 2888
rect 2535 2688 2735 2888
rect 2815 2688 3015 2888
rect 3095 2688 3295 2888
rect 3375 2688 3575 2888
rect 3655 2688 3855 2888
rect 3935 2688 4135 2888
rect 4215 2688 4415 2888
rect 4495 2688 4695 2888
rect 4775 2688 4975 2888
rect 5055 2688 5255 2888
rect 5335 2688 5535 2888
rect 5615 2688 5815 2888
rect 5895 2688 6095 2888
rect 6175 2688 6375 2888
rect 6455 2688 6655 2888
rect 6735 2688 6935 2888
rect 7015 2688 7215 2888
rect 7295 2688 7495 2888
rect 7575 2688 7775 2888
rect 7855 2688 8055 2888
rect 8135 2688 8335 2888
rect 8415 2688 8615 2888
rect 8695 2688 8895 2888
rect 8975 2688 9175 2888
rect 9255 2688 9455 2888
rect 9535 2688 9735 2888
rect 295 2036 495 2236
rect 575 2036 775 2236
rect 855 2036 1055 2236
rect 1135 2036 1335 2236
rect 1415 2036 1615 2236
rect 1695 2036 1895 2236
rect 1975 2036 2175 2236
rect 2255 2036 2455 2236
rect 2535 2036 2735 2236
rect 2815 2036 3015 2236
rect 3095 2036 3295 2236
rect 3375 2036 3575 2236
rect 3655 2036 3855 2236
rect 3935 2036 4135 2236
rect 4215 2036 4415 2236
rect 4495 2036 4695 2236
rect 4775 2036 4975 2236
rect 5055 2036 5255 2236
rect 5335 2036 5535 2236
rect 5615 2036 5815 2236
rect 5895 2036 6095 2236
rect 6175 2036 6375 2236
rect 6455 2036 6655 2236
rect 6735 2036 6935 2236
rect 7015 2036 7215 2236
rect 7295 2036 7495 2236
rect 7575 2036 7775 2236
rect 7855 2036 8055 2236
rect 8135 2036 8335 2236
rect 8415 2036 8615 2236
rect 8695 2036 8895 2236
rect 8975 2036 9175 2236
rect 9255 2036 9455 2236
rect 9535 2036 9735 2236
rect 295 1384 495 1584
rect 575 1384 775 1584
rect 855 1384 1055 1584
rect 1135 1384 1335 1584
rect 1415 1384 1615 1584
rect 1695 1384 1895 1584
rect 1975 1384 2175 1584
rect 2255 1384 2455 1584
rect 2535 1384 2735 1584
rect 2815 1384 3015 1584
rect 3095 1384 3295 1584
rect 3375 1384 3575 1584
rect 3655 1384 3855 1584
rect 3935 1384 4135 1584
rect 4215 1384 4415 1584
rect 4495 1384 4695 1584
rect 4775 1384 4975 1584
rect 5055 1384 5255 1584
rect 5335 1384 5535 1584
rect 5615 1384 5815 1584
rect 5895 1384 6095 1584
rect 6175 1384 6375 1584
rect 6455 1384 6655 1584
rect 6735 1384 6935 1584
rect 7015 1384 7215 1584
rect 7295 1384 7495 1584
rect 7575 1384 7775 1584
rect 7855 1384 8055 1584
rect 8135 1384 8335 1584
rect 8415 1384 8615 1584
rect 8695 1384 8895 1584
rect 8975 1384 9175 1584
rect 9255 1384 9455 1584
rect 9535 1384 9735 1584
<< metal1 >>
rect -39 5698 10069 5715
rect -39 5648 -22 5698
rect 24 5652 76 5698
rect 122 5652 174 5698
rect 220 5652 272 5698
rect 318 5652 370 5698
rect 416 5652 468 5698
rect 514 5652 566 5698
rect 612 5652 664 5698
rect 710 5652 762 5698
rect 808 5652 860 5698
rect 906 5652 958 5698
rect 1004 5652 1056 5698
rect 1102 5652 1154 5698
rect 1200 5652 1252 5698
rect 1298 5652 1350 5698
rect 1396 5652 1448 5698
rect 1494 5652 1546 5698
rect 1592 5652 1644 5698
rect 1690 5652 1742 5698
rect 1788 5652 1840 5698
rect 1886 5652 1938 5698
rect 1984 5652 2036 5698
rect 2082 5652 2134 5698
rect 2180 5652 2232 5698
rect 2278 5652 2330 5698
rect 2376 5652 2428 5698
rect 2474 5652 2526 5698
rect 2572 5652 2624 5698
rect 2670 5652 2722 5698
rect 2768 5652 2820 5698
rect 2866 5652 2918 5698
rect 2964 5652 3016 5698
rect 3062 5652 3114 5698
rect 3160 5652 3212 5698
rect 3258 5652 3310 5698
rect 3356 5652 3408 5698
rect 3454 5652 3506 5698
rect 3552 5652 3604 5698
rect 3650 5652 3702 5698
rect 3748 5652 3800 5698
rect 3846 5652 3898 5698
rect 3944 5652 3996 5698
rect 4042 5652 4094 5698
rect 4140 5652 4192 5698
rect 4238 5652 4290 5698
rect 4336 5652 4388 5698
rect 4434 5652 4486 5698
rect 4532 5652 4584 5698
rect 4630 5652 4682 5698
rect 4728 5652 4780 5698
rect 4826 5652 4878 5698
rect 4924 5652 4976 5698
rect 5022 5652 5074 5698
rect 5120 5652 5172 5698
rect 5218 5652 5270 5698
rect 5316 5652 5368 5698
rect 5414 5652 5466 5698
rect 5512 5652 5564 5698
rect 5610 5652 5662 5698
rect 5708 5652 5760 5698
rect 5806 5652 5858 5698
rect 5904 5652 5956 5698
rect 6002 5652 6054 5698
rect 6100 5652 6152 5698
rect 6198 5652 6250 5698
rect 6296 5652 6348 5698
rect 6394 5652 6446 5698
rect 6492 5652 6544 5698
rect 6590 5652 6642 5698
rect 6688 5652 6740 5698
rect 6786 5652 6838 5698
rect 6884 5652 6936 5698
rect 6982 5652 7034 5698
rect 7080 5652 7132 5698
rect 7178 5652 7230 5698
rect 7276 5652 7328 5698
rect 7374 5652 7426 5698
rect 7472 5652 7524 5698
rect 7570 5652 7622 5698
rect 7668 5652 7720 5698
rect 7766 5652 7818 5698
rect 7864 5652 7916 5698
rect 7962 5652 8014 5698
rect 8060 5652 8112 5698
rect 8158 5652 8210 5698
rect 8256 5652 8308 5698
rect 8354 5652 8406 5698
rect 8452 5652 8504 5698
rect 8550 5652 8602 5698
rect 8648 5652 8700 5698
rect 8746 5652 8798 5698
rect 8844 5652 8896 5698
rect 8942 5652 8994 5698
rect 9040 5652 9092 5698
rect 9138 5652 9190 5698
rect 9236 5652 9288 5698
rect 9334 5652 9386 5698
rect 9432 5652 9484 5698
rect 9530 5652 9582 5698
rect 9628 5652 9680 5698
rect 9726 5652 9778 5698
rect 9824 5652 9876 5698
rect 9922 5652 10006 5698
rect 24 5648 10006 5652
rect 10052 5648 10069 5698
rect -39 5635 10069 5648
rect -39 5596 41 5635
rect -39 5550 -22 5596
rect 24 5550 41 5596
rect -39 5498 41 5550
rect -39 5452 -22 5498
rect 24 5452 41 5498
rect -39 5400 41 5452
rect 369 5406 438 5635
rect 9989 5596 10069 5635
rect 9989 5550 10006 5596
rect 10052 5550 10069 5596
rect 2454 5512 2644 5516
rect 2454 5503 2466 5512
rect 1556 5457 2466 5503
rect 1556 5406 1602 5457
rect 2454 5456 2466 5457
rect 2522 5456 2576 5512
rect 2632 5456 2644 5512
rect 2454 5452 2644 5456
rect 2906 5512 3096 5516
rect 2906 5456 2918 5512
rect 2974 5456 3028 5512
rect 3084 5503 3096 5512
rect 6934 5512 7124 5516
rect 6934 5503 6946 5512
rect 3084 5457 3994 5503
rect 3084 5456 3096 5457
rect 2906 5452 3096 5456
rect 1695 5406 1895 5410
rect 2052 5406 2102 5408
rect 3448 5406 3498 5408
rect 3655 5406 3855 5410
rect 3948 5406 3994 5457
rect 6036 5457 6946 5503
rect 6036 5406 6082 5457
rect 6934 5456 6946 5457
rect 7002 5456 7056 5512
rect 7112 5456 7124 5512
rect 6934 5452 7124 5456
rect 7386 5512 7576 5516
rect 7386 5456 7398 5512
rect 7454 5456 7508 5512
rect 7564 5503 7576 5512
rect 7564 5457 8474 5503
rect 7564 5456 7576 5457
rect 7386 5452 7576 5456
rect 6175 5406 6375 5410
rect 6532 5406 6582 5408
rect 7928 5406 7978 5408
rect 8135 5406 8335 5410
rect 8428 5406 8474 5457
rect 9989 5498 10069 5550
rect 9989 5452 10006 5498
rect 10052 5452 10069 5498
rect 9989 5412 10069 5452
rect 9720 5406 10069 5412
rect -39 5354 -22 5400
rect 24 5354 41 5400
rect 297 5360 308 5406
rect 482 5360 493 5406
rect 577 5360 588 5406
rect 762 5360 868 5406
rect 1042 5360 1064 5406
rect 1137 5360 1148 5406
rect 1322 5360 1333 5406
rect 1417 5360 1428 5406
rect 1602 5360 1613 5406
rect 1695 5360 1708 5406
rect 1882 5360 1895 5406
rect 1977 5360 1988 5406
rect 2162 5360 2173 5406
rect 2257 5360 2268 5406
rect 2442 5360 2548 5406
rect 2722 5360 2733 5406
rect 2817 5360 2828 5406
rect 3002 5360 3108 5406
rect 3282 5360 3293 5406
rect 3377 5360 3388 5406
rect 3562 5360 3573 5406
rect 3655 5360 3668 5406
rect 3842 5360 3855 5406
rect 3937 5360 3948 5406
rect 4122 5360 4133 5406
rect 4217 5360 4228 5406
rect 4402 5360 4413 5406
rect 4486 5360 4508 5406
rect 4682 5360 4788 5406
rect 4962 5360 4973 5406
rect 5057 5360 5068 5406
rect 5242 5360 5348 5406
rect 5522 5360 5544 5406
rect 5617 5360 5628 5406
rect 5802 5360 5813 5406
rect 5897 5360 5908 5406
rect 6082 5360 6093 5406
rect 6175 5360 6188 5406
rect 6362 5360 6375 5406
rect 6457 5360 6468 5406
rect 6642 5360 6653 5406
rect 6737 5360 6748 5406
rect 6922 5360 7028 5406
rect 7202 5360 7213 5406
rect 7297 5360 7308 5406
rect 7482 5360 7588 5406
rect 7762 5360 7773 5406
rect 7857 5360 7868 5406
rect 8042 5360 8053 5406
rect 8135 5360 8148 5406
rect 8322 5360 8335 5406
rect 8417 5360 8428 5406
rect 8602 5360 8613 5406
rect 8697 5360 8708 5406
rect 8882 5360 8893 5406
rect 8966 5360 8988 5406
rect 9162 5360 9268 5406
rect 9442 5360 9453 5406
rect 9537 5360 9548 5406
rect 9722 5400 10069 5406
rect 9722 5360 10006 5400
rect -39 5302 41 5354
rect -39 5256 -22 5302
rect 24 5256 41 5302
rect -39 5204 41 5256
rect -39 5158 -22 5204
rect 24 5158 41 5204
rect -39 5106 41 5158
rect -39 5060 -22 5106
rect 24 5060 41 5106
rect 369 5074 438 5360
rect 588 5074 669 5360
rect 1192 5208 1249 5360
rect 1695 5345 1709 5360
rect 1765 5345 1819 5360
rect 1875 5345 1895 5360
rect 1695 5333 1895 5345
rect 2052 5304 2102 5360
rect 3448 5304 3498 5360
rect 3655 5345 3675 5360
rect 3731 5345 3785 5360
rect 3841 5345 3855 5360
rect 3655 5333 3855 5345
rect 2052 5254 3498 5304
rect 4301 5208 4358 5360
rect 1192 5151 4358 5208
rect 5672 5208 5729 5360
rect 6175 5345 6189 5360
rect 6245 5345 6299 5360
rect 6355 5345 6375 5360
rect 6175 5333 6375 5345
rect 6532 5304 6582 5360
rect 7928 5304 7978 5360
rect 8135 5345 8155 5360
rect 8211 5345 8265 5360
rect 8321 5345 8335 5360
rect 8135 5333 8335 5345
rect 6532 5254 7978 5304
rect 8781 5208 8838 5360
rect 9720 5355 10006 5360
rect 5672 5151 8838 5208
rect 9989 5354 10006 5355
rect 10052 5354 10069 5400
rect 9989 5302 10069 5354
rect 9989 5256 10006 5302
rect 10052 5256 10069 5302
rect 9989 5204 10069 5256
rect 9989 5158 10006 5204
rect 10052 5158 10069 5204
rect 9989 5106 10069 5158
rect 855 5086 1055 5100
rect -39 5008 41 5060
rect 297 5028 308 5074
rect 482 5028 493 5074
rect 577 5028 588 5074
rect 762 5028 773 5074
rect 855 5030 867 5086
rect 923 5074 975 5086
rect 1031 5074 1055 5086
rect 1415 5093 1615 5101
rect 855 5028 868 5030
rect 1042 5028 1055 5074
rect 1137 5028 1148 5074
rect 1322 5028 1333 5074
rect 1415 5028 1428 5093
rect 1484 5074 1538 5093
rect 1594 5074 1615 5093
rect 1602 5028 1615 5074
rect -39 4962 -22 5008
rect 24 4962 41 5008
rect -39 4910 41 4962
rect -39 4864 -22 4910
rect 24 4864 41 4910
rect 333 4967 530 4972
rect 333 4911 349 4967
rect 405 4911 459 4967
rect 515 4962 530 4967
rect 588 4962 634 5028
rect 855 5023 1055 5028
rect 515 4916 634 4962
rect 515 4911 530 4916
rect 333 4906 530 4911
rect -39 4812 41 4864
rect -236 4752 -170 4767
rect -236 4696 -231 4752
rect -175 4696 -170 4752
rect -236 4642 -170 4696
rect -236 4586 -231 4642
rect -175 4586 -170 4642
rect -236 4570 -170 4586
rect -39 4766 -22 4812
rect 24 4766 41 4812
rect -39 4763 41 4766
rect 714 4900 1029 4904
rect 714 4844 851 4900
rect 907 4844 961 4900
rect 1017 4844 1029 4900
rect 714 4838 1029 4844
rect 1155 4857 1201 5028
rect 1415 5024 1615 5028
rect 1695 5090 1895 5101
rect 1695 5074 1709 5090
rect 1765 5074 1819 5090
rect 1875 5074 1895 5090
rect 2255 5087 2455 5101
rect 1695 5028 1708 5074
rect 1882 5028 1895 5074
rect 1977 5028 1988 5074
rect 2162 5028 2173 5074
rect 2255 5031 2267 5087
rect 2323 5074 2377 5087
rect 2433 5074 2455 5087
rect 3095 5087 3295 5101
rect 3095 5074 3117 5087
rect 3173 5074 3227 5087
rect 2255 5028 2268 5031
rect 2442 5028 2455 5074
rect 2537 5028 2548 5074
rect 2722 5028 2828 5074
rect 3002 5028 3013 5074
rect 3095 5028 3108 5074
rect 3283 5031 3295 5087
rect 3655 5090 3855 5101
rect 3655 5074 3675 5090
rect 3731 5074 3785 5090
rect 3841 5074 3855 5090
rect 3282 5028 3295 5031
rect 3377 5028 3388 5074
rect 3562 5028 3573 5074
rect 3655 5028 3668 5074
rect 3842 5028 3855 5074
rect 1695 5024 1895 5028
rect 1250 4966 1442 4968
rect 1988 4966 2038 5028
rect 2255 5024 2455 5028
rect 3095 5024 3295 5028
rect 1250 4965 2038 4966
rect 1250 4909 1262 4965
rect 1318 4909 1372 4965
rect 1428 4920 2038 4965
rect 3512 4966 3562 5028
rect 3655 5024 3855 5028
rect 3935 5093 4135 5101
rect 3935 5074 3956 5093
rect 4012 5074 4066 5093
rect 3935 5028 3948 5074
rect 4122 5028 4135 5093
rect 4495 5086 4695 5100
rect 4495 5074 4519 5086
rect 4575 5074 4627 5086
rect 4217 5028 4228 5074
rect 4402 5028 4413 5074
rect 4495 5028 4508 5074
rect 4683 5030 4695 5086
rect 5335 5086 5535 5100
rect 4682 5028 4695 5030
rect 4777 5028 4788 5074
rect 4962 5028 4973 5074
rect 5057 5028 5068 5074
rect 5242 5028 5253 5074
rect 5335 5030 5347 5086
rect 5403 5074 5455 5086
rect 5511 5074 5535 5086
rect 5895 5093 6095 5101
rect 5335 5028 5348 5030
rect 5522 5028 5535 5074
rect 5617 5028 5628 5074
rect 5802 5028 5813 5074
rect 5895 5028 5908 5093
rect 5964 5074 6018 5093
rect 6074 5074 6095 5093
rect 6082 5028 6095 5074
rect 3935 5024 4135 5028
rect 4108 4966 4300 4968
rect 3512 4965 4300 4966
rect 3512 4920 4122 4965
rect 1428 4909 1442 4920
rect 1250 4906 1442 4909
rect 4108 4909 4122 4920
rect 4178 4909 4232 4965
rect 4288 4909 4300 4965
rect 4108 4906 4300 4909
rect 4349 4857 4395 5028
rect 4495 5023 4695 5028
rect 4916 4982 4962 5028
rect 5068 4982 5114 5028
rect 5335 5023 5535 5028
rect 4884 4936 5114 4982
rect -39 4754 348 4763
rect 714 4754 762 4838
rect 1155 4811 2038 4857
rect 855 4754 1055 4756
rect -39 4714 308 4754
rect -39 4668 -22 4714
rect 24 4708 308 4714
rect 482 4708 493 4754
rect 577 4708 588 4754
rect 762 4708 773 4754
rect 855 4708 868 4754
rect 1042 4708 1055 4754
rect 24 4697 348 4708
rect 24 4668 41 4697
rect 855 4688 870 4708
rect 926 4688 980 4708
rect 1036 4688 1055 4708
rect 855 4678 1055 4688
rect 1135 4754 1335 4758
rect 1491 4754 1541 4755
rect 1775 4754 1825 4755
rect 1988 4754 2038 4811
rect 3512 4811 4395 4857
rect 4519 4899 4836 4904
rect 4519 4843 4531 4899
rect 4587 4843 4641 4899
rect 4697 4843 4836 4899
rect 4519 4838 4836 4843
rect 2255 4754 2455 4757
rect 1135 4708 1148 4754
rect 1322 4708 1335 4754
rect 1417 4708 1428 4754
rect 1602 4708 1613 4754
rect 1697 4708 1708 4754
rect 1882 4708 1893 4754
rect 1977 4708 1988 4754
rect 2162 4708 2173 4754
rect 2255 4708 2268 4754
rect 2442 4708 2455 4754
rect 1135 4694 1150 4708
rect 1206 4694 1260 4708
rect 1316 4694 1335 4708
rect 1135 4681 1335 4694
rect -39 4616 41 4668
rect -39 4570 -22 4616
rect 24 4570 41 4616
rect 96 4632 293 4636
rect 1491 4632 1541 4708
rect 96 4631 1541 4632
rect 96 4575 109 4631
rect 165 4575 219 4631
rect 275 4582 1541 4631
rect 1775 4630 1825 4708
rect 2255 4687 2269 4708
rect 2325 4687 2379 4708
rect 2435 4687 2455 4708
rect 2255 4677 2455 4687
rect 2535 4754 2735 4758
rect 2535 4689 2548 4754
rect 2722 4708 2735 4754
rect 2604 4689 2658 4708
rect 2714 4689 2735 4708
rect 2535 4681 2735 4689
rect 2815 4754 3015 4758
rect 2815 4708 2828 4754
rect 2815 4689 2836 4708
rect 2892 4689 2946 4708
rect 3002 4689 3015 4754
rect 2815 4681 3015 4689
rect 3095 4754 3295 4757
rect 3512 4754 3562 4811
rect 3725 4754 3775 4755
rect 4009 4754 4059 4755
rect 4215 4754 4415 4758
rect 3095 4708 3108 4754
rect 3282 4708 3295 4754
rect 3377 4708 3388 4754
rect 3562 4708 3573 4754
rect 3657 4708 3668 4754
rect 3842 4708 3853 4754
rect 3937 4708 3948 4754
rect 4122 4708 4133 4754
rect 4215 4708 4228 4754
rect 4402 4708 4415 4754
rect 3095 4687 3115 4708
rect 3171 4687 3225 4708
rect 3281 4687 3295 4708
rect 3095 4677 3295 4687
rect 3725 4630 3775 4708
rect 275 4575 293 4582
rect 1775 4580 3775 4630
rect 4009 4632 4059 4708
rect 4215 4694 4234 4708
rect 4290 4694 4344 4708
rect 4400 4694 4415 4708
rect 4215 4681 4415 4694
rect 4495 4754 4695 4756
rect 4788 4754 4836 4838
rect 5194 4900 5509 4904
rect 5194 4844 5331 4900
rect 5387 4844 5441 4900
rect 5497 4844 5509 4900
rect 5194 4838 5509 4844
rect 5635 4857 5681 5028
rect 5895 5024 6095 5028
rect 6175 5090 6375 5101
rect 6175 5074 6189 5090
rect 6245 5074 6299 5090
rect 6355 5074 6375 5090
rect 6735 5087 6935 5101
rect 6175 5028 6188 5074
rect 6362 5028 6375 5074
rect 6457 5028 6468 5074
rect 6642 5028 6653 5074
rect 6735 5031 6747 5087
rect 6803 5074 6857 5087
rect 6913 5074 6935 5087
rect 7575 5087 7775 5101
rect 7575 5074 7597 5087
rect 7653 5074 7707 5087
rect 6735 5028 6748 5031
rect 6922 5028 6935 5074
rect 7017 5028 7028 5074
rect 7202 5028 7308 5074
rect 7482 5028 7493 5074
rect 7575 5028 7588 5074
rect 7763 5031 7775 5087
rect 8135 5090 8335 5101
rect 8135 5074 8155 5090
rect 8211 5074 8265 5090
rect 8321 5074 8335 5090
rect 7762 5028 7775 5031
rect 7857 5028 7868 5074
rect 8042 5028 8053 5074
rect 8135 5028 8148 5074
rect 8322 5028 8335 5074
rect 6175 5024 6375 5028
rect 5730 4966 5922 4968
rect 6468 4966 6518 5028
rect 6735 5024 6935 5028
rect 7575 5024 7775 5028
rect 5730 4965 6518 4966
rect 5730 4909 5742 4965
rect 5798 4909 5852 4965
rect 5908 4920 6518 4965
rect 7992 4966 8042 5028
rect 8135 5024 8335 5028
rect 8415 5093 8615 5101
rect 8415 5074 8436 5093
rect 8492 5074 8546 5093
rect 8415 5028 8428 5074
rect 8602 5028 8615 5093
rect 8975 5086 9175 5100
rect 9989 5086 10006 5106
rect 8975 5074 8999 5086
rect 9055 5074 9107 5086
rect 8697 5028 8708 5074
rect 8882 5028 8893 5074
rect 8975 5028 8988 5074
rect 9163 5030 9175 5086
rect 9720 5074 10006 5086
rect 9162 5028 9175 5030
rect 9257 5028 9268 5074
rect 9442 5028 9453 5074
rect 9537 5028 9548 5074
rect 9722 5060 10006 5074
rect 10052 5060 10069 5106
rect 9722 5029 10069 5060
rect 9722 5028 9733 5029
rect 8415 5024 8615 5028
rect 8588 4966 8780 4968
rect 7992 4965 8780 4966
rect 7992 4920 8602 4965
rect 5908 4909 5922 4920
rect 5730 4906 5922 4909
rect 8588 4909 8602 4920
rect 8658 4909 8712 4965
rect 8768 4909 8780 4965
rect 8588 4906 8780 4909
rect 8829 4857 8875 5028
rect 8975 5023 9175 5028
rect 9396 4962 9442 5028
rect 9989 5008 10069 5029
rect 9700 4967 9897 4972
rect 9700 4962 9713 4967
rect 9396 4916 9713 4962
rect 9700 4911 9713 4916
rect 9771 4911 9823 4967
rect 9881 4911 9897 4967
rect 9700 4906 9897 4911
rect 9989 4962 10006 5008
rect 10052 4962 10069 5008
rect 9989 4910 10069 4962
rect 5194 4754 5242 4838
rect 5635 4811 6518 4857
rect 5335 4754 5535 4756
rect 4495 4708 4508 4754
rect 4682 4708 4695 4754
rect 4777 4708 4788 4754
rect 4962 4708 4973 4754
rect 5057 4708 5068 4754
rect 5242 4708 5253 4754
rect 5335 4708 5348 4754
rect 5522 4708 5535 4754
rect 4495 4688 4514 4708
rect 4570 4688 4624 4708
rect 4680 4688 4695 4708
rect 4495 4678 4695 4688
rect 5335 4688 5350 4708
rect 5406 4688 5460 4708
rect 5516 4688 5535 4708
rect 5335 4678 5535 4688
rect 5615 4754 5815 4758
rect 5971 4754 6021 4755
rect 6255 4754 6305 4755
rect 6468 4754 6518 4811
rect 7992 4811 8875 4857
rect 8999 4899 9316 4904
rect 8999 4843 9011 4899
rect 9067 4843 9121 4899
rect 9177 4843 9316 4899
rect 8999 4838 9316 4843
rect 6735 4754 6935 4757
rect 5615 4708 5628 4754
rect 5802 4708 5815 4754
rect 5897 4708 5908 4754
rect 6082 4708 6093 4754
rect 6177 4708 6188 4754
rect 6362 4708 6373 4754
rect 6457 4708 6468 4754
rect 6642 4708 6653 4754
rect 6735 4708 6748 4754
rect 6922 4708 6935 4754
rect 5615 4694 5630 4708
rect 5686 4694 5740 4708
rect 5796 4694 5815 4708
rect 5615 4681 5815 4694
rect 5971 4632 6021 4708
rect 4009 4582 6021 4632
rect 6255 4630 6305 4708
rect 6735 4687 6749 4708
rect 6805 4687 6859 4708
rect 6915 4687 6935 4708
rect 6735 4677 6935 4687
rect 7015 4754 7215 4758
rect 7015 4689 7028 4754
rect 7202 4708 7215 4754
rect 7084 4689 7138 4708
rect 7194 4689 7215 4708
rect 7015 4681 7215 4689
rect 7295 4754 7495 4758
rect 7295 4708 7308 4754
rect 7295 4689 7316 4708
rect 7372 4689 7426 4708
rect 7482 4689 7495 4754
rect 7295 4681 7495 4689
rect 7575 4754 7775 4757
rect 7992 4754 8042 4811
rect 8205 4754 8255 4755
rect 8489 4754 8539 4755
rect 8695 4754 8895 4758
rect 7575 4708 7588 4754
rect 7762 4708 7775 4754
rect 7857 4708 7868 4754
rect 8042 4708 8053 4754
rect 8137 4708 8148 4754
rect 8322 4708 8333 4754
rect 8417 4708 8428 4754
rect 8602 4708 8613 4754
rect 8695 4708 8708 4754
rect 8882 4708 8895 4754
rect 7575 4687 7595 4708
rect 7651 4687 7705 4708
rect 7761 4687 7775 4708
rect 7575 4677 7775 4687
rect 8205 4630 8255 4708
rect 6255 4580 8255 4630
rect 8489 4632 8539 4708
rect 8695 4694 8714 4708
rect 8770 4694 8824 4708
rect 8880 4694 8895 4708
rect 8695 4681 8895 4694
rect 8975 4754 9175 4756
rect 9268 4754 9316 4838
rect 9989 4864 10006 4910
rect 10052 4864 10069 4910
rect 9989 4812 10069 4864
rect 9989 4766 10006 4812
rect 10052 4766 10069 4812
rect 9989 4763 10069 4766
rect 9718 4754 10069 4763
rect 8975 4708 8988 4754
rect 9162 4708 9175 4754
rect 9257 4708 9268 4754
rect 9442 4708 9453 4754
rect 9537 4708 9548 4754
rect 9722 4714 10069 4754
rect 9722 4708 10006 4714
rect 8975 4688 8994 4708
rect 9050 4688 9104 4708
rect 9160 4688 9175 4708
rect 9718 4706 10006 4708
rect 8975 4678 9175 4688
rect 9989 4668 10006 4706
rect 10052 4668 10069 4714
rect 9485 4632 9682 4636
rect 8489 4631 9682 4632
rect 8489 4582 9503 4631
rect 96 4570 293 4575
rect -346 4447 -280 4462
rect -346 4391 -341 4447
rect -285 4391 -280 4447
rect -468 4325 -402 4340
rect -468 4269 -463 4325
rect -407 4269 -402 4325
rect -468 4215 -402 4269
rect -468 4159 -463 4215
rect -407 4159 -402 4215
rect -468 4153 -402 4159
rect -469 4143 -402 4153
rect -346 4337 -280 4391
rect -346 4281 -341 4337
rect -285 4281 -280 4337
rect -346 4265 -280 4281
rect -582 3733 -516 3748
rect -582 3677 -577 3733
rect -521 3677 -516 3733
rect -582 3623 -516 3677
rect -582 3567 -577 3623
rect -521 3567 -516 3623
rect -582 3553 -516 3567
rect -582 3551 -517 3553
rect -580 1319 -517 3551
rect -469 1911 -406 4143
rect -346 2033 -283 4265
rect -234 2338 -171 4570
rect -39 4518 41 4570
rect -39 4472 -22 4518
rect 24 4472 41 4518
rect -39 4443 41 4472
rect -39 4422 349 4443
rect 855 4438 1055 4448
rect -39 4420 308 4422
rect -39 4374 -22 4420
rect 24 4377 308 4420
rect 24 4374 41 4377
rect 297 4376 308 4377
rect 482 4376 493 4422
rect 577 4376 588 4422
rect 762 4376 773 4422
rect 855 4376 868 4438
rect 924 4422 978 4438
rect 1034 4422 1055 4438
rect 1042 4376 1055 4422
rect -39 4322 41 4374
rect -39 4276 -22 4322
rect 24 4276 41 4322
rect -39 4224 41 4276
rect 87 4326 284 4331
rect 87 4270 100 4326
rect 156 4270 210 4326
rect 266 4323 284 4326
rect 588 4323 634 4376
rect 855 4371 1055 4376
rect 1135 4439 1335 4449
rect 1135 4376 1148 4439
rect 1204 4422 1258 4439
rect 1314 4422 1335 4439
rect 2255 4437 2455 4449
rect 1987 4422 2037 4423
rect 2255 4422 2270 4437
rect 2326 4422 2380 4437
rect 2436 4422 2455 4437
rect 1322 4376 1335 4422
rect 1417 4376 1428 4422
rect 1602 4376 1708 4422
rect 1882 4376 1893 4422
rect 1977 4376 1988 4422
rect 2162 4376 2173 4422
rect 2255 4376 2268 4422
rect 2442 4376 2455 4422
rect 2537 4437 2734 4442
rect 2537 4422 2553 4437
rect 2609 4422 2663 4437
rect 2719 4422 2734 4437
rect 2817 4437 3014 4442
rect 2817 4422 2833 4437
rect 2889 4422 2943 4437
rect 2999 4422 3014 4437
rect 2537 4376 2548 4422
rect 2722 4376 2828 4422
rect 3002 4376 3014 4422
rect 3095 4437 3295 4449
rect 3095 4422 3114 4437
rect 3170 4422 3224 4437
rect 3280 4422 3295 4437
rect 4215 4439 4415 4449
rect 3513 4422 3563 4423
rect 4215 4422 4236 4439
rect 4292 4422 4346 4439
rect 3095 4376 3108 4422
rect 3282 4376 3295 4422
rect 3377 4376 3388 4422
rect 3562 4376 3573 4422
rect 3657 4376 3668 4422
rect 3842 4376 3948 4422
rect 4122 4376 4133 4422
rect 4215 4376 4228 4422
rect 4402 4376 4415 4439
rect 1135 4372 1335 4376
rect 266 4277 634 4323
rect 1987 4320 2037 4376
rect 2255 4371 2455 4376
rect 3095 4371 3295 4376
rect 266 4270 284 4277
rect 87 4265 284 4270
rect 1154 4274 2037 4320
rect 3513 4320 3563 4376
rect 4215 4372 4415 4376
rect 4495 4438 4695 4448
rect 4495 4422 4516 4438
rect 4572 4422 4626 4438
rect 4495 4376 4508 4422
rect 4682 4376 4695 4438
rect 5335 4438 5535 4448
rect 4777 4376 4788 4422
rect 4962 4376 4973 4422
rect 5057 4376 5068 4422
rect 5242 4376 5253 4422
rect 5335 4376 5348 4438
rect 5404 4422 5458 4438
rect 5514 4422 5535 4438
rect 5522 4376 5535 4422
rect 4495 4371 4695 4376
rect 4916 4330 4962 4376
rect 5068 4330 5114 4376
rect 5335 4371 5535 4376
rect 5615 4439 5815 4449
rect 5615 4376 5628 4439
rect 5684 4422 5738 4439
rect 5794 4422 5815 4439
rect 6735 4437 6935 4449
rect 6467 4422 6517 4423
rect 6735 4422 6750 4437
rect 6806 4422 6860 4437
rect 6916 4422 6935 4437
rect 7575 4437 7775 4449
rect 7575 4422 7594 4437
rect 7650 4422 7704 4437
rect 7760 4422 7775 4437
rect 8695 4439 8895 4449
rect 7993 4422 8043 4423
rect 8695 4422 8716 4439
rect 8772 4422 8826 4439
rect 5802 4376 5815 4422
rect 5897 4376 5908 4422
rect 6082 4376 6188 4422
rect 6362 4376 6373 4422
rect 6457 4376 6468 4422
rect 6642 4376 6653 4422
rect 6735 4376 6748 4422
rect 6922 4376 6935 4422
rect 7017 4376 7028 4422
rect 7202 4376 7308 4422
rect 7482 4376 7493 4422
rect 7575 4376 7588 4422
rect 7762 4376 7775 4422
rect 7857 4376 7868 4422
rect 8042 4376 8053 4422
rect 8137 4376 8148 4422
rect 8322 4376 8428 4422
rect 8602 4376 8613 4422
rect 8695 4376 8708 4422
rect 8882 4376 8895 4439
rect 5615 4372 5815 4376
rect 3513 4274 4396 4320
rect 4884 4284 5114 4330
rect 6467 4320 6517 4376
rect 6735 4371 6935 4376
rect 7575 4371 7775 4376
rect -39 4178 -22 4224
rect 24 4178 41 4224
rect -39 4126 41 4178
rect 350 4209 547 4214
rect 350 4153 366 4209
rect 422 4153 476 4209
rect 532 4194 547 4209
rect 532 4153 634 4194
rect 350 4148 634 4153
rect -39 4080 -22 4126
rect 24 4103 41 4126
rect 24 4102 313 4103
rect 588 4102 634 4148
rect 855 4102 1055 4106
rect 1154 4102 1200 4274
rect 1249 4210 1329 4215
rect 1249 4154 1261 4210
rect 1317 4204 1329 4210
rect 4221 4210 4301 4215
rect 4221 4204 4233 4210
rect 1317 4158 2038 4204
rect 1317 4154 1329 4158
rect 1249 4148 1329 4154
rect 1415 4102 1615 4106
rect 24 4080 308 4102
rect -39 4056 308 4080
rect 482 4056 493 4102
rect 577 4056 588 4102
rect 762 4056 773 4102
rect -39 4028 41 4056
rect 855 4040 868 4102
rect 1042 4056 1055 4102
rect 1137 4056 1148 4102
rect 1322 4056 1333 4102
rect 1415 4056 1428 4102
rect 1602 4056 1615 4102
rect 924 4040 978 4056
rect 1034 4040 1055 4056
rect 855 4029 1055 4040
rect 1415 4039 1429 4056
rect 1485 4039 1539 4056
rect 1595 4039 1615 4056
rect 1415 4029 1615 4039
rect 1695 4102 1895 4106
rect 1988 4102 2038 4158
rect 3512 4158 4233 4204
rect 3512 4102 3562 4158
rect 4221 4154 4233 4158
rect 4289 4154 4301 4210
rect 4221 4148 4301 4154
rect 3655 4102 3855 4106
rect 1695 4056 1708 4102
rect 1882 4056 1895 4102
rect 1977 4056 1988 4102
rect 2162 4056 2173 4102
rect 2257 4056 2268 4102
rect 2442 4056 2548 4102
rect 2722 4056 2733 4102
rect 2817 4056 2828 4102
rect 3002 4056 3108 4102
rect 3282 4056 3293 4102
rect 3377 4056 3388 4102
rect 3562 4056 3573 4102
rect 3655 4056 3668 4102
rect 3842 4056 3855 4102
rect 1695 4040 1710 4056
rect 1766 4040 1820 4056
rect 1876 4040 1895 4056
rect 1695 4029 1895 4040
rect 3655 4040 3674 4056
rect 3730 4040 3784 4056
rect 3840 4040 3855 4056
rect 3655 4029 3855 4040
rect 3935 4102 4135 4106
rect 4350 4102 4396 4274
rect 5634 4274 6517 4320
rect 7993 4320 8043 4376
rect 8695 4372 8895 4376
rect 8975 4438 9175 4448
rect 8975 4422 8996 4438
rect 9052 4422 9106 4438
rect 8975 4376 8988 4422
rect 9162 4376 9175 4438
rect 9268 4422 9326 4582
rect 9485 4575 9503 4582
rect 9559 4575 9613 4631
rect 9669 4575 9682 4631
rect 9485 4570 9682 4575
rect 9989 4616 10069 4668
rect 9989 4570 10006 4616
rect 10052 4570 10069 4616
rect 9989 4518 10069 4570
rect 9989 4472 10006 4518
rect 10052 4472 10069 4518
rect 9989 4425 10069 4472
rect 9717 4422 10069 4425
rect 9257 4376 9268 4422
rect 9442 4376 9453 4422
rect 9537 4376 9548 4422
rect 9722 4420 10069 4422
rect 9722 4376 10006 4420
rect 8975 4371 9175 4376
rect 9717 4374 10006 4376
rect 10052 4374 10069 4420
rect 9717 4368 10069 4374
rect 9989 4322 10069 4368
rect 7993 4274 8876 4320
rect 4884 4148 5114 4194
rect 4495 4102 4695 4106
rect 4916 4102 4962 4148
rect 5068 4102 5114 4148
rect 5335 4102 5535 4106
rect 5634 4102 5680 4274
rect 5729 4210 5809 4215
rect 5729 4154 5741 4210
rect 5797 4204 5809 4210
rect 8701 4210 8781 4215
rect 8701 4204 8713 4210
rect 5797 4158 6518 4204
rect 5797 4154 5809 4158
rect 5729 4148 5809 4154
rect 5895 4102 6095 4106
rect 3935 4056 3948 4102
rect 4122 4056 4135 4102
rect 4217 4056 4228 4102
rect 4402 4056 4413 4102
rect 4495 4056 4508 4102
rect 3935 4039 3955 4056
rect 4011 4039 4065 4056
rect 4121 4039 4135 4056
rect 3935 4029 4135 4039
rect 4495 4040 4516 4056
rect 4572 4040 4626 4056
rect 4682 4040 4695 4102
rect 4777 4056 4788 4102
rect 4962 4056 4973 4102
rect 5057 4056 5068 4102
rect 5242 4056 5253 4102
rect 4495 4029 4695 4040
rect 5335 4040 5348 4102
rect 5522 4056 5535 4102
rect 5617 4056 5628 4102
rect 5802 4056 5813 4102
rect 5895 4056 5908 4102
rect 6082 4056 6095 4102
rect 5404 4040 5458 4056
rect 5514 4040 5535 4056
rect 5335 4029 5535 4040
rect 5895 4039 5909 4056
rect 5965 4039 6019 4056
rect 6075 4039 6095 4056
rect 5895 4029 6095 4039
rect 6175 4102 6375 4106
rect 6468 4102 6518 4158
rect 7992 4158 8713 4204
rect 7992 4102 8042 4158
rect 8701 4154 8713 4158
rect 8769 4154 8781 4210
rect 8701 4148 8781 4154
rect 8135 4102 8335 4106
rect 6175 4056 6188 4102
rect 6362 4056 6375 4102
rect 6457 4056 6468 4102
rect 6642 4056 6653 4102
rect 6737 4056 6748 4102
rect 6922 4056 7028 4102
rect 7202 4056 7213 4102
rect 7297 4056 7308 4102
rect 7482 4056 7588 4102
rect 7762 4056 7773 4102
rect 7857 4056 7868 4102
rect 8042 4056 8053 4102
rect 8135 4056 8148 4102
rect 8322 4056 8335 4102
rect 6175 4040 6190 4056
rect 6246 4040 6300 4056
rect 6356 4040 6375 4056
rect 6175 4029 6375 4040
rect 8135 4040 8154 4056
rect 8210 4040 8264 4056
rect 8320 4040 8335 4056
rect 8135 4029 8335 4040
rect 8415 4102 8615 4106
rect 8830 4102 8876 4274
rect 9989 4276 10006 4322
rect 10052 4276 10069 4322
rect 9989 4224 10069 4276
rect 9484 4209 9681 4214
rect 9484 4195 9502 4209
rect 9442 4194 9502 4195
rect 9396 4153 9502 4194
rect 9558 4153 9612 4209
rect 9668 4153 9681 4209
rect 9396 4148 9681 4153
rect 9989 4178 10006 4224
rect 10052 4178 10069 4224
rect 8975 4102 9175 4106
rect 9396 4102 9442 4148
rect 9989 4126 10069 4178
rect 9989 4107 10006 4126
rect 8415 4056 8428 4102
rect 8602 4056 8615 4102
rect 8697 4056 8708 4102
rect 8882 4056 8893 4102
rect 8975 4056 8988 4102
rect 8415 4039 8435 4056
rect 8491 4039 8545 4056
rect 8601 4039 8615 4056
rect 8415 4029 8615 4039
rect 8975 4040 8996 4056
rect 9052 4040 9106 4056
rect 9162 4040 9175 4102
rect 9257 4056 9268 4102
rect 9442 4056 9453 4102
rect 9537 4056 9548 4102
rect 9722 4080 10006 4107
rect 10052 4080 10069 4126
rect 9722 4050 10069 4080
rect 8975 4029 9175 4040
rect -39 3982 -22 4028
rect 24 3982 41 4028
rect 9989 4028 10069 4050
rect -39 3930 41 3982
rect -39 3884 -22 3930
rect 24 3884 41 3930
rect 88 3985 285 3990
rect 88 3929 101 3985
rect 157 3929 211 3985
rect 267 3983 285 3985
rect 9733 3985 9935 3990
rect 9733 3983 9751 3985
rect 267 3933 2038 3983
rect 267 3929 285 3933
rect 88 3924 285 3929
rect -39 3832 41 3884
rect -39 3786 -22 3832
rect 24 3786 41 3832
rect -39 3777 41 3786
rect 857 3793 1054 3798
rect -39 3770 327 3777
rect 857 3770 870 3793
rect 926 3770 980 3793
rect 1036 3770 1054 3793
rect 1415 3795 1612 3800
rect -39 3734 308 3770
rect -39 3688 -22 3734
rect 24 3724 308 3734
rect 482 3724 493 3770
rect 577 3724 588 3770
rect 762 3724 868 3770
rect 1042 3732 1054 3770
rect 1042 3724 1053 3732
rect 1137 3724 1148 3770
rect 1322 3724 1333 3770
rect 1415 3734 1428 3795
rect 1484 3770 1538 3795
rect 1594 3770 1612 3795
rect 1988 3770 2038 3933
rect 3512 3933 6518 3983
rect 2255 3782 2455 3797
rect 1417 3724 1428 3734
rect 1602 3724 1613 3770
rect 1697 3724 1708 3770
rect 1882 3724 1893 3770
rect 1977 3724 1988 3770
rect 2162 3724 2173 3770
rect 2255 3726 2267 3782
rect 2323 3770 2377 3782
rect 2433 3770 2455 3782
rect 3095 3782 3295 3797
rect 3095 3770 3117 3782
rect 3173 3770 3227 3782
rect 2255 3724 2268 3726
rect 2442 3724 2455 3770
rect 2537 3724 2548 3770
rect 2722 3724 2828 3770
rect 3002 3724 3013 3770
rect 3095 3724 3108 3770
rect 3283 3726 3295 3782
rect 3512 3770 3562 3933
rect 4333 3822 5697 3872
rect 4333 3796 4402 3822
rect 4332 3770 4402 3796
rect 5628 3796 5697 3822
rect 5628 3770 5698 3796
rect 6468 3770 6518 3933
rect 7992 3933 9751 3983
rect 6735 3782 6935 3797
rect 3282 3724 3295 3726
rect 3377 3724 3388 3770
rect 3562 3724 3573 3770
rect 3657 3724 3668 3770
rect 3842 3724 3853 3770
rect 3937 3724 3948 3770
rect 4122 3724 4133 3770
rect 4217 3724 4228 3770
rect 4402 3724 4413 3770
rect 4497 3724 4508 3770
rect 4682 3724 4788 3770
rect 4962 3724 4973 3770
rect 5057 3724 5068 3770
rect 5242 3724 5348 3770
rect 5522 3724 5533 3770
rect 5617 3724 5628 3770
rect 5802 3724 5813 3770
rect 5897 3724 5908 3770
rect 6082 3724 6093 3770
rect 6177 3724 6188 3770
rect 6362 3724 6373 3770
rect 6457 3724 6468 3770
rect 6642 3724 6653 3770
rect 6735 3726 6747 3782
rect 6803 3770 6857 3782
rect 6913 3770 6935 3782
rect 7575 3782 7775 3797
rect 7575 3770 7597 3782
rect 7653 3770 7707 3782
rect 6735 3724 6748 3726
rect 6922 3724 6935 3770
rect 7017 3724 7028 3770
rect 7202 3724 7308 3770
rect 7482 3724 7493 3770
rect 7575 3724 7588 3770
rect 7763 3726 7775 3782
rect 7992 3770 8042 3933
rect 9733 3929 9751 3933
rect 9807 3929 9861 3985
rect 9917 3929 9935 3985
rect 9733 3924 9935 3929
rect 9989 3982 10006 4028
rect 10052 3982 10069 4028
rect 9989 3930 10069 3982
rect 9483 3882 9680 3887
rect 9483 3872 9501 3882
rect 8813 3826 9501 3872
rect 9557 3826 9611 3882
rect 9667 3826 9680 3882
rect 8813 3822 9680 3826
rect 8813 3796 8882 3822
rect 9483 3821 9680 3822
rect 9989 3884 10006 3930
rect 10052 3884 10069 3930
rect 9989 3832 10069 3884
rect 8812 3770 8882 3796
rect 9989 3786 10006 3832
rect 10052 3786 10069 3832
rect 9989 3777 10069 3786
rect 9710 3770 10069 3777
rect 7762 3724 7775 3726
rect 7857 3724 7868 3770
rect 8042 3724 8053 3770
rect 8137 3724 8148 3770
rect 8322 3724 8333 3770
rect 8417 3724 8428 3770
rect 8602 3724 8613 3770
rect 8697 3724 8708 3770
rect 8882 3724 8893 3770
rect 8977 3724 8988 3770
rect 9162 3724 9268 3770
rect 9442 3724 9453 3770
rect 9537 3724 9548 3770
rect 9722 3734 10069 3770
rect 9722 3724 10006 3734
rect 24 3720 327 3724
rect 24 3688 41 3720
rect -39 3636 41 3688
rect -39 3590 -22 3636
rect 24 3590 41 3636
rect -39 3538 41 3590
rect 92 3612 289 3617
rect 92 3556 105 3612
rect 161 3556 215 3612
rect 271 3610 289 3612
rect 1232 3610 1322 3724
rect 1429 3610 1482 3724
rect 271 3557 1482 3610
rect 271 3556 289 3557
rect 92 3551 289 3556
rect 1429 3550 1482 3557
rect 1827 3605 1880 3724
rect 2255 3720 2455 3724
rect 3095 3720 3295 3724
rect 3670 3605 3723 3724
rect 1827 3552 3723 3605
rect 4068 3610 4121 3724
rect 5909 3610 5962 3724
rect 4068 3557 5962 3610
rect 4068 3550 4121 3557
rect 5909 3550 5962 3557
rect 6307 3605 6360 3724
rect 6735 3720 6935 3724
rect 7575 3720 7775 3724
rect 8150 3605 8203 3724
rect 6307 3552 8203 3605
rect 8548 3610 8601 3724
rect 9710 3720 10006 3724
rect 9989 3688 10006 3720
rect 10052 3688 10069 3734
rect 9989 3636 10069 3688
rect 9713 3612 9910 3617
rect 9713 3610 9731 3612
rect 8548 3557 9731 3610
rect 8548 3550 8601 3557
rect 9713 3556 9731 3557
rect 9787 3556 9841 3612
rect 9897 3556 9910 3612
rect 9713 3551 9910 3556
rect 9989 3590 10006 3636
rect 10052 3590 10069 3636
rect -39 3492 -22 3538
rect 24 3492 41 3538
rect -39 3457 41 3492
rect 9989 3538 10069 3590
rect 9989 3492 10006 3538
rect 10052 3492 10069 3538
rect 9989 3457 10069 3492
rect -39 3440 10069 3457
rect -39 3394 -22 3440
rect 24 3394 76 3440
rect 122 3394 174 3440
rect 220 3394 272 3440
rect 318 3394 370 3440
rect 416 3394 468 3440
rect 514 3394 566 3440
rect 612 3394 664 3440
rect 710 3394 762 3440
rect 808 3394 860 3440
rect 906 3394 958 3440
rect 1004 3394 1056 3440
rect 1102 3394 1154 3440
rect 1200 3394 1252 3440
rect 1298 3394 1350 3440
rect 1396 3394 1448 3440
rect 1494 3394 1546 3440
rect 1592 3394 1644 3440
rect 1690 3394 1742 3440
rect 1788 3394 1840 3440
rect 1886 3394 1938 3440
rect 1984 3394 2036 3440
rect 2082 3394 2134 3440
rect 2180 3394 2232 3440
rect 2278 3394 2330 3440
rect 2376 3394 2428 3440
rect 2474 3394 2526 3440
rect 2572 3394 2624 3440
rect 2670 3394 2722 3440
rect 2768 3394 2820 3440
rect 2866 3394 2918 3440
rect 2964 3394 3016 3440
rect 3062 3394 3114 3440
rect 3160 3394 3212 3440
rect 3258 3394 3310 3440
rect 3356 3394 3408 3440
rect 3454 3394 3506 3440
rect 3552 3394 3604 3440
rect 3650 3394 3702 3440
rect 3748 3394 3800 3440
rect 3846 3394 3898 3440
rect 3944 3394 3996 3440
rect 4042 3394 4094 3440
rect 4140 3394 4192 3440
rect 4238 3394 4290 3440
rect 4336 3394 4388 3440
rect 4434 3394 4486 3440
rect 4532 3394 4584 3440
rect 4630 3394 4682 3440
rect 4728 3394 4780 3440
rect 4826 3394 4878 3440
rect 4924 3394 4976 3440
rect 5022 3394 5074 3440
rect 5120 3394 5172 3440
rect 5218 3394 5270 3440
rect 5316 3394 5368 3440
rect 5414 3394 5466 3440
rect 5512 3394 5564 3440
rect 5610 3394 5662 3440
rect 5708 3394 5760 3440
rect 5806 3394 5858 3440
rect 5904 3394 5956 3440
rect 6002 3394 6054 3440
rect 6100 3394 6152 3440
rect 6198 3394 6250 3440
rect 6296 3394 6348 3440
rect 6394 3394 6446 3440
rect 6492 3394 6544 3440
rect 6590 3394 6642 3440
rect 6688 3394 6740 3440
rect 6786 3394 6838 3440
rect 6884 3394 6936 3440
rect 6982 3394 7034 3440
rect 7080 3394 7132 3440
rect 7178 3394 7230 3440
rect 7276 3394 7328 3440
rect 7374 3394 7426 3440
rect 7472 3394 7524 3440
rect 7570 3394 7622 3440
rect 7668 3394 7720 3440
rect 7766 3394 7818 3440
rect 7864 3394 7916 3440
rect 7962 3394 8014 3440
rect 8060 3394 8112 3440
rect 8158 3394 8210 3440
rect 8256 3394 8308 3440
rect 8354 3394 8406 3440
rect 8452 3394 8504 3440
rect 8550 3394 8602 3440
rect 8648 3394 8700 3440
rect 8746 3394 8798 3440
rect 8844 3394 8896 3440
rect 8942 3394 8994 3440
rect 9040 3394 9092 3440
rect 9138 3394 9190 3440
rect 9236 3394 9288 3440
rect 9334 3394 9386 3440
rect 9432 3394 9484 3440
rect 9530 3394 9582 3440
rect 9628 3394 9680 3440
rect 9726 3394 9778 3440
rect 9824 3394 9876 3440
rect 9922 3394 10006 3440
rect 10052 3394 10069 3440
rect -39 3377 10069 3394
rect 10122 4645 10185 4660
rect 10122 4589 10127 4645
rect 10183 4589 10185 4645
rect 10122 4535 10185 4589
rect 10122 4479 10127 4535
rect 10183 4479 10185 4535
rect 54 3286 9950 3377
rect -39 3269 10069 3286
rect -39 3219 -22 3269
rect 24 3223 76 3269
rect 122 3223 174 3269
rect 220 3223 272 3269
rect 318 3223 370 3269
rect 416 3223 468 3269
rect 514 3223 566 3269
rect 612 3223 664 3269
rect 710 3223 762 3269
rect 808 3223 860 3269
rect 906 3223 958 3269
rect 1004 3223 1056 3269
rect 1102 3223 1154 3269
rect 1200 3223 1252 3269
rect 1298 3223 1350 3269
rect 1396 3223 1448 3269
rect 1494 3223 1546 3269
rect 1592 3223 1644 3269
rect 1690 3223 1742 3269
rect 1788 3223 1840 3269
rect 1886 3223 1938 3269
rect 1984 3223 2036 3269
rect 2082 3223 2134 3269
rect 2180 3223 2232 3269
rect 2278 3223 2330 3269
rect 2376 3223 2428 3269
rect 2474 3223 2526 3269
rect 2572 3223 2624 3269
rect 2670 3223 2722 3269
rect 2768 3223 2820 3269
rect 2866 3223 2918 3269
rect 2964 3223 3016 3269
rect 3062 3223 3114 3269
rect 3160 3223 3212 3269
rect 3258 3223 3310 3269
rect 3356 3223 3408 3269
rect 3454 3223 3506 3269
rect 3552 3223 3604 3269
rect 3650 3223 3702 3269
rect 3748 3223 3800 3269
rect 3846 3223 3898 3269
rect 3944 3223 3996 3269
rect 4042 3223 4094 3269
rect 4140 3223 4192 3269
rect 4238 3223 4290 3269
rect 4336 3223 4388 3269
rect 4434 3223 4486 3269
rect 4532 3223 4584 3269
rect 4630 3223 4682 3269
rect 4728 3223 4780 3269
rect 4826 3223 4878 3269
rect 4924 3223 4976 3269
rect 5022 3223 5074 3269
rect 5120 3223 5172 3269
rect 5218 3223 5270 3269
rect 5316 3223 5368 3269
rect 5414 3223 5466 3269
rect 5512 3223 5564 3269
rect 5610 3223 5662 3269
rect 5708 3223 5760 3269
rect 5806 3223 5858 3269
rect 5904 3223 5956 3269
rect 6002 3223 6054 3269
rect 6100 3223 6152 3269
rect 6198 3223 6250 3269
rect 6296 3223 6348 3269
rect 6394 3223 6446 3269
rect 6492 3223 6544 3269
rect 6590 3223 6642 3269
rect 6688 3223 6740 3269
rect 6786 3223 6838 3269
rect 6884 3223 6936 3269
rect 6982 3223 7034 3269
rect 7080 3223 7132 3269
rect 7178 3223 7230 3269
rect 7276 3223 7328 3269
rect 7374 3223 7426 3269
rect 7472 3223 7524 3269
rect 7570 3223 7622 3269
rect 7668 3223 7720 3269
rect 7766 3223 7818 3269
rect 7864 3223 7916 3269
rect 7962 3223 8014 3269
rect 8060 3223 8112 3269
rect 8158 3223 8210 3269
rect 8256 3223 8308 3269
rect 8354 3223 8406 3269
rect 8452 3223 8504 3269
rect 8550 3223 8602 3269
rect 8648 3223 8700 3269
rect 8746 3223 8798 3269
rect 8844 3223 8896 3269
rect 8942 3223 8994 3269
rect 9040 3223 9092 3269
rect 9138 3223 9190 3269
rect 9236 3223 9288 3269
rect 9334 3223 9386 3269
rect 9432 3223 9484 3269
rect 9530 3223 9582 3269
rect 9628 3223 9680 3269
rect 9726 3223 9778 3269
rect 9824 3223 9876 3269
rect 9922 3223 10006 3269
rect 24 3219 10006 3223
rect 10052 3219 10069 3269
rect -39 3206 10069 3219
rect -39 3167 41 3206
rect -39 3121 -22 3167
rect 24 3121 41 3167
rect -39 3069 41 3121
rect -39 3023 -22 3069
rect 24 3023 41 3069
rect -39 2971 41 3023
rect 369 2977 438 3206
rect 9989 3167 10069 3206
rect 9989 3121 10006 3167
rect 10052 3121 10069 3167
rect 2454 3083 2644 3087
rect 2454 3074 2466 3083
rect 1556 3028 2466 3074
rect 1556 2977 1602 3028
rect 2454 3027 2466 3028
rect 2522 3027 2576 3083
rect 2632 3027 2644 3083
rect 2454 3023 2644 3027
rect 2906 3083 3096 3087
rect 2906 3027 2918 3083
rect 2974 3027 3028 3083
rect 3084 3074 3096 3083
rect 6934 3083 7124 3087
rect 6934 3074 6946 3083
rect 3084 3028 3994 3074
rect 3084 3027 3096 3028
rect 2906 3023 3096 3027
rect 1695 2977 1895 2981
rect 2052 2977 2102 2979
rect 3448 2977 3498 2979
rect 3655 2977 3855 2981
rect 3948 2977 3994 3028
rect 6036 3028 6946 3074
rect 6036 2977 6082 3028
rect 6934 3027 6946 3028
rect 7002 3027 7056 3083
rect 7112 3027 7124 3083
rect 6934 3023 7124 3027
rect 7386 3083 7576 3087
rect 7386 3027 7398 3083
rect 7454 3027 7508 3083
rect 7564 3074 7576 3083
rect 7564 3028 8474 3074
rect 7564 3027 7576 3028
rect 7386 3023 7576 3027
rect 6175 2977 6375 2981
rect 6532 2977 6582 2979
rect 7928 2977 7978 2979
rect 8135 2977 8335 2981
rect 8428 2977 8474 3028
rect 9989 3069 10069 3121
rect 9989 3023 10006 3069
rect 10052 3023 10069 3069
rect 9989 2983 10069 3023
rect 9720 2977 10069 2983
rect -39 2925 -22 2971
rect 24 2925 41 2971
rect 297 2931 308 2977
rect 482 2931 493 2977
rect 577 2931 588 2977
rect 762 2931 868 2977
rect 1042 2931 1064 2977
rect 1137 2931 1148 2977
rect 1322 2931 1333 2977
rect 1417 2931 1428 2977
rect 1602 2931 1613 2977
rect 1695 2931 1708 2977
rect 1882 2931 1895 2977
rect 1977 2931 1988 2977
rect 2162 2931 2173 2977
rect 2257 2931 2268 2977
rect 2442 2931 2548 2977
rect 2722 2931 2733 2977
rect 2817 2931 2828 2977
rect 3002 2931 3108 2977
rect 3282 2931 3293 2977
rect 3377 2931 3388 2977
rect 3562 2931 3573 2977
rect 3655 2931 3668 2977
rect 3842 2931 3855 2977
rect 3937 2931 3948 2977
rect 4122 2931 4133 2977
rect 4217 2931 4228 2977
rect 4402 2931 4413 2977
rect 4486 2931 4508 2977
rect 4682 2931 4788 2977
rect 4962 2931 4973 2977
rect 5057 2931 5068 2977
rect 5242 2931 5348 2977
rect 5522 2931 5544 2977
rect 5617 2931 5628 2977
rect 5802 2931 5813 2977
rect 5897 2931 5908 2977
rect 6082 2931 6093 2977
rect 6175 2931 6188 2977
rect 6362 2931 6375 2977
rect 6457 2931 6468 2977
rect 6642 2931 6653 2977
rect 6737 2931 6748 2977
rect 6922 2931 7028 2977
rect 7202 2931 7213 2977
rect 7297 2931 7308 2977
rect 7482 2931 7588 2977
rect 7762 2931 7773 2977
rect 7857 2931 7868 2977
rect 8042 2931 8053 2977
rect 8135 2931 8148 2977
rect 8322 2931 8335 2977
rect 8417 2931 8428 2977
rect 8602 2931 8613 2977
rect 8697 2931 8708 2977
rect 8882 2931 8893 2977
rect 8966 2931 8988 2977
rect 9162 2931 9268 2977
rect 9442 2931 9453 2977
rect 9537 2931 9548 2977
rect 9722 2971 10069 2977
rect 9722 2931 10006 2971
rect -39 2873 41 2925
rect -39 2827 -22 2873
rect 24 2827 41 2873
rect -39 2775 41 2827
rect -39 2729 -22 2775
rect 24 2729 41 2775
rect -39 2677 41 2729
rect -39 2631 -22 2677
rect 24 2631 41 2677
rect 369 2645 438 2931
rect 588 2645 669 2931
rect 1192 2779 1249 2931
rect 1695 2916 1709 2931
rect 1765 2916 1819 2931
rect 1875 2916 1895 2931
rect 1695 2904 1895 2916
rect 2052 2875 2102 2931
rect 3448 2875 3498 2931
rect 3655 2916 3675 2931
rect 3731 2916 3785 2931
rect 3841 2916 3855 2931
rect 3655 2904 3855 2916
rect 2052 2825 3498 2875
rect 4301 2779 4358 2931
rect 1192 2722 4358 2779
rect 5672 2779 5729 2931
rect 6175 2916 6189 2931
rect 6245 2916 6299 2931
rect 6355 2916 6375 2931
rect 6175 2904 6375 2916
rect 6532 2875 6582 2931
rect 7928 2875 7978 2931
rect 8135 2916 8155 2931
rect 8211 2916 8265 2931
rect 8321 2916 8335 2931
rect 8135 2904 8335 2916
rect 6532 2825 7978 2875
rect 8781 2779 8838 2931
rect 9720 2926 10006 2931
rect 5672 2722 8838 2779
rect 9989 2925 10006 2926
rect 10052 2925 10069 2971
rect 9989 2873 10069 2925
rect 9989 2827 10006 2873
rect 10052 2827 10069 2873
rect 9989 2775 10069 2827
rect 9989 2729 10006 2775
rect 10052 2729 10069 2775
rect 9989 2677 10069 2729
rect 855 2657 1055 2671
rect -39 2579 41 2631
rect 297 2599 308 2645
rect 482 2599 493 2645
rect 577 2599 588 2645
rect 762 2599 773 2645
rect 855 2601 867 2657
rect 923 2645 975 2657
rect 1031 2645 1055 2657
rect 1415 2664 1615 2672
rect 855 2599 868 2601
rect 1042 2599 1055 2645
rect 1137 2599 1148 2645
rect 1322 2599 1333 2645
rect 1415 2599 1428 2664
rect 1484 2645 1538 2664
rect 1594 2645 1615 2664
rect 1602 2599 1615 2645
rect -39 2533 -22 2579
rect 24 2533 41 2579
rect -39 2481 41 2533
rect -39 2435 -22 2481
rect 24 2435 41 2481
rect 333 2538 530 2543
rect 333 2482 349 2538
rect 405 2482 459 2538
rect 515 2533 530 2538
rect 588 2533 634 2599
rect 855 2594 1055 2599
rect 515 2487 634 2533
rect 515 2482 530 2487
rect 333 2477 530 2482
rect -39 2383 41 2435
rect -234 2323 -168 2338
rect -234 2267 -229 2323
rect -173 2267 -168 2323
rect -234 2213 -168 2267
rect -234 2157 -229 2213
rect -173 2157 -168 2213
rect -234 2141 -168 2157
rect -39 2337 -22 2383
rect 24 2337 41 2383
rect -39 2334 41 2337
rect 714 2471 1029 2475
rect 714 2415 851 2471
rect 907 2415 961 2471
rect 1017 2415 1029 2471
rect 714 2409 1029 2415
rect 1155 2428 1201 2599
rect 1415 2595 1615 2599
rect 1695 2661 1895 2672
rect 1695 2645 1709 2661
rect 1765 2645 1819 2661
rect 1875 2645 1895 2661
rect 2255 2658 2455 2672
rect 1695 2599 1708 2645
rect 1882 2599 1895 2645
rect 1977 2599 1988 2645
rect 2162 2599 2173 2645
rect 2255 2602 2267 2658
rect 2323 2645 2377 2658
rect 2433 2645 2455 2658
rect 3095 2658 3295 2672
rect 3095 2645 3117 2658
rect 3173 2645 3227 2658
rect 2255 2599 2268 2602
rect 2442 2599 2455 2645
rect 2537 2599 2548 2645
rect 2722 2599 2828 2645
rect 3002 2599 3013 2645
rect 3095 2599 3108 2645
rect 3283 2602 3295 2658
rect 3655 2661 3855 2672
rect 3655 2645 3675 2661
rect 3731 2645 3785 2661
rect 3841 2645 3855 2661
rect 3282 2599 3295 2602
rect 3377 2599 3388 2645
rect 3562 2599 3573 2645
rect 3655 2599 3668 2645
rect 3842 2599 3855 2645
rect 1695 2595 1895 2599
rect 1250 2537 1442 2539
rect 1988 2537 2038 2599
rect 2255 2595 2455 2599
rect 3095 2595 3295 2599
rect 1250 2536 2038 2537
rect 1250 2480 1262 2536
rect 1318 2480 1372 2536
rect 1428 2491 2038 2536
rect 3512 2537 3562 2599
rect 3655 2595 3855 2599
rect 3935 2664 4135 2672
rect 3935 2645 3956 2664
rect 4012 2645 4066 2664
rect 3935 2599 3948 2645
rect 4122 2599 4135 2664
rect 4495 2657 4695 2671
rect 4495 2645 4519 2657
rect 4575 2645 4627 2657
rect 4217 2599 4228 2645
rect 4402 2599 4413 2645
rect 4495 2599 4508 2645
rect 4683 2601 4695 2657
rect 5335 2657 5535 2671
rect 4682 2599 4695 2601
rect 4777 2599 4788 2645
rect 4962 2599 4973 2645
rect 5057 2599 5068 2645
rect 5242 2599 5253 2645
rect 5335 2601 5347 2657
rect 5403 2645 5455 2657
rect 5511 2645 5535 2657
rect 5895 2664 6095 2672
rect 5335 2599 5348 2601
rect 5522 2599 5535 2645
rect 5617 2599 5628 2645
rect 5802 2599 5813 2645
rect 5895 2599 5908 2664
rect 5964 2645 6018 2664
rect 6074 2645 6095 2664
rect 6082 2599 6095 2645
rect 3935 2595 4135 2599
rect 4108 2537 4300 2539
rect 3512 2536 4300 2537
rect 3512 2491 4122 2536
rect 1428 2480 1442 2491
rect 1250 2477 1442 2480
rect 4108 2480 4122 2491
rect 4178 2480 4232 2536
rect 4288 2480 4300 2536
rect 4108 2477 4300 2480
rect 4349 2428 4395 2599
rect 4495 2594 4695 2599
rect 4916 2553 4962 2599
rect 5068 2553 5114 2599
rect 5335 2594 5535 2599
rect 4884 2507 5114 2553
rect -39 2325 348 2334
rect 714 2325 762 2409
rect 1155 2382 2038 2428
rect 855 2325 1055 2327
rect -39 2285 308 2325
rect -39 2239 -22 2285
rect 24 2279 308 2285
rect 482 2279 493 2325
rect 577 2279 588 2325
rect 762 2279 773 2325
rect 855 2279 868 2325
rect 1042 2279 1055 2325
rect 24 2268 348 2279
rect 24 2239 41 2268
rect 855 2259 870 2279
rect 926 2259 980 2279
rect 1036 2259 1055 2279
rect 855 2249 1055 2259
rect 1135 2325 1335 2329
rect 1491 2325 1541 2326
rect 1775 2325 1825 2326
rect 1988 2325 2038 2382
rect 3512 2382 4395 2428
rect 4519 2470 4836 2475
rect 4519 2414 4531 2470
rect 4587 2414 4641 2470
rect 4697 2414 4836 2470
rect 4519 2409 4836 2414
rect 2255 2325 2455 2328
rect 1135 2279 1148 2325
rect 1322 2279 1335 2325
rect 1417 2279 1428 2325
rect 1602 2279 1613 2325
rect 1697 2279 1708 2325
rect 1882 2279 1893 2325
rect 1977 2279 1988 2325
rect 2162 2279 2173 2325
rect 2255 2279 2268 2325
rect 2442 2279 2455 2325
rect 1135 2265 1150 2279
rect 1206 2265 1260 2279
rect 1316 2265 1335 2279
rect 1135 2252 1335 2265
rect -39 2187 41 2239
rect -39 2141 -22 2187
rect 24 2141 41 2187
rect 96 2203 293 2207
rect 1491 2203 1541 2279
rect 96 2202 1541 2203
rect 96 2146 109 2202
rect 165 2146 219 2202
rect 275 2153 1541 2202
rect 1775 2201 1825 2279
rect 2255 2258 2269 2279
rect 2325 2258 2379 2279
rect 2435 2258 2455 2279
rect 2255 2248 2455 2258
rect 2535 2325 2735 2329
rect 2535 2260 2548 2325
rect 2722 2279 2735 2325
rect 2604 2260 2658 2279
rect 2714 2260 2735 2279
rect 2535 2252 2735 2260
rect 2815 2325 3015 2329
rect 2815 2279 2828 2325
rect 2815 2260 2836 2279
rect 2892 2260 2946 2279
rect 3002 2260 3015 2325
rect 2815 2252 3015 2260
rect 3095 2325 3295 2328
rect 3512 2325 3562 2382
rect 3725 2325 3775 2326
rect 4009 2325 4059 2326
rect 4215 2325 4415 2329
rect 3095 2279 3108 2325
rect 3282 2279 3295 2325
rect 3377 2279 3388 2325
rect 3562 2279 3573 2325
rect 3657 2279 3668 2325
rect 3842 2279 3853 2325
rect 3937 2279 3948 2325
rect 4122 2279 4133 2325
rect 4215 2279 4228 2325
rect 4402 2279 4415 2325
rect 3095 2258 3115 2279
rect 3171 2258 3225 2279
rect 3281 2258 3295 2279
rect 3095 2248 3295 2258
rect 3725 2201 3775 2279
rect 275 2146 293 2153
rect 1775 2151 3775 2201
rect 4009 2203 4059 2279
rect 4215 2265 4234 2279
rect 4290 2265 4344 2279
rect 4400 2265 4415 2279
rect 4215 2252 4415 2265
rect 4495 2325 4695 2327
rect 4788 2325 4836 2409
rect 5194 2471 5509 2475
rect 5194 2415 5331 2471
rect 5387 2415 5441 2471
rect 5497 2415 5509 2471
rect 5194 2409 5509 2415
rect 5635 2428 5681 2599
rect 5895 2595 6095 2599
rect 6175 2661 6375 2672
rect 6175 2645 6189 2661
rect 6245 2645 6299 2661
rect 6355 2645 6375 2661
rect 6735 2658 6935 2672
rect 6175 2599 6188 2645
rect 6362 2599 6375 2645
rect 6457 2599 6468 2645
rect 6642 2599 6653 2645
rect 6735 2602 6747 2658
rect 6803 2645 6857 2658
rect 6913 2645 6935 2658
rect 7575 2658 7775 2672
rect 7575 2645 7597 2658
rect 7653 2645 7707 2658
rect 6735 2599 6748 2602
rect 6922 2599 6935 2645
rect 7017 2599 7028 2645
rect 7202 2599 7308 2645
rect 7482 2599 7493 2645
rect 7575 2599 7588 2645
rect 7763 2602 7775 2658
rect 8135 2661 8335 2672
rect 8135 2645 8155 2661
rect 8211 2645 8265 2661
rect 8321 2645 8335 2661
rect 7762 2599 7775 2602
rect 7857 2599 7868 2645
rect 8042 2599 8053 2645
rect 8135 2599 8148 2645
rect 8322 2599 8335 2645
rect 6175 2595 6375 2599
rect 5730 2537 5922 2539
rect 6468 2537 6518 2599
rect 6735 2595 6935 2599
rect 7575 2595 7775 2599
rect 5730 2536 6518 2537
rect 5730 2480 5742 2536
rect 5798 2480 5852 2536
rect 5908 2491 6518 2536
rect 7992 2537 8042 2599
rect 8135 2595 8335 2599
rect 8415 2664 8615 2672
rect 8415 2645 8436 2664
rect 8492 2645 8546 2664
rect 8415 2599 8428 2645
rect 8602 2599 8615 2664
rect 8975 2657 9175 2671
rect 9989 2657 10006 2677
rect 8975 2645 8999 2657
rect 9055 2645 9107 2657
rect 8697 2599 8708 2645
rect 8882 2599 8893 2645
rect 8975 2599 8988 2645
rect 9163 2601 9175 2657
rect 9720 2645 10006 2657
rect 9162 2599 9175 2601
rect 9257 2599 9268 2645
rect 9442 2599 9453 2645
rect 9537 2599 9548 2645
rect 9722 2631 10006 2645
rect 10052 2631 10069 2677
rect 9722 2600 10069 2631
rect 9722 2599 9733 2600
rect 8415 2595 8615 2599
rect 8588 2537 8780 2539
rect 7992 2536 8780 2537
rect 7992 2491 8602 2536
rect 5908 2480 5922 2491
rect 5730 2477 5922 2480
rect 8588 2480 8602 2491
rect 8658 2480 8712 2536
rect 8768 2480 8780 2536
rect 8588 2477 8780 2480
rect 8829 2428 8875 2599
rect 8975 2594 9175 2599
rect 9396 2533 9442 2599
rect 9989 2579 10069 2600
rect 9700 2538 9897 2543
rect 9700 2533 9713 2538
rect 9396 2487 9713 2533
rect 9700 2482 9713 2487
rect 9771 2482 9823 2538
rect 9881 2482 9897 2538
rect 9700 2477 9897 2482
rect 9989 2533 10006 2579
rect 10052 2533 10069 2579
rect 9989 2481 10069 2533
rect 5194 2325 5242 2409
rect 5635 2382 6518 2428
rect 5335 2325 5535 2327
rect 4495 2279 4508 2325
rect 4682 2279 4695 2325
rect 4777 2279 4788 2325
rect 4962 2279 4973 2325
rect 5057 2279 5068 2325
rect 5242 2279 5253 2325
rect 5335 2279 5348 2325
rect 5522 2279 5535 2325
rect 4495 2259 4514 2279
rect 4570 2259 4624 2279
rect 4680 2259 4695 2279
rect 4495 2249 4695 2259
rect 5335 2259 5350 2279
rect 5406 2259 5460 2279
rect 5516 2259 5535 2279
rect 5335 2249 5535 2259
rect 5615 2325 5815 2329
rect 5971 2325 6021 2326
rect 6255 2325 6305 2326
rect 6468 2325 6518 2382
rect 7992 2382 8875 2428
rect 8999 2470 9316 2475
rect 8999 2414 9011 2470
rect 9067 2414 9121 2470
rect 9177 2414 9316 2470
rect 8999 2409 9316 2414
rect 6735 2325 6935 2328
rect 5615 2279 5628 2325
rect 5802 2279 5815 2325
rect 5897 2279 5908 2325
rect 6082 2279 6093 2325
rect 6177 2279 6188 2325
rect 6362 2279 6373 2325
rect 6457 2279 6468 2325
rect 6642 2279 6653 2325
rect 6735 2279 6748 2325
rect 6922 2279 6935 2325
rect 5615 2265 5630 2279
rect 5686 2265 5740 2279
rect 5796 2265 5815 2279
rect 5615 2252 5815 2265
rect 5971 2203 6021 2279
rect 4009 2153 6021 2203
rect 6255 2201 6305 2279
rect 6735 2258 6749 2279
rect 6805 2258 6859 2279
rect 6915 2258 6935 2279
rect 6735 2248 6935 2258
rect 7015 2325 7215 2329
rect 7015 2260 7028 2325
rect 7202 2279 7215 2325
rect 7084 2260 7138 2279
rect 7194 2260 7215 2279
rect 7015 2252 7215 2260
rect 7295 2325 7495 2329
rect 7295 2279 7308 2325
rect 7295 2260 7316 2279
rect 7372 2260 7426 2279
rect 7482 2260 7495 2325
rect 7295 2252 7495 2260
rect 7575 2325 7775 2328
rect 7992 2325 8042 2382
rect 8205 2325 8255 2326
rect 8489 2325 8539 2326
rect 8695 2325 8895 2329
rect 7575 2279 7588 2325
rect 7762 2279 7775 2325
rect 7857 2279 7868 2325
rect 8042 2279 8053 2325
rect 8137 2279 8148 2325
rect 8322 2279 8333 2325
rect 8417 2279 8428 2325
rect 8602 2279 8613 2325
rect 8695 2279 8708 2325
rect 8882 2279 8895 2325
rect 7575 2258 7595 2279
rect 7651 2258 7705 2279
rect 7761 2258 7775 2279
rect 7575 2248 7775 2258
rect 8205 2201 8255 2279
rect 6255 2151 8255 2201
rect 8489 2203 8539 2279
rect 8695 2265 8714 2279
rect 8770 2265 8824 2279
rect 8880 2265 8895 2279
rect 8695 2252 8895 2265
rect 8975 2325 9175 2327
rect 9268 2325 9316 2409
rect 9989 2435 10006 2481
rect 10052 2435 10069 2481
rect 9989 2383 10069 2435
rect 9989 2337 10006 2383
rect 10052 2337 10069 2383
rect 10122 2338 10185 4479
rect 9989 2334 10069 2337
rect 9718 2325 10069 2334
rect 8975 2279 8988 2325
rect 9162 2279 9175 2325
rect 9257 2279 9268 2325
rect 9442 2279 9453 2325
rect 9537 2279 9548 2325
rect 9722 2285 10069 2325
rect 9722 2279 10006 2285
rect 8975 2259 8994 2279
rect 9050 2259 9104 2279
rect 9160 2259 9175 2279
rect 9718 2277 10006 2279
rect 8975 2249 9175 2259
rect 9989 2239 10006 2277
rect 10052 2239 10069 2285
rect 9485 2203 9682 2207
rect 8489 2202 9682 2203
rect 8489 2153 9503 2202
rect 96 2141 293 2146
rect -39 2089 41 2141
rect -39 2043 -22 2089
rect 24 2043 41 2089
rect -346 2018 -280 2033
rect -346 1962 -341 2018
rect -285 1962 -280 2018
rect -469 1896 -403 1911
rect -469 1840 -464 1896
rect -408 1840 -403 1896
rect -469 1786 -403 1840
rect -346 1908 -280 1962
rect -346 1852 -341 1908
rect -285 1852 -280 1908
rect -346 1836 -280 1852
rect -39 2014 41 2043
rect -39 1993 349 2014
rect 855 2009 1055 2019
rect -39 1991 308 1993
rect -39 1945 -22 1991
rect 24 1948 308 1991
rect 24 1945 41 1948
rect 297 1947 308 1948
rect 482 1947 493 1993
rect 577 1947 588 1993
rect 762 1947 773 1993
rect 855 1947 868 2009
rect 924 1993 978 2009
rect 1034 1993 1055 2009
rect 1042 1947 1055 1993
rect -39 1893 41 1945
rect -39 1847 -22 1893
rect 24 1847 41 1893
rect -469 1730 -464 1786
rect -408 1730 -403 1786
rect -469 1714 -403 1730
rect -39 1795 41 1847
rect 87 1897 284 1902
rect 87 1841 100 1897
rect 156 1841 210 1897
rect 266 1894 284 1897
rect 588 1894 634 1947
rect 855 1942 1055 1947
rect 1135 2010 1335 2020
rect 1135 1947 1148 2010
rect 1204 1993 1258 2010
rect 1314 1993 1335 2010
rect 2255 2008 2455 2020
rect 1987 1993 2037 1994
rect 2255 1993 2270 2008
rect 2326 1993 2380 2008
rect 2436 1993 2455 2008
rect 1322 1947 1335 1993
rect 1417 1947 1428 1993
rect 1602 1947 1708 1993
rect 1882 1947 1893 1993
rect 1977 1947 1988 1993
rect 2162 1947 2173 1993
rect 2255 1947 2268 1993
rect 2442 1947 2455 1993
rect 2537 2008 2734 2013
rect 2537 1993 2553 2008
rect 2609 1993 2663 2008
rect 2719 1993 2734 2008
rect 2817 2008 3014 2013
rect 2817 1993 2833 2008
rect 2889 1993 2943 2008
rect 2999 1993 3014 2008
rect 2537 1947 2548 1993
rect 2722 1947 2828 1993
rect 3002 1947 3014 1993
rect 3095 2008 3295 2020
rect 3095 1993 3114 2008
rect 3170 1993 3224 2008
rect 3280 1993 3295 2008
rect 4215 2010 4415 2020
rect 3513 1993 3563 1994
rect 4215 1993 4236 2010
rect 4292 1993 4346 2010
rect 3095 1947 3108 1993
rect 3282 1947 3295 1993
rect 3377 1947 3388 1993
rect 3562 1947 3573 1993
rect 3657 1947 3668 1993
rect 3842 1947 3948 1993
rect 4122 1947 4133 1993
rect 4215 1947 4228 1993
rect 4402 1947 4415 2010
rect 1135 1943 1335 1947
rect 266 1848 634 1894
rect 1987 1891 2037 1947
rect 2255 1942 2455 1947
rect 3095 1942 3295 1947
rect 266 1841 284 1848
rect 87 1836 284 1841
rect 1154 1845 2037 1891
rect 3513 1891 3563 1947
rect 4215 1943 4415 1947
rect 4495 2009 4695 2019
rect 4495 1993 4516 2009
rect 4572 1993 4626 2009
rect 4495 1947 4508 1993
rect 4682 1947 4695 2009
rect 5335 2009 5535 2019
rect 4777 1947 4788 1993
rect 4962 1947 4973 1993
rect 5057 1947 5068 1993
rect 5242 1947 5253 1993
rect 5335 1947 5348 2009
rect 5404 1993 5458 2009
rect 5514 1993 5535 2009
rect 5522 1947 5535 1993
rect 4495 1942 4695 1947
rect 4916 1901 4962 1947
rect 5068 1901 5114 1947
rect 5335 1942 5535 1947
rect 5615 2010 5815 2020
rect 5615 1947 5628 2010
rect 5684 1993 5738 2010
rect 5794 1993 5815 2010
rect 6735 2008 6935 2020
rect 6467 1993 6517 1994
rect 6735 1993 6750 2008
rect 6806 1993 6860 2008
rect 6916 1993 6935 2008
rect 7575 2008 7775 2020
rect 7575 1993 7594 2008
rect 7650 1993 7704 2008
rect 7760 1993 7775 2008
rect 8695 2010 8895 2020
rect 7993 1993 8043 1994
rect 8695 1993 8716 2010
rect 8772 1993 8826 2010
rect 5802 1947 5815 1993
rect 5897 1947 5908 1993
rect 6082 1947 6188 1993
rect 6362 1947 6373 1993
rect 6457 1947 6468 1993
rect 6642 1947 6653 1993
rect 6735 1947 6748 1993
rect 6922 1947 6935 1993
rect 7017 1947 7028 1993
rect 7202 1947 7308 1993
rect 7482 1947 7493 1993
rect 7575 1947 7588 1993
rect 7762 1947 7775 1993
rect 7857 1947 7868 1993
rect 8042 1947 8053 1993
rect 8137 1947 8148 1993
rect 8322 1947 8428 1993
rect 8602 1947 8613 1993
rect 8695 1947 8708 1993
rect 8882 1947 8895 2010
rect 5615 1943 5815 1947
rect 3513 1845 4396 1891
rect 4884 1855 5114 1901
rect 6467 1891 6517 1947
rect 6735 1942 6935 1947
rect 7575 1942 7775 1947
rect -39 1749 -22 1795
rect 24 1749 41 1795
rect -39 1697 41 1749
rect 350 1780 547 1785
rect 350 1724 366 1780
rect 422 1724 476 1780
rect 532 1765 547 1780
rect 532 1724 634 1765
rect 350 1719 634 1724
rect -39 1651 -22 1697
rect 24 1674 41 1697
rect 24 1673 313 1674
rect 588 1673 634 1719
rect 855 1673 1055 1677
rect 1154 1673 1200 1845
rect 1249 1781 1329 1786
rect 1249 1725 1261 1781
rect 1317 1775 1329 1781
rect 4221 1781 4301 1786
rect 4221 1775 4233 1781
rect 1317 1729 2038 1775
rect 1317 1725 1329 1729
rect 1249 1719 1329 1725
rect 1415 1673 1615 1677
rect 24 1651 308 1673
rect -39 1627 308 1651
rect 482 1627 493 1673
rect 577 1627 588 1673
rect 762 1627 773 1673
rect -39 1599 41 1627
rect 855 1611 868 1673
rect 1042 1627 1055 1673
rect 1137 1627 1148 1673
rect 1322 1627 1333 1673
rect 1415 1627 1428 1673
rect 1602 1627 1615 1673
rect 924 1611 978 1627
rect 1034 1611 1055 1627
rect 855 1600 1055 1611
rect 1415 1610 1429 1627
rect 1485 1610 1539 1627
rect 1595 1610 1615 1627
rect 1415 1600 1615 1610
rect 1695 1673 1895 1677
rect 1988 1673 2038 1729
rect 3512 1729 4233 1775
rect 3512 1673 3562 1729
rect 4221 1725 4233 1729
rect 4289 1725 4301 1781
rect 4221 1719 4301 1725
rect 3655 1673 3855 1677
rect 1695 1627 1708 1673
rect 1882 1627 1895 1673
rect 1977 1627 1988 1673
rect 2162 1627 2173 1673
rect 2257 1627 2268 1673
rect 2442 1627 2548 1673
rect 2722 1627 2733 1673
rect 2817 1627 2828 1673
rect 3002 1627 3108 1673
rect 3282 1627 3293 1673
rect 3377 1627 3388 1673
rect 3562 1627 3573 1673
rect 3655 1627 3668 1673
rect 3842 1627 3855 1673
rect 1695 1611 1710 1627
rect 1766 1611 1820 1627
rect 1876 1611 1895 1627
rect 1695 1600 1895 1611
rect 3655 1611 3674 1627
rect 3730 1611 3784 1627
rect 3840 1611 3855 1627
rect 3655 1600 3855 1611
rect 3935 1673 4135 1677
rect 4350 1673 4396 1845
rect 5634 1845 6517 1891
rect 7993 1891 8043 1947
rect 8695 1943 8895 1947
rect 8975 2009 9175 2019
rect 8975 1993 8996 2009
rect 9052 1993 9106 2009
rect 8975 1947 8988 1993
rect 9162 1947 9175 2009
rect 9268 1993 9326 2153
rect 9485 2146 9503 2153
rect 9559 2146 9613 2202
rect 9669 2146 9682 2202
rect 9485 2141 9682 2146
rect 9989 2187 10069 2239
rect 9989 2141 10006 2187
rect 10052 2141 10069 2187
rect 9989 2089 10069 2141
rect 10121 2323 10185 2338
rect 10121 2267 10126 2323
rect 10182 2267 10185 2323
rect 10121 2213 10185 2267
rect 10121 2157 10126 2213
rect 10182 2212 10185 2213
rect 10231 4106 10297 4121
rect 10231 4050 10236 4106
rect 10292 4050 10297 4106
rect 10231 3996 10297 4050
rect 10231 3940 10236 3996
rect 10292 3940 10297 3996
rect 10231 3924 10297 3940
rect 10182 2157 10184 2212
rect 10121 2140 10184 2157
rect 9989 2043 10006 2089
rect 10052 2043 10069 2089
rect 9989 1996 10069 2043
rect 9717 1993 10069 1996
rect 9257 1947 9268 1993
rect 9442 1947 9453 1993
rect 9537 1947 9548 1993
rect 9722 1991 10069 1993
rect 9722 1947 10006 1991
rect 8975 1942 9175 1947
rect 9717 1945 10006 1947
rect 10052 1945 10069 1991
rect 9717 1939 10069 1945
rect 9989 1893 10069 1939
rect 7993 1845 8876 1891
rect 4884 1719 5114 1765
rect 4495 1673 4695 1677
rect 4916 1673 4962 1719
rect 5068 1673 5114 1719
rect 5335 1673 5535 1677
rect 5634 1673 5680 1845
rect 5729 1781 5809 1786
rect 5729 1725 5741 1781
rect 5797 1775 5809 1781
rect 8701 1781 8781 1786
rect 8701 1775 8713 1781
rect 5797 1729 6518 1775
rect 5797 1725 5809 1729
rect 5729 1719 5809 1725
rect 5895 1673 6095 1677
rect 3935 1627 3948 1673
rect 4122 1627 4135 1673
rect 4217 1627 4228 1673
rect 4402 1627 4413 1673
rect 4495 1627 4508 1673
rect 3935 1610 3955 1627
rect 4011 1610 4065 1627
rect 4121 1610 4135 1627
rect 3935 1600 4135 1610
rect 4495 1611 4516 1627
rect 4572 1611 4626 1627
rect 4682 1611 4695 1673
rect 4777 1627 4788 1673
rect 4962 1627 4973 1673
rect 5057 1627 5068 1673
rect 5242 1627 5253 1673
rect 4495 1600 4695 1611
rect 5335 1611 5348 1673
rect 5522 1627 5535 1673
rect 5617 1627 5628 1673
rect 5802 1627 5813 1673
rect 5895 1627 5908 1673
rect 6082 1627 6095 1673
rect 5404 1611 5458 1627
rect 5514 1611 5535 1627
rect 5335 1600 5535 1611
rect 5895 1610 5909 1627
rect 5965 1610 6019 1627
rect 6075 1610 6095 1627
rect 5895 1600 6095 1610
rect 6175 1673 6375 1677
rect 6468 1673 6518 1729
rect 7992 1729 8713 1775
rect 7992 1673 8042 1729
rect 8701 1725 8713 1729
rect 8769 1725 8781 1781
rect 8701 1719 8781 1725
rect 8135 1673 8335 1677
rect 6175 1627 6188 1673
rect 6362 1627 6375 1673
rect 6457 1627 6468 1673
rect 6642 1627 6653 1673
rect 6737 1627 6748 1673
rect 6922 1627 7028 1673
rect 7202 1627 7213 1673
rect 7297 1627 7308 1673
rect 7482 1627 7588 1673
rect 7762 1627 7773 1673
rect 7857 1627 7868 1673
rect 8042 1627 8053 1673
rect 8135 1627 8148 1673
rect 8322 1627 8335 1673
rect 6175 1611 6190 1627
rect 6246 1611 6300 1627
rect 6356 1611 6375 1627
rect 6175 1600 6375 1611
rect 8135 1611 8154 1627
rect 8210 1611 8264 1627
rect 8320 1611 8335 1627
rect 8135 1600 8335 1611
rect 8415 1673 8615 1677
rect 8830 1673 8876 1845
rect 9989 1847 10006 1893
rect 10052 1847 10069 1893
rect 9989 1795 10069 1847
rect 9484 1780 9681 1785
rect 9484 1766 9502 1780
rect 9442 1765 9502 1766
rect 9396 1724 9502 1765
rect 9558 1724 9612 1780
rect 9668 1724 9681 1780
rect 9396 1719 9681 1724
rect 9989 1749 10006 1795
rect 10052 1749 10069 1795
rect 8975 1673 9175 1677
rect 9396 1673 9442 1719
rect 9989 1697 10069 1749
rect 9989 1678 10006 1697
rect 8415 1627 8428 1673
rect 8602 1627 8615 1673
rect 8697 1627 8708 1673
rect 8882 1627 8893 1673
rect 8975 1627 8988 1673
rect 8415 1610 8435 1627
rect 8491 1610 8545 1627
rect 8601 1610 8615 1627
rect 8415 1600 8615 1610
rect 8975 1611 8996 1627
rect 9052 1611 9106 1627
rect 9162 1611 9175 1673
rect 9257 1627 9268 1673
rect 9442 1627 9453 1673
rect 9537 1627 9548 1673
rect 9722 1651 10006 1678
rect 10052 1651 10069 1697
rect 9722 1621 10069 1651
rect 8975 1600 9175 1611
rect -39 1553 -22 1599
rect 24 1553 41 1599
rect 9989 1599 10069 1621
rect -39 1501 41 1553
rect -39 1455 -22 1501
rect 24 1455 41 1501
rect 88 1556 285 1561
rect 88 1500 101 1556
rect 157 1500 211 1556
rect 267 1554 285 1556
rect 9733 1556 9935 1561
rect 9733 1554 9751 1556
rect 267 1504 2038 1554
rect 267 1500 285 1504
rect 88 1495 285 1500
rect -39 1403 41 1455
rect -39 1357 -22 1403
rect 24 1357 41 1403
rect -39 1348 41 1357
rect 857 1364 1054 1369
rect -39 1341 327 1348
rect 857 1341 870 1364
rect 926 1341 980 1364
rect 1036 1341 1054 1364
rect 1415 1367 1612 1372
rect -580 1304 -514 1319
rect -580 1248 -575 1304
rect -519 1248 -514 1304
rect -580 1194 -514 1248
rect -580 1138 -575 1194
rect -519 1138 -514 1194
rect -580 1122 -514 1138
rect -39 1305 308 1341
rect -39 1259 -22 1305
rect 24 1295 308 1305
rect 482 1295 493 1341
rect 577 1295 588 1341
rect 762 1295 868 1341
rect 1042 1303 1054 1341
rect 1042 1295 1053 1303
rect 1137 1295 1148 1341
rect 1322 1295 1333 1341
rect 1415 1306 1428 1367
rect 1484 1341 1538 1367
rect 1594 1341 1612 1367
rect 1988 1341 2038 1504
rect 3512 1504 6518 1554
rect 2255 1353 2455 1368
rect 1417 1295 1428 1306
rect 1602 1295 1613 1341
rect 1697 1295 1708 1341
rect 1882 1295 1893 1341
rect 1977 1295 1988 1341
rect 2162 1295 2173 1341
rect 2255 1297 2267 1353
rect 2323 1341 2377 1353
rect 2433 1341 2455 1353
rect 3095 1353 3295 1368
rect 3095 1341 3117 1353
rect 3173 1341 3227 1353
rect 2255 1295 2268 1297
rect 2442 1295 2455 1341
rect 2537 1295 2548 1341
rect 2722 1295 2828 1341
rect 3002 1295 3013 1341
rect 3095 1295 3108 1341
rect 3283 1297 3295 1353
rect 3512 1341 3562 1504
rect 4333 1393 5697 1443
rect 4333 1367 4402 1393
rect 4332 1341 4402 1367
rect 5628 1367 5697 1393
rect 5628 1341 5698 1367
rect 6468 1341 6518 1504
rect 7992 1504 9751 1554
rect 6735 1353 6935 1368
rect 3282 1295 3295 1297
rect 3377 1295 3388 1341
rect 3562 1295 3573 1341
rect 3657 1295 3668 1341
rect 3842 1295 3853 1341
rect 3937 1295 3948 1341
rect 4122 1295 4133 1341
rect 4217 1295 4228 1341
rect 4402 1295 4413 1341
rect 4497 1295 4508 1341
rect 4682 1295 4788 1341
rect 4962 1295 4973 1341
rect 5057 1295 5068 1341
rect 5242 1295 5348 1341
rect 5522 1295 5533 1341
rect 5617 1295 5628 1341
rect 5802 1295 5813 1341
rect 5897 1295 5908 1341
rect 6082 1295 6093 1341
rect 6177 1295 6188 1341
rect 6362 1295 6373 1341
rect 6457 1295 6468 1341
rect 6642 1295 6653 1341
rect 6735 1297 6747 1353
rect 6803 1341 6857 1353
rect 6913 1341 6935 1353
rect 7575 1353 7775 1368
rect 7575 1341 7597 1353
rect 7653 1341 7707 1353
rect 6735 1295 6748 1297
rect 6922 1295 6935 1341
rect 7017 1295 7028 1341
rect 7202 1295 7308 1341
rect 7482 1295 7493 1341
rect 7575 1295 7588 1341
rect 7763 1297 7775 1353
rect 7992 1341 8042 1504
rect 9733 1500 9751 1504
rect 9807 1500 9861 1556
rect 9917 1500 9935 1556
rect 9733 1495 9935 1500
rect 9989 1553 10006 1599
rect 10052 1553 10069 1599
rect 9989 1501 10069 1553
rect 9483 1453 9680 1458
rect 9483 1443 9501 1453
rect 8813 1397 9501 1443
rect 9557 1397 9611 1453
rect 9667 1397 9680 1453
rect 8813 1393 9680 1397
rect 8813 1367 8882 1393
rect 9483 1392 9680 1393
rect 9989 1455 10006 1501
rect 10052 1455 10069 1501
rect 10231 1678 10294 3924
rect 10231 1622 10236 1678
rect 10292 1622 10294 1678
rect 10231 1568 10294 1622
rect 10231 1512 10236 1568
rect 10292 1512 10294 1568
rect 10231 1495 10294 1512
rect 10360 3904 10423 3919
rect 10360 3848 10365 3904
rect 10421 3848 10423 3904
rect 10360 3794 10423 3848
rect 10360 3738 10365 3794
rect 10421 3738 10423 3794
rect 9989 1403 10069 1455
rect 8812 1341 8882 1367
rect 9989 1357 10006 1403
rect 10052 1357 10069 1403
rect 9989 1348 10069 1357
rect 9710 1341 10069 1348
rect 7762 1295 7775 1297
rect 7857 1295 7868 1341
rect 8042 1295 8053 1341
rect 8137 1295 8148 1341
rect 8322 1295 8333 1341
rect 8417 1295 8428 1341
rect 8602 1295 8613 1341
rect 8697 1295 8708 1341
rect 8882 1295 8893 1341
rect 8977 1295 8988 1341
rect 9162 1295 9268 1341
rect 9442 1295 9453 1341
rect 9537 1295 9548 1341
rect 9722 1305 10069 1341
rect 9722 1295 10006 1305
rect 24 1291 327 1295
rect 24 1259 41 1291
rect -39 1207 41 1259
rect -39 1161 -22 1207
rect 24 1161 41 1207
rect -39 1109 41 1161
rect 92 1183 289 1188
rect 92 1127 105 1183
rect 161 1127 215 1183
rect 271 1181 289 1183
rect 1232 1181 1322 1295
rect 1429 1181 1482 1295
rect 271 1128 1482 1181
rect 271 1127 289 1128
rect 92 1122 289 1127
rect 1429 1121 1482 1128
rect 1827 1176 1880 1295
rect 2255 1291 2455 1295
rect 3095 1291 3295 1295
rect 3670 1176 3723 1295
rect 1827 1123 3723 1176
rect 4068 1181 4121 1295
rect 5909 1181 5962 1295
rect 4068 1128 5962 1181
rect 4068 1121 4121 1128
rect 5909 1121 5962 1128
rect 6307 1176 6360 1295
rect 6735 1291 6935 1295
rect 7575 1291 7775 1295
rect 8150 1176 8203 1295
rect 6307 1123 8203 1176
rect 8548 1181 8601 1295
rect 9710 1291 10006 1295
rect 9989 1259 10006 1291
rect 10052 1259 10069 1305
rect 10360 1476 10423 3738
rect 10481 3733 10545 3748
rect 10481 3677 10484 3733
rect 10540 3677 10545 3733
rect 10481 3623 10545 3677
rect 10481 3617 10484 3623
rect 10360 1420 10365 1476
rect 10421 1420 10423 1476
rect 10360 1366 10423 1420
rect 10360 1310 10365 1366
rect 10421 1310 10423 1366
rect 10360 1293 10423 1310
rect 10479 3567 10484 3617
rect 10540 3567 10545 3623
rect 10479 3551 10545 3567
rect 10479 1305 10542 3551
rect 9989 1207 10069 1259
rect 9713 1183 9910 1188
rect 9713 1181 9731 1183
rect 8548 1128 9731 1181
rect 8548 1121 8601 1128
rect 9713 1127 9731 1128
rect 9787 1127 9841 1183
rect 9897 1127 9910 1183
rect 9713 1122 9910 1127
rect 9989 1161 10006 1207
rect 10052 1161 10069 1207
rect -39 1063 -22 1109
rect 24 1063 41 1109
rect -39 1028 41 1063
rect 9989 1109 10069 1161
rect 10479 1249 10484 1305
rect 10540 1249 10542 1305
rect 10479 1195 10542 1249
rect 10479 1139 10484 1195
rect 10540 1139 10542 1195
rect 10479 1122 10542 1139
rect 9989 1063 10006 1109
rect 10052 1063 10069 1109
rect 9989 1028 10069 1063
rect -39 1011 10069 1028
rect -39 965 -22 1011
rect 24 965 76 1011
rect 122 965 174 1011
rect 220 965 272 1011
rect 318 965 370 1011
rect 416 965 468 1011
rect 514 965 566 1011
rect 612 965 664 1011
rect 710 965 762 1011
rect 808 965 860 1011
rect 906 965 958 1011
rect 1004 965 1056 1011
rect 1102 965 1154 1011
rect 1200 965 1252 1011
rect 1298 965 1350 1011
rect 1396 965 1448 1011
rect 1494 965 1546 1011
rect 1592 965 1644 1011
rect 1690 965 1742 1011
rect 1788 965 1840 1011
rect 1886 965 1938 1011
rect 1984 965 2036 1011
rect 2082 965 2134 1011
rect 2180 965 2232 1011
rect 2278 965 2330 1011
rect 2376 965 2428 1011
rect 2474 965 2526 1011
rect 2572 965 2624 1011
rect 2670 965 2722 1011
rect 2768 965 2820 1011
rect 2866 965 2918 1011
rect 2964 965 3016 1011
rect 3062 965 3114 1011
rect 3160 965 3212 1011
rect 3258 965 3310 1011
rect 3356 965 3408 1011
rect 3454 965 3506 1011
rect 3552 965 3604 1011
rect 3650 965 3702 1011
rect 3748 965 3800 1011
rect 3846 965 3898 1011
rect 3944 965 3996 1011
rect 4042 965 4094 1011
rect 4140 965 4192 1011
rect 4238 965 4290 1011
rect 4336 965 4388 1011
rect 4434 965 4486 1011
rect 4532 965 4584 1011
rect 4630 965 4682 1011
rect 4728 965 4780 1011
rect 4826 965 4878 1011
rect 4924 965 4976 1011
rect 5022 965 5074 1011
rect 5120 965 5172 1011
rect 5218 965 5270 1011
rect 5316 965 5368 1011
rect 5414 965 5466 1011
rect 5512 965 5564 1011
rect 5610 965 5662 1011
rect 5708 965 5760 1011
rect 5806 965 5858 1011
rect 5904 965 5956 1011
rect 6002 965 6054 1011
rect 6100 965 6152 1011
rect 6198 965 6250 1011
rect 6296 965 6348 1011
rect 6394 965 6446 1011
rect 6492 965 6544 1011
rect 6590 965 6642 1011
rect 6688 965 6740 1011
rect 6786 965 6838 1011
rect 6884 965 6936 1011
rect 6982 965 7034 1011
rect 7080 965 7132 1011
rect 7178 965 7230 1011
rect 7276 965 7328 1011
rect 7374 965 7426 1011
rect 7472 965 7524 1011
rect 7570 965 7622 1011
rect 7668 965 7720 1011
rect 7766 965 7818 1011
rect 7864 965 7916 1011
rect 7962 965 8014 1011
rect 8060 965 8112 1011
rect 8158 965 8210 1011
rect 8256 965 8308 1011
rect 8354 965 8406 1011
rect 8452 965 8504 1011
rect 8550 965 8602 1011
rect 8648 965 8700 1011
rect 8746 965 8798 1011
rect 8844 965 8896 1011
rect 8942 965 8994 1011
rect 9040 965 9092 1011
rect 9138 965 9190 1011
rect 9236 965 9288 1011
rect 9334 965 9386 1011
rect 9432 965 9484 1011
rect 9530 965 9582 1011
rect 9628 965 9680 1011
rect 9726 965 9778 1011
rect 9824 965 9876 1011
rect 9922 965 10006 1011
rect 10052 965 10069 1011
rect -39 948 10069 965
<< via1 >>
rect 2466 5456 2522 5512
rect 2576 5456 2632 5512
rect 2918 5456 2974 5512
rect 3028 5456 3084 5512
rect 6946 5456 7002 5512
rect 7056 5456 7112 5512
rect 7398 5456 7454 5512
rect 7508 5456 7564 5512
rect 1709 5360 1765 5401
rect 1819 5360 1875 5401
rect 3675 5360 3731 5401
rect 3785 5360 3841 5401
rect 6189 5360 6245 5401
rect 6299 5360 6355 5401
rect 8155 5360 8211 5401
rect 8265 5360 8321 5401
rect 1709 5345 1765 5360
rect 1819 5345 1875 5360
rect 3675 5345 3731 5360
rect 3785 5345 3841 5360
rect 6189 5345 6245 5360
rect 6299 5345 6355 5360
rect 8155 5345 8211 5360
rect 8265 5345 8321 5360
rect 867 5074 923 5086
rect 975 5074 1031 5086
rect 867 5030 868 5074
rect 868 5030 923 5074
rect 975 5030 1031 5074
rect 1428 5074 1484 5093
rect 1538 5074 1594 5093
rect 1428 5037 1484 5074
rect 1538 5037 1594 5074
rect 349 4911 405 4967
rect 459 4911 515 4967
rect -231 4696 -175 4752
rect -231 4586 -175 4642
rect 851 4844 907 4900
rect 961 4844 1017 4900
rect 1709 5074 1765 5090
rect 1819 5074 1875 5090
rect 1709 5034 1765 5074
rect 1819 5034 1875 5074
rect 2267 5074 2323 5087
rect 2377 5074 2433 5087
rect 3117 5074 3173 5087
rect 3227 5074 3283 5087
rect 2267 5031 2268 5074
rect 2268 5031 2323 5074
rect 2377 5031 2433 5074
rect 3117 5031 3173 5074
rect 3227 5031 3282 5074
rect 3282 5031 3283 5074
rect 3675 5074 3731 5090
rect 3785 5074 3841 5090
rect 3675 5034 3731 5074
rect 3785 5034 3841 5074
rect 1262 4909 1318 4965
rect 1372 4909 1428 4965
rect 3956 5074 4012 5093
rect 4066 5074 4122 5093
rect 3956 5037 4012 5074
rect 4066 5037 4122 5074
rect 4519 5074 4575 5086
rect 4627 5074 4683 5086
rect 4519 5030 4575 5074
rect 4627 5030 4682 5074
rect 4682 5030 4683 5074
rect 5347 5074 5403 5086
rect 5455 5074 5511 5086
rect 5347 5030 5348 5074
rect 5348 5030 5403 5074
rect 5455 5030 5511 5074
rect 5908 5074 5964 5093
rect 6018 5074 6074 5093
rect 5908 5037 5964 5074
rect 6018 5037 6074 5074
rect 4122 4909 4178 4965
rect 4232 4909 4288 4965
rect 870 4708 926 4744
rect 980 4708 1036 4744
rect 870 4688 926 4708
rect 980 4688 1036 4708
rect 4531 4843 4587 4899
rect 4641 4843 4697 4899
rect 1150 4708 1206 4750
rect 1260 4708 1316 4750
rect 2269 4708 2325 4743
rect 2379 4708 2435 4743
rect 1150 4694 1206 4708
rect 1260 4694 1316 4708
rect 109 4575 165 4631
rect 219 4575 275 4631
rect 2269 4687 2325 4708
rect 2379 4687 2435 4708
rect 2548 4708 2604 4745
rect 2658 4708 2714 4745
rect 2548 4689 2604 4708
rect 2658 4689 2714 4708
rect 2836 4708 2892 4745
rect 2946 4708 3002 4745
rect 2836 4689 2892 4708
rect 2946 4689 3002 4708
rect 3115 4708 3171 4743
rect 3225 4708 3281 4743
rect 4234 4708 4290 4750
rect 4344 4708 4400 4750
rect 3115 4687 3171 4708
rect 3225 4687 3281 4708
rect 4234 4694 4290 4708
rect 4344 4694 4400 4708
rect 5331 4844 5387 4900
rect 5441 4844 5497 4900
rect 6189 5074 6245 5090
rect 6299 5074 6355 5090
rect 6189 5034 6245 5074
rect 6299 5034 6355 5074
rect 6747 5074 6803 5087
rect 6857 5074 6913 5087
rect 7597 5074 7653 5087
rect 7707 5074 7763 5087
rect 6747 5031 6748 5074
rect 6748 5031 6803 5074
rect 6857 5031 6913 5074
rect 7597 5031 7653 5074
rect 7707 5031 7762 5074
rect 7762 5031 7763 5074
rect 8155 5074 8211 5090
rect 8265 5074 8321 5090
rect 8155 5034 8211 5074
rect 8265 5034 8321 5074
rect 5742 4909 5798 4965
rect 5852 4909 5908 4965
rect 8436 5074 8492 5093
rect 8546 5074 8602 5093
rect 8436 5037 8492 5074
rect 8546 5037 8602 5074
rect 8999 5074 9055 5086
rect 9107 5074 9163 5086
rect 8999 5030 9055 5074
rect 9107 5030 9162 5074
rect 9162 5030 9163 5074
rect 8602 4909 8658 4965
rect 8712 4909 8768 4965
rect 9713 4911 9771 4967
rect 9823 4911 9881 4967
rect 4514 4708 4570 4744
rect 4624 4708 4680 4744
rect 5350 4708 5406 4744
rect 5460 4708 5516 4744
rect 4514 4688 4570 4708
rect 4624 4688 4680 4708
rect 5350 4688 5406 4708
rect 5460 4688 5516 4708
rect 9011 4843 9067 4899
rect 9121 4843 9177 4899
rect 5630 4708 5686 4750
rect 5740 4708 5796 4750
rect 6749 4708 6805 4743
rect 6859 4708 6915 4743
rect 5630 4694 5686 4708
rect 5740 4694 5796 4708
rect 6749 4687 6805 4708
rect 6859 4687 6915 4708
rect 7028 4708 7084 4745
rect 7138 4708 7194 4745
rect 7028 4689 7084 4708
rect 7138 4689 7194 4708
rect 7316 4708 7372 4745
rect 7426 4708 7482 4745
rect 7316 4689 7372 4708
rect 7426 4689 7482 4708
rect 7595 4708 7651 4743
rect 7705 4708 7761 4743
rect 8714 4708 8770 4750
rect 8824 4708 8880 4750
rect 7595 4687 7651 4708
rect 7705 4687 7761 4708
rect 8714 4694 8770 4708
rect 8824 4694 8880 4708
rect 8994 4708 9050 4744
rect 9104 4708 9160 4744
rect 8994 4688 9050 4708
rect 9104 4688 9160 4708
rect -341 4391 -285 4447
rect -463 4269 -407 4325
rect -463 4159 -407 4215
rect -341 4281 -285 4337
rect -577 3677 -521 3733
rect -577 3567 -521 3623
rect 868 4422 924 4438
rect 978 4422 1034 4438
rect 868 4382 924 4422
rect 978 4382 1034 4422
rect 100 4270 156 4326
rect 210 4270 266 4326
rect 1148 4422 1204 4439
rect 1258 4422 1314 4439
rect 2270 4422 2326 4437
rect 2380 4422 2436 4437
rect 1148 4383 1204 4422
rect 1258 4383 1314 4422
rect 2270 4381 2326 4422
rect 2380 4381 2436 4422
rect 2553 4422 2609 4437
rect 2663 4422 2719 4437
rect 2833 4422 2889 4437
rect 2943 4422 2999 4437
rect 2553 4381 2609 4422
rect 2663 4381 2719 4422
rect 2833 4381 2889 4422
rect 2943 4381 2999 4422
rect 3114 4422 3170 4437
rect 3224 4422 3280 4437
rect 4236 4422 4292 4439
rect 4346 4422 4402 4439
rect 3114 4381 3170 4422
rect 3224 4381 3280 4422
rect 4236 4383 4292 4422
rect 4346 4383 4402 4422
rect 4516 4422 4572 4438
rect 4626 4422 4682 4438
rect 4516 4382 4572 4422
rect 4626 4382 4682 4422
rect 5348 4422 5404 4438
rect 5458 4422 5514 4438
rect 5348 4382 5404 4422
rect 5458 4382 5514 4422
rect 5628 4422 5684 4439
rect 5738 4422 5794 4439
rect 6750 4422 6806 4437
rect 6860 4422 6916 4437
rect 7594 4422 7650 4437
rect 7704 4422 7760 4437
rect 8716 4422 8772 4439
rect 8826 4422 8882 4439
rect 5628 4383 5684 4422
rect 5738 4383 5794 4422
rect 6750 4381 6806 4422
rect 6860 4381 6916 4422
rect 7594 4381 7650 4422
rect 7704 4381 7760 4422
rect 8716 4383 8772 4422
rect 8826 4383 8882 4422
rect 366 4153 422 4209
rect 476 4153 532 4209
rect 1261 4154 1317 4210
rect 868 4056 924 4096
rect 978 4056 1034 4096
rect 1429 4056 1485 4095
rect 1539 4056 1595 4095
rect 868 4040 924 4056
rect 978 4040 1034 4056
rect 1429 4039 1485 4056
rect 1539 4039 1595 4056
rect 4233 4154 4289 4210
rect 1710 4056 1766 4096
rect 1820 4056 1876 4096
rect 3674 4056 3730 4096
rect 3784 4056 3840 4096
rect 1710 4040 1766 4056
rect 1820 4040 1876 4056
rect 3674 4040 3730 4056
rect 3784 4040 3840 4056
rect 8996 4422 9052 4438
rect 9106 4422 9162 4438
rect 8996 4382 9052 4422
rect 9106 4382 9162 4422
rect 9503 4575 9559 4631
rect 9613 4575 9669 4631
rect 5741 4154 5797 4210
rect 3955 4056 4011 4095
rect 4065 4056 4121 4095
rect 4516 4056 4572 4096
rect 4626 4056 4682 4096
rect 3955 4039 4011 4056
rect 4065 4039 4121 4056
rect 4516 4040 4572 4056
rect 4626 4040 4682 4056
rect 5348 4056 5404 4096
rect 5458 4056 5514 4096
rect 5909 4056 5965 4095
rect 6019 4056 6075 4095
rect 5348 4040 5404 4056
rect 5458 4040 5514 4056
rect 5909 4039 5965 4056
rect 6019 4039 6075 4056
rect 8713 4154 8769 4210
rect 6190 4056 6246 4096
rect 6300 4056 6356 4096
rect 8154 4056 8210 4096
rect 8264 4056 8320 4096
rect 6190 4040 6246 4056
rect 6300 4040 6356 4056
rect 8154 4040 8210 4056
rect 8264 4040 8320 4056
rect 9502 4153 9558 4209
rect 9612 4153 9668 4209
rect 8435 4056 8491 4095
rect 8545 4056 8601 4095
rect 8996 4056 9052 4096
rect 9106 4056 9162 4096
rect 8435 4039 8491 4056
rect 8545 4039 8601 4056
rect 8996 4040 9052 4056
rect 9106 4040 9162 4056
rect 101 3929 157 3985
rect 211 3929 267 3985
rect 870 3770 926 3793
rect 980 3770 1036 3793
rect 870 3737 926 3770
rect 980 3737 1036 3770
rect 1428 3770 1484 3795
rect 1538 3770 1594 3795
rect 1428 3739 1484 3770
rect 1538 3739 1594 3770
rect 2267 3770 2323 3782
rect 2377 3770 2433 3782
rect 3117 3770 3173 3782
rect 3227 3770 3283 3782
rect 2267 3726 2268 3770
rect 2268 3726 2323 3770
rect 2377 3726 2433 3770
rect 3117 3726 3173 3770
rect 3227 3726 3282 3770
rect 3282 3726 3283 3770
rect 6747 3770 6803 3782
rect 6857 3770 6913 3782
rect 7597 3770 7653 3782
rect 7707 3770 7763 3782
rect 6747 3726 6748 3770
rect 6748 3726 6803 3770
rect 6857 3726 6913 3770
rect 7597 3726 7653 3770
rect 7707 3726 7762 3770
rect 7762 3726 7763 3770
rect 9751 3929 9807 3985
rect 9861 3929 9917 3985
rect 9501 3826 9557 3882
rect 9611 3826 9667 3882
rect 105 3556 161 3612
rect 215 3556 271 3612
rect 9731 3556 9787 3612
rect 9841 3556 9897 3612
rect 10127 4589 10183 4645
rect 10127 4479 10183 4535
rect 2466 3027 2522 3083
rect 2576 3027 2632 3083
rect 2918 3027 2974 3083
rect 3028 3027 3084 3083
rect 6946 3027 7002 3083
rect 7056 3027 7112 3083
rect 7398 3027 7454 3083
rect 7508 3027 7564 3083
rect 1709 2931 1765 2972
rect 1819 2931 1875 2972
rect 3675 2931 3731 2972
rect 3785 2931 3841 2972
rect 6189 2931 6245 2972
rect 6299 2931 6355 2972
rect 8155 2931 8211 2972
rect 8265 2931 8321 2972
rect 1709 2916 1765 2931
rect 1819 2916 1875 2931
rect 3675 2916 3731 2931
rect 3785 2916 3841 2931
rect 6189 2916 6245 2931
rect 6299 2916 6355 2931
rect 8155 2916 8211 2931
rect 8265 2916 8321 2931
rect 867 2645 923 2657
rect 975 2645 1031 2657
rect 867 2601 868 2645
rect 868 2601 923 2645
rect 975 2601 1031 2645
rect 1428 2645 1484 2664
rect 1538 2645 1594 2664
rect 1428 2608 1484 2645
rect 1538 2608 1594 2645
rect 349 2482 405 2538
rect 459 2482 515 2538
rect -229 2267 -173 2323
rect -229 2157 -173 2213
rect 851 2415 907 2471
rect 961 2415 1017 2471
rect 1709 2645 1765 2661
rect 1819 2645 1875 2661
rect 1709 2605 1765 2645
rect 1819 2605 1875 2645
rect 2267 2645 2323 2658
rect 2377 2645 2433 2658
rect 3117 2645 3173 2658
rect 3227 2645 3283 2658
rect 2267 2602 2268 2645
rect 2268 2602 2323 2645
rect 2377 2602 2433 2645
rect 3117 2602 3173 2645
rect 3227 2602 3282 2645
rect 3282 2602 3283 2645
rect 3675 2645 3731 2661
rect 3785 2645 3841 2661
rect 3675 2605 3731 2645
rect 3785 2605 3841 2645
rect 1262 2480 1318 2536
rect 1372 2480 1428 2536
rect 3956 2645 4012 2664
rect 4066 2645 4122 2664
rect 3956 2608 4012 2645
rect 4066 2608 4122 2645
rect 4519 2645 4575 2657
rect 4627 2645 4683 2657
rect 4519 2601 4575 2645
rect 4627 2601 4682 2645
rect 4682 2601 4683 2645
rect 5347 2645 5403 2657
rect 5455 2645 5511 2657
rect 5347 2601 5348 2645
rect 5348 2601 5403 2645
rect 5455 2601 5511 2645
rect 5908 2645 5964 2664
rect 6018 2645 6074 2664
rect 5908 2608 5964 2645
rect 6018 2608 6074 2645
rect 4122 2480 4178 2536
rect 4232 2480 4288 2536
rect 870 2279 926 2315
rect 980 2279 1036 2315
rect 870 2259 926 2279
rect 980 2259 1036 2279
rect 4531 2414 4587 2470
rect 4641 2414 4697 2470
rect 1150 2279 1206 2321
rect 1260 2279 1316 2321
rect 2269 2279 2325 2314
rect 2379 2279 2435 2314
rect 1150 2265 1206 2279
rect 1260 2265 1316 2279
rect 109 2146 165 2202
rect 219 2146 275 2202
rect 2269 2258 2325 2279
rect 2379 2258 2435 2279
rect 2548 2279 2604 2316
rect 2658 2279 2714 2316
rect 2548 2260 2604 2279
rect 2658 2260 2714 2279
rect 2836 2279 2892 2316
rect 2946 2279 3002 2316
rect 2836 2260 2892 2279
rect 2946 2260 3002 2279
rect 3115 2279 3171 2314
rect 3225 2279 3281 2314
rect 4234 2279 4290 2321
rect 4344 2279 4400 2321
rect 3115 2258 3171 2279
rect 3225 2258 3281 2279
rect 4234 2265 4290 2279
rect 4344 2265 4400 2279
rect 5331 2415 5387 2471
rect 5441 2415 5497 2471
rect 6189 2645 6245 2661
rect 6299 2645 6355 2661
rect 6189 2605 6245 2645
rect 6299 2605 6355 2645
rect 6747 2645 6803 2658
rect 6857 2645 6913 2658
rect 7597 2645 7653 2658
rect 7707 2645 7763 2658
rect 6747 2602 6748 2645
rect 6748 2602 6803 2645
rect 6857 2602 6913 2645
rect 7597 2602 7653 2645
rect 7707 2602 7762 2645
rect 7762 2602 7763 2645
rect 8155 2645 8211 2661
rect 8265 2645 8321 2661
rect 8155 2605 8211 2645
rect 8265 2605 8321 2645
rect 5742 2480 5798 2536
rect 5852 2480 5908 2536
rect 8436 2645 8492 2664
rect 8546 2645 8602 2664
rect 8436 2608 8492 2645
rect 8546 2608 8602 2645
rect 8999 2645 9055 2657
rect 9107 2645 9163 2657
rect 8999 2601 9055 2645
rect 9107 2601 9162 2645
rect 9162 2601 9163 2645
rect 8602 2480 8658 2536
rect 8712 2480 8768 2536
rect 9713 2482 9771 2538
rect 9823 2482 9881 2538
rect 4514 2279 4570 2315
rect 4624 2279 4680 2315
rect 5350 2279 5406 2315
rect 5460 2279 5516 2315
rect 4514 2259 4570 2279
rect 4624 2259 4680 2279
rect 5350 2259 5406 2279
rect 5460 2259 5516 2279
rect 9011 2414 9067 2470
rect 9121 2414 9177 2470
rect 5630 2279 5686 2321
rect 5740 2279 5796 2321
rect 6749 2279 6805 2314
rect 6859 2279 6915 2314
rect 5630 2265 5686 2279
rect 5740 2265 5796 2279
rect 6749 2258 6805 2279
rect 6859 2258 6915 2279
rect 7028 2279 7084 2316
rect 7138 2279 7194 2316
rect 7028 2260 7084 2279
rect 7138 2260 7194 2279
rect 7316 2279 7372 2316
rect 7426 2279 7482 2316
rect 7316 2260 7372 2279
rect 7426 2260 7482 2279
rect 7595 2279 7651 2314
rect 7705 2279 7761 2314
rect 8714 2279 8770 2321
rect 8824 2279 8880 2321
rect 7595 2258 7651 2279
rect 7705 2258 7761 2279
rect 8714 2265 8770 2279
rect 8824 2265 8880 2279
rect 8994 2279 9050 2315
rect 9104 2279 9160 2315
rect 8994 2259 9050 2279
rect 9104 2259 9160 2279
rect -341 1962 -285 2018
rect -464 1840 -408 1896
rect -341 1852 -285 1908
rect 868 1993 924 2009
rect 978 1993 1034 2009
rect 868 1953 924 1993
rect 978 1953 1034 1993
rect -464 1730 -408 1786
rect 100 1841 156 1897
rect 210 1841 266 1897
rect 1148 1993 1204 2010
rect 1258 1993 1314 2010
rect 2270 1993 2326 2008
rect 2380 1993 2436 2008
rect 1148 1954 1204 1993
rect 1258 1954 1314 1993
rect 2270 1952 2326 1993
rect 2380 1952 2436 1993
rect 2553 1993 2609 2008
rect 2663 1993 2719 2008
rect 2833 1993 2889 2008
rect 2943 1993 2999 2008
rect 2553 1952 2609 1993
rect 2663 1952 2719 1993
rect 2833 1952 2889 1993
rect 2943 1952 2999 1993
rect 3114 1993 3170 2008
rect 3224 1993 3280 2008
rect 4236 1993 4292 2010
rect 4346 1993 4402 2010
rect 3114 1952 3170 1993
rect 3224 1952 3280 1993
rect 4236 1954 4292 1993
rect 4346 1954 4402 1993
rect 4516 1993 4572 2009
rect 4626 1993 4682 2009
rect 4516 1953 4572 1993
rect 4626 1953 4682 1993
rect 5348 1993 5404 2009
rect 5458 1993 5514 2009
rect 5348 1953 5404 1993
rect 5458 1953 5514 1993
rect 5628 1993 5684 2010
rect 5738 1993 5794 2010
rect 6750 1993 6806 2008
rect 6860 1993 6916 2008
rect 7594 1993 7650 2008
rect 7704 1993 7760 2008
rect 8716 1993 8772 2010
rect 8826 1993 8882 2010
rect 5628 1954 5684 1993
rect 5738 1954 5794 1993
rect 6750 1952 6806 1993
rect 6860 1952 6916 1993
rect 7594 1952 7650 1993
rect 7704 1952 7760 1993
rect 8716 1954 8772 1993
rect 8826 1954 8882 1993
rect 366 1724 422 1780
rect 476 1724 532 1780
rect 1261 1725 1317 1781
rect 868 1627 924 1667
rect 978 1627 1034 1667
rect 1429 1627 1485 1666
rect 1539 1627 1595 1666
rect 868 1611 924 1627
rect 978 1611 1034 1627
rect 1429 1610 1485 1627
rect 1539 1610 1595 1627
rect 4233 1725 4289 1781
rect 1710 1627 1766 1667
rect 1820 1627 1876 1667
rect 3674 1627 3730 1667
rect 3784 1627 3840 1667
rect 1710 1611 1766 1627
rect 1820 1611 1876 1627
rect 3674 1611 3730 1627
rect 3784 1611 3840 1627
rect 8996 1993 9052 2009
rect 9106 1993 9162 2009
rect 8996 1953 9052 1993
rect 9106 1953 9162 1993
rect 9503 2146 9559 2202
rect 9613 2146 9669 2202
rect 10126 2267 10182 2323
rect 10126 2157 10182 2213
rect 10236 4050 10292 4106
rect 10236 3940 10292 3996
rect 5741 1725 5797 1781
rect 3955 1627 4011 1666
rect 4065 1627 4121 1666
rect 4516 1627 4572 1667
rect 4626 1627 4682 1667
rect 3955 1610 4011 1627
rect 4065 1610 4121 1627
rect 4516 1611 4572 1627
rect 4626 1611 4682 1627
rect 5348 1627 5404 1667
rect 5458 1627 5514 1667
rect 5909 1627 5965 1666
rect 6019 1627 6075 1666
rect 5348 1611 5404 1627
rect 5458 1611 5514 1627
rect 5909 1610 5965 1627
rect 6019 1610 6075 1627
rect 8713 1725 8769 1781
rect 6190 1627 6246 1667
rect 6300 1627 6356 1667
rect 8154 1627 8210 1667
rect 8264 1627 8320 1667
rect 6190 1611 6246 1627
rect 6300 1611 6356 1627
rect 8154 1611 8210 1627
rect 8264 1611 8320 1627
rect 9502 1724 9558 1780
rect 9612 1724 9668 1780
rect 8435 1627 8491 1666
rect 8545 1627 8601 1666
rect 8996 1627 9052 1667
rect 9106 1627 9162 1667
rect 8435 1610 8491 1627
rect 8545 1610 8601 1627
rect 8996 1611 9052 1627
rect 9106 1611 9162 1627
rect 101 1500 157 1556
rect 211 1500 267 1556
rect 870 1341 926 1364
rect 980 1341 1036 1364
rect -575 1248 -519 1304
rect -575 1138 -519 1194
rect 870 1308 926 1341
rect 980 1308 1036 1341
rect 1428 1341 1484 1367
rect 1538 1341 1594 1367
rect 1428 1311 1484 1341
rect 1538 1311 1594 1341
rect 2267 1341 2323 1353
rect 2377 1341 2433 1353
rect 3117 1341 3173 1353
rect 3227 1341 3283 1353
rect 2267 1297 2268 1341
rect 2268 1297 2323 1341
rect 2377 1297 2433 1341
rect 3117 1297 3173 1341
rect 3227 1297 3282 1341
rect 3282 1297 3283 1341
rect 6747 1341 6803 1353
rect 6857 1341 6913 1353
rect 7597 1341 7653 1353
rect 7707 1341 7763 1353
rect 6747 1297 6748 1341
rect 6748 1297 6803 1341
rect 6857 1297 6913 1341
rect 7597 1297 7653 1341
rect 7707 1297 7762 1341
rect 7762 1297 7763 1341
rect 9751 1500 9807 1556
rect 9861 1500 9917 1556
rect 9501 1397 9557 1453
rect 9611 1397 9667 1453
rect 10236 1622 10292 1678
rect 10236 1512 10292 1568
rect 10365 3848 10421 3904
rect 10365 3738 10421 3794
rect 105 1127 161 1183
rect 215 1127 271 1183
rect 10484 3677 10540 3733
rect 10365 1420 10421 1476
rect 10365 1310 10421 1366
rect 10484 3567 10540 3623
rect 9731 1127 9787 1183
rect 9841 1127 9897 1183
rect 10484 1249 10540 1305
rect 10484 1139 10540 1195
<< metal2 >>
rect 2454 5512 2644 5516
rect 2454 5456 2466 5512
rect 2522 5456 2576 5512
rect 2632 5456 2644 5512
rect 2454 5452 2644 5456
rect 2906 5512 3096 5516
rect 2906 5456 2918 5512
rect 2974 5456 3028 5512
rect 3084 5456 3096 5512
rect 2906 5452 3096 5456
rect 6934 5512 7124 5516
rect 6934 5456 6946 5512
rect 7002 5456 7056 5512
rect 7112 5456 7124 5512
rect 6934 5452 7124 5456
rect 7386 5512 7576 5516
rect 7386 5456 7398 5512
rect 7454 5456 7508 5512
rect 7564 5456 7576 5512
rect 7386 5452 7576 5456
rect 1709 5410 1765 5411
rect 1695 5401 1895 5410
rect 1695 5345 1709 5401
rect 1765 5345 1819 5401
rect 1875 5345 1895 5401
rect 1695 5333 1895 5345
rect 1428 5101 1484 5103
rect 855 5091 1055 5100
rect 603 5086 1055 5091
rect 603 5030 867 5086
rect 923 5030 975 5086
rect 1031 5030 1055 5086
rect 603 5025 1055 5030
rect 333 4967 530 4972
rect 333 4911 349 4967
rect 405 4911 459 4967
rect 515 4911 530 4967
rect 333 4906 530 4911
rect -236 4752 -170 4767
rect -236 4696 -231 4752
rect -175 4696 -170 4752
rect -236 4642 -170 4696
rect -236 4586 -231 4642
rect -175 4636 -170 4642
rect -175 4631 293 4636
rect -175 4586 109 4631
rect -236 4575 109 4586
rect 165 4575 219 4631
rect 275 4575 293 4631
rect -236 4570 293 4575
rect -346 4447 -280 4462
rect -346 4391 -341 4447
rect -285 4391 -280 4447
rect -468 4325 -402 4340
rect -468 4269 -463 4325
rect -407 4269 -402 4325
rect -468 4215 -402 4269
rect -346 4337 -280 4391
rect -346 4281 -341 4337
rect -285 4331 -280 4337
rect -285 4326 284 4331
rect -285 4281 100 4326
rect -346 4270 100 4281
rect 156 4270 210 4326
rect 266 4270 284 4326
rect -346 4265 284 4270
rect -468 4159 -463 4215
rect -407 4209 -402 4215
rect 430 4214 496 4906
rect 350 4209 547 4214
rect -407 4159 366 4209
rect -468 4153 366 4159
rect 422 4153 476 4209
rect 532 4153 547 4209
rect -468 4148 547 4153
rect -468 4143 350 4148
rect 88 3985 285 3990
rect 88 3929 101 3985
rect 157 3929 211 3985
rect 267 3929 285 3985
rect 88 3924 285 3929
rect -582 3733 -516 3748
rect -582 3677 -577 3733
rect -521 3677 -516 3733
rect -582 3623 -516 3677
rect -582 3567 -577 3623
rect -521 3617 -516 3623
rect 603 3676 669 5025
rect 855 5023 1055 5025
rect 1415 5093 1615 5101
rect 1415 5037 1428 5093
rect 1484 5037 1538 5093
rect 1594 5037 1615 5093
rect 1415 5024 1615 5037
rect 1695 5090 1895 5101
rect 1695 5034 1709 5090
rect 1765 5034 1819 5090
rect 1875 5034 1895 5090
rect 1695 5024 1895 5034
rect 2255 5087 2455 5101
rect 2255 5031 2267 5087
rect 2323 5031 2377 5087
rect 2433 5031 2455 5087
rect 2255 5024 2455 5031
rect 865 5020 921 5023
rect 1250 4965 1442 4968
rect 1250 4909 1262 4965
rect 1318 4909 1372 4965
rect 1428 4909 1442 4965
rect 1250 4906 1442 4909
rect 839 4900 1029 4904
rect 839 4844 851 4900
rect 907 4844 961 4900
rect 1017 4844 1029 4900
rect 839 4839 1029 4844
rect 851 4838 1029 4839
rect 1256 4758 1322 4906
rect 855 4744 1055 4756
rect 855 4688 870 4744
rect 926 4688 980 4744
rect 1036 4688 1055 4744
rect 855 4678 1055 4688
rect 1135 4750 1335 4758
rect 1135 4694 1150 4750
rect 1206 4694 1260 4750
rect 1316 4694 1335 4750
rect 1135 4681 1335 4694
rect 1812 4700 1884 5024
rect 2542 4758 2608 5452
rect 2942 4758 3008 5452
rect 3785 5410 3841 5411
rect 6189 5410 6245 5411
rect 3655 5401 3855 5410
rect 3655 5345 3675 5401
rect 3731 5345 3785 5401
rect 3841 5345 3855 5401
rect 3655 5333 3855 5345
rect 6175 5401 6375 5410
rect 6175 5345 6189 5401
rect 6245 5345 6299 5401
rect 6355 5345 6375 5401
rect 6175 5333 6375 5345
rect 4066 5101 4122 5103
rect 5908 5101 5964 5103
rect 3095 5087 3295 5101
rect 3095 5031 3117 5087
rect 3173 5031 3227 5087
rect 3283 5031 3295 5087
rect 3095 5024 3295 5031
rect 3655 5090 3855 5101
rect 3655 5034 3675 5090
rect 3731 5034 3785 5090
rect 3841 5034 3855 5090
rect 3655 5024 3855 5034
rect 3935 5093 4135 5101
rect 3935 5037 3956 5093
rect 4012 5037 4066 5093
rect 4122 5037 4135 5093
rect 3935 5024 4135 5037
rect 4495 5091 4695 5100
rect 5335 5091 5535 5100
rect 4495 5086 4947 5091
rect 4495 5030 4519 5086
rect 4575 5030 4627 5086
rect 4683 5030 4947 5086
rect 4495 5025 4947 5030
rect 2255 4743 2455 4757
rect 2255 4700 2269 4743
rect 1812 4687 2269 4700
rect 2325 4687 2379 4743
rect 2435 4687 2455 4743
rect 1812 4677 2455 4687
rect 2535 4745 2735 4758
rect 2535 4689 2548 4745
rect 2604 4689 2658 4745
rect 2714 4689 2735 4745
rect 2535 4681 2735 4689
rect 2815 4745 3015 4758
rect 2815 4689 2836 4745
rect 2892 4689 2946 4745
rect 3002 4689 3015 4745
rect 2815 4681 3015 4689
rect 3095 4743 3295 4757
rect 3095 4687 3115 4743
rect 3171 4687 3225 4743
rect 3281 4700 3295 4743
rect 3666 4700 3738 5024
rect 4495 5023 4695 5025
rect 4629 5020 4685 5023
rect 4108 4965 4300 4968
rect 4108 4909 4122 4965
rect 4178 4909 4232 4965
rect 4288 4909 4300 4965
rect 4108 4906 4300 4909
rect 4228 4758 4294 4906
rect 4519 4899 4709 4904
rect 4519 4843 4531 4899
rect 4587 4843 4641 4899
rect 4697 4843 4709 4899
rect 4519 4838 4709 4843
rect 3281 4687 3738 4700
rect 2548 4679 2675 4681
rect 1812 4628 2370 4677
rect 855 4438 1055 4448
rect 855 4382 868 4438
rect 924 4382 978 4438
rect 1034 4382 1055 4438
rect 855 4371 1055 4382
rect 1135 4439 1335 4449
rect 1135 4383 1148 4439
rect 1204 4383 1258 4439
rect 1314 4383 1335 4439
rect 1135 4372 1335 4383
rect 2255 4437 2455 4449
rect 2599 4442 2675 4679
rect 2890 4679 3002 4681
rect 2890 4442 2966 4679
rect 3095 4677 3738 4687
rect 4215 4750 4415 4758
rect 4215 4694 4234 4750
rect 4290 4694 4344 4750
rect 4400 4694 4415 4750
rect 4215 4681 4415 4694
rect 4495 4744 4695 4756
rect 4495 4688 4514 4744
rect 4570 4688 4624 4744
rect 4680 4688 4695 4744
rect 4495 4678 4695 4688
rect 3180 4628 3738 4677
rect 2255 4381 2270 4437
rect 2326 4381 2380 4437
rect 2436 4381 2455 4437
rect 1256 4215 1322 4372
rect 2255 4371 2455 4381
rect 2537 4437 2734 4442
rect 2537 4381 2553 4437
rect 2609 4381 2663 4437
rect 2719 4381 2734 4437
rect 2537 4376 2734 4381
rect 2817 4437 3014 4442
rect 2817 4381 2833 4437
rect 2889 4381 2943 4437
rect 2999 4381 3014 4437
rect 2817 4376 3014 4381
rect 3095 4437 3295 4449
rect 3095 4381 3114 4437
rect 3170 4381 3224 4437
rect 3280 4381 3295 4437
rect 3095 4371 3295 4381
rect 4215 4439 4415 4449
rect 4215 4383 4236 4439
rect 4292 4383 4346 4439
rect 4402 4383 4415 4439
rect 4215 4372 4415 4383
rect 4495 4438 4695 4448
rect 4495 4382 4516 4438
rect 4572 4382 4626 4438
rect 4682 4382 4695 4438
rect 2272 4249 2340 4371
rect 1249 4210 1329 4215
rect 1249 4154 1261 4210
rect 1317 4154 1329 4210
rect 1249 4148 1329 4154
rect 1777 4181 2340 4249
rect 3210 4249 3278 4371
rect 3210 4181 3773 4249
rect 4228 4215 4294 4372
rect 4495 4371 4695 4382
rect 1777 4106 1845 4181
rect 3705 4106 3773 4181
rect 4221 4210 4301 4215
rect 4221 4154 4233 4210
rect 4289 4154 4301 4210
rect 4221 4148 4301 4154
rect 855 4096 1055 4106
rect 855 4040 868 4096
rect 924 4040 978 4096
rect 1034 4040 1055 4096
rect 855 4029 1055 4040
rect 1415 4095 1615 4106
rect 1415 4039 1429 4095
rect 1485 4039 1539 4095
rect 1595 4039 1615 4095
rect 1415 4029 1615 4039
rect 1695 4096 1895 4106
rect 1695 4040 1710 4096
rect 1766 4040 1820 4096
rect 1876 4040 1895 4096
rect 1695 4029 1895 4040
rect 3655 4096 3855 4106
rect 3655 4040 3674 4096
rect 3730 4040 3784 4096
rect 3840 4040 3855 4096
rect 3655 4029 3855 4040
rect 3935 4095 4135 4106
rect 3935 4039 3955 4095
rect 4011 4039 4065 4095
rect 4121 4039 4135 4095
rect 3935 4029 4135 4039
rect 4495 4096 4695 4106
rect 4495 4040 4516 4096
rect 4572 4040 4626 4096
rect 4682 4040 4695 4096
rect 4495 4029 4695 4040
rect 1477 3800 1547 4029
rect 857 3793 1054 3798
rect 857 3737 870 3793
rect 926 3737 980 3793
rect 1036 3737 1054 3793
rect 857 3732 1054 3737
rect 1415 3795 1612 3800
rect 1415 3739 1428 3795
rect 1484 3739 1538 3795
rect 1594 3739 1612 3795
rect 1415 3734 1612 3739
rect 2255 3782 2455 3797
rect 2255 3726 2267 3782
rect 2323 3726 2377 3782
rect 2433 3726 2455 3782
rect 2255 3720 2455 3726
rect 3095 3782 3295 3797
rect 3095 3726 3117 3782
rect 3173 3726 3227 3782
rect 3283 3726 3295 3782
rect 3095 3720 3295 3726
rect 2255 3716 2323 3720
rect 3227 3716 3295 3720
rect 2255 3676 2321 3716
rect -521 3612 289 3617
rect -521 3567 105 3612
rect -582 3556 105 3567
rect 161 3556 215 3612
rect 271 3556 289 3612
rect 603 3610 2321 3676
rect 3229 3676 3295 3716
rect 4881 3676 4947 5025
rect 3229 3610 4947 3676
rect 5083 5086 5535 5091
rect 5083 5030 5347 5086
rect 5403 5030 5455 5086
rect 5511 5030 5535 5086
rect 5083 5025 5535 5030
rect 5083 3676 5149 5025
rect 5335 5023 5535 5025
rect 5895 5093 6095 5101
rect 5895 5037 5908 5093
rect 5964 5037 6018 5093
rect 6074 5037 6095 5093
rect 5895 5024 6095 5037
rect 6175 5090 6375 5101
rect 6175 5034 6189 5090
rect 6245 5034 6299 5090
rect 6355 5034 6375 5090
rect 6175 5024 6375 5034
rect 6735 5087 6935 5101
rect 6735 5031 6747 5087
rect 6803 5031 6857 5087
rect 6913 5031 6935 5087
rect 6735 5024 6935 5031
rect 5345 5020 5401 5023
rect 5730 4965 5922 4968
rect 5730 4909 5742 4965
rect 5798 4909 5852 4965
rect 5908 4909 5922 4965
rect 5730 4906 5922 4909
rect 5319 4900 5509 4904
rect 5319 4844 5331 4900
rect 5387 4844 5441 4900
rect 5497 4844 5509 4900
rect 5319 4839 5509 4844
rect 5331 4838 5509 4839
rect 5736 4758 5802 4906
rect 5335 4744 5535 4756
rect 5335 4688 5350 4744
rect 5406 4688 5460 4744
rect 5516 4688 5535 4744
rect 5335 4678 5535 4688
rect 5615 4750 5815 4758
rect 5615 4694 5630 4750
rect 5686 4694 5740 4750
rect 5796 4694 5815 4750
rect 5615 4681 5815 4694
rect 6292 4700 6364 5024
rect 7022 4758 7088 5452
rect 7422 4758 7488 5452
rect 8265 5410 8321 5411
rect 8135 5401 8335 5410
rect 8135 5345 8155 5401
rect 8211 5345 8265 5401
rect 8321 5345 8335 5401
rect 8135 5333 8335 5345
rect 8546 5101 8602 5103
rect 7575 5087 7775 5101
rect 7575 5031 7597 5087
rect 7653 5031 7707 5087
rect 7763 5031 7775 5087
rect 7575 5024 7775 5031
rect 8135 5090 8335 5101
rect 8135 5034 8155 5090
rect 8211 5034 8265 5090
rect 8321 5034 8335 5090
rect 8135 5024 8335 5034
rect 8415 5093 8615 5101
rect 8415 5037 8436 5093
rect 8492 5037 8546 5093
rect 8602 5037 8615 5093
rect 8415 5024 8615 5037
rect 8975 5091 9175 5100
rect 8975 5086 9427 5091
rect 8975 5030 8999 5086
rect 9055 5030 9107 5086
rect 9163 5030 9427 5086
rect 8975 5025 9427 5030
rect 6735 4743 6935 4757
rect 6735 4700 6749 4743
rect 6292 4687 6749 4700
rect 6805 4687 6859 4743
rect 6915 4687 6935 4743
rect 6292 4677 6935 4687
rect 7015 4745 7215 4758
rect 7015 4689 7028 4745
rect 7084 4689 7138 4745
rect 7194 4689 7215 4745
rect 7015 4681 7215 4689
rect 7295 4745 7495 4758
rect 7295 4689 7316 4745
rect 7372 4689 7426 4745
rect 7482 4689 7495 4745
rect 7295 4681 7495 4689
rect 7575 4743 7775 4757
rect 7575 4687 7595 4743
rect 7651 4687 7705 4743
rect 7761 4700 7775 4743
rect 8146 4700 8218 5024
rect 8975 5023 9175 5025
rect 9109 5020 9165 5023
rect 8588 4965 8780 4968
rect 8588 4909 8602 4965
rect 8658 4909 8712 4965
rect 8768 4909 8780 4965
rect 8588 4906 8780 4909
rect 8708 4758 8774 4906
rect 8999 4899 9189 4904
rect 8999 4843 9011 4899
rect 9067 4843 9121 4899
rect 9177 4843 9189 4899
rect 8999 4838 9189 4843
rect 7761 4687 8218 4700
rect 7028 4679 7084 4681
rect 7426 4679 7482 4681
rect 7575 4677 8218 4687
rect 8695 4750 8895 4758
rect 8695 4694 8714 4750
rect 8770 4694 8824 4750
rect 8880 4694 8895 4750
rect 8695 4681 8895 4694
rect 8975 4744 9175 4756
rect 8975 4688 8994 4744
rect 9050 4688 9104 4744
rect 9160 4688 9175 4744
rect 8975 4678 9175 4688
rect 6292 4628 6850 4677
rect 7660 4628 8218 4677
rect 5335 4438 5535 4448
rect 5335 4382 5348 4438
rect 5404 4382 5458 4438
rect 5514 4382 5535 4438
rect 5335 4371 5535 4382
rect 5615 4439 5815 4449
rect 5615 4383 5628 4439
rect 5684 4383 5738 4439
rect 5794 4383 5815 4439
rect 5615 4372 5815 4383
rect 6735 4437 6935 4449
rect 6735 4381 6750 4437
rect 6806 4381 6860 4437
rect 6916 4381 6935 4437
rect 5736 4215 5802 4372
rect 6735 4371 6935 4381
rect 7575 4437 7775 4449
rect 7575 4381 7594 4437
rect 7650 4381 7704 4437
rect 7760 4381 7775 4437
rect 7575 4371 7775 4381
rect 8695 4439 8895 4449
rect 8695 4383 8716 4439
rect 8772 4383 8826 4439
rect 8882 4383 8895 4439
rect 8695 4372 8895 4383
rect 8975 4438 9175 4448
rect 8975 4382 8996 4438
rect 9052 4382 9106 4438
rect 9162 4382 9175 4438
rect 6752 4249 6820 4371
rect 5729 4210 5809 4215
rect 5729 4154 5741 4210
rect 5797 4154 5809 4210
rect 5729 4148 5809 4154
rect 6257 4181 6820 4249
rect 7690 4249 7758 4371
rect 7690 4181 8253 4249
rect 8708 4215 8774 4372
rect 8975 4371 9175 4382
rect 6257 4106 6325 4181
rect 8185 4106 8253 4181
rect 8701 4210 8781 4215
rect 8701 4154 8713 4210
rect 8769 4154 8781 4210
rect 8701 4148 8781 4154
rect 5335 4096 5535 4106
rect 5335 4040 5348 4096
rect 5404 4040 5458 4096
rect 5514 4040 5535 4096
rect 5335 4029 5535 4040
rect 5895 4095 6095 4106
rect 5895 4039 5909 4095
rect 5965 4039 6019 4095
rect 6075 4039 6095 4095
rect 5895 4029 6095 4039
rect 6175 4096 6375 4106
rect 6175 4040 6190 4096
rect 6246 4040 6300 4096
rect 6356 4040 6375 4096
rect 6175 4029 6375 4040
rect 8135 4096 8335 4106
rect 8135 4040 8154 4096
rect 8210 4040 8264 4096
rect 8320 4040 8335 4096
rect 8135 4029 8335 4040
rect 8415 4095 8615 4106
rect 8415 4039 8435 4095
rect 8491 4039 8545 4095
rect 8601 4039 8615 4095
rect 8415 4029 8615 4039
rect 8975 4096 9175 4106
rect 8975 4040 8996 4096
rect 9052 4040 9106 4096
rect 9162 4040 9175 4096
rect 8975 4029 9175 4040
rect 6735 3782 6935 3797
rect 6735 3726 6747 3782
rect 6803 3726 6857 3782
rect 6913 3726 6935 3782
rect 6735 3720 6935 3726
rect 7575 3782 7775 3797
rect 7575 3726 7597 3782
rect 7653 3726 7707 3782
rect 7763 3726 7775 3782
rect 7575 3720 7775 3726
rect 6735 3716 6803 3720
rect 7707 3716 7775 3720
rect 6735 3676 6801 3716
rect 5083 3610 6801 3676
rect 7709 3676 7775 3716
rect 9361 3676 9427 5025
rect 9700 4967 9897 4972
rect 9700 4911 9713 4967
rect 9771 4911 9823 4967
rect 9881 4911 9897 4967
rect 9700 4906 9897 4911
rect 10122 4645 10185 4660
rect 10122 4636 10127 4645
rect 9485 4631 10127 4636
rect 9485 4575 9503 4631
rect 9559 4575 9613 4631
rect 9669 4589 10127 4631
rect 10183 4636 10185 4645
rect 10183 4589 10311 4636
rect 9669 4575 10311 4589
rect 9485 4570 10311 4575
rect 10122 4535 10185 4570
rect 10122 4479 10127 4535
rect 10183 4479 10185 4535
rect 10122 4462 10185 4479
rect 9484 4209 9681 4214
rect 9484 4153 9502 4209
rect 9558 4153 9612 4209
rect 9668 4153 9681 4209
rect 9484 4148 9681 4153
rect 9555 3887 9621 4148
rect 10231 4106 10297 4121
rect 10231 4050 10236 4106
rect 10292 4050 10297 4106
rect 10231 3996 10297 4050
rect 10231 3990 10236 3996
rect 9733 3985 10236 3990
rect 9733 3929 9751 3985
rect 9807 3929 9861 3985
rect 9917 3940 10236 3985
rect 10292 3940 10297 3996
rect 9917 3929 10297 3940
rect 9733 3924 10297 3929
rect 10360 3904 10423 3919
rect 9483 3882 9680 3887
rect 9483 3826 9501 3882
rect 9557 3826 9611 3882
rect 9667 3826 9680 3882
rect 9483 3821 9680 3826
rect 9614 3788 9680 3821
rect 10360 3848 10365 3904
rect 10421 3848 10423 3904
rect 10360 3794 10423 3848
rect 10360 3788 10365 3794
rect 9614 3738 10365 3788
rect 10421 3738 10423 3794
rect 9614 3722 10423 3738
rect 10481 3733 10545 3748
rect 7709 3610 9427 3676
rect 10481 3677 10484 3733
rect 10540 3677 10545 3733
rect 10481 3623 10545 3677
rect 10481 3617 10484 3623
rect 9713 3612 10484 3617
rect -582 3551 289 3556
rect 9713 3556 9731 3612
rect 9787 3556 9841 3612
rect 9897 3567 10484 3612
rect 10540 3567 10545 3623
rect 9897 3556 10545 3567
rect 9713 3551 10545 3556
rect 2454 3083 2644 3087
rect 2454 3027 2466 3083
rect 2522 3027 2576 3083
rect 2632 3027 2644 3083
rect 2454 3023 2644 3027
rect 2906 3083 3096 3087
rect 2906 3027 2918 3083
rect 2974 3027 3028 3083
rect 3084 3027 3096 3083
rect 2906 3023 3096 3027
rect 6934 3083 7124 3087
rect 6934 3027 6946 3083
rect 7002 3027 7056 3083
rect 7112 3027 7124 3083
rect 6934 3023 7124 3027
rect 7386 3083 7576 3087
rect 7386 3027 7398 3083
rect 7454 3027 7508 3083
rect 7564 3027 7576 3083
rect 7386 3023 7576 3027
rect 1709 2981 1765 2982
rect 1695 2972 1895 2981
rect 1695 2916 1709 2972
rect 1765 2916 1819 2972
rect 1875 2916 1895 2972
rect 1695 2904 1895 2916
rect 1428 2672 1484 2674
rect 855 2662 1055 2671
rect 603 2657 1055 2662
rect 603 2601 867 2657
rect 923 2601 975 2657
rect 1031 2601 1055 2657
rect 603 2596 1055 2601
rect 333 2538 530 2543
rect 333 2482 349 2538
rect 405 2482 459 2538
rect 515 2482 530 2538
rect 333 2477 530 2482
rect -234 2323 -168 2338
rect -234 2267 -229 2323
rect -173 2267 -168 2323
rect -234 2213 -168 2267
rect -234 2207 -229 2213
rect -236 2157 -229 2207
rect -173 2207 -168 2213
rect -173 2202 293 2207
rect -173 2157 109 2202
rect -236 2146 109 2157
rect 165 2146 219 2202
rect 275 2146 293 2202
rect -236 2141 293 2146
rect -346 2018 -280 2033
rect -346 1962 -341 2018
rect -285 1962 -280 2018
rect -469 1896 -403 1911
rect -469 1840 -464 1896
rect -408 1840 -403 1896
rect -469 1786 -403 1840
rect -346 1908 -280 1962
rect -346 1852 -341 1908
rect -285 1902 -280 1908
rect -285 1897 284 1902
rect -285 1852 100 1897
rect -346 1841 100 1852
rect 156 1841 210 1897
rect 266 1841 284 1897
rect -346 1836 284 1841
rect -469 1730 -464 1786
rect -408 1780 -403 1786
rect 430 1785 496 2477
rect 350 1780 547 1785
rect -408 1730 366 1780
rect -469 1724 366 1730
rect 422 1724 476 1780
rect 532 1724 547 1780
rect -469 1719 547 1724
rect -469 1714 350 1719
rect 88 1556 285 1561
rect 88 1500 101 1556
rect 157 1500 211 1556
rect 267 1500 285 1556
rect 88 1495 285 1500
rect -580 1304 -514 1319
rect -580 1248 -575 1304
rect -519 1248 -514 1304
rect -580 1194 -514 1248
rect -580 1138 -575 1194
rect -519 1188 -514 1194
rect 603 1247 669 2596
rect 855 2594 1055 2596
rect 1415 2664 1615 2672
rect 1415 2608 1428 2664
rect 1484 2608 1538 2664
rect 1594 2608 1615 2664
rect 1415 2595 1615 2608
rect 1695 2661 1895 2672
rect 1695 2605 1709 2661
rect 1765 2605 1819 2661
rect 1875 2605 1895 2661
rect 1695 2595 1895 2605
rect 2255 2658 2455 2672
rect 2255 2602 2267 2658
rect 2323 2602 2377 2658
rect 2433 2602 2455 2658
rect 2255 2595 2455 2602
rect 865 2591 921 2594
rect 1250 2536 1442 2539
rect 1250 2480 1262 2536
rect 1318 2480 1372 2536
rect 1428 2480 1442 2536
rect 1250 2477 1442 2480
rect 839 2471 1029 2475
rect 839 2415 851 2471
rect 907 2415 961 2471
rect 1017 2415 1029 2471
rect 839 2410 1029 2415
rect 851 2409 1029 2410
rect 1256 2329 1322 2477
rect 855 2315 1055 2327
rect 855 2259 870 2315
rect 926 2259 980 2315
rect 1036 2259 1055 2315
rect 855 2249 1055 2259
rect 1135 2321 1335 2329
rect 1135 2265 1150 2321
rect 1206 2265 1260 2321
rect 1316 2265 1335 2321
rect 1135 2252 1335 2265
rect 1812 2271 1884 2595
rect 2542 2329 2608 3023
rect 2942 2329 3008 3023
rect 3785 2981 3841 2982
rect 6189 2981 6245 2982
rect 3655 2972 3855 2981
rect 3655 2916 3675 2972
rect 3731 2916 3785 2972
rect 3841 2916 3855 2972
rect 3655 2904 3855 2916
rect 6175 2972 6375 2981
rect 6175 2916 6189 2972
rect 6245 2916 6299 2972
rect 6355 2916 6375 2972
rect 6175 2904 6375 2916
rect 4066 2672 4122 2674
rect 5908 2672 5964 2674
rect 3095 2658 3295 2672
rect 3095 2602 3117 2658
rect 3173 2602 3227 2658
rect 3283 2602 3295 2658
rect 3095 2595 3295 2602
rect 3655 2661 3855 2672
rect 3655 2605 3675 2661
rect 3731 2605 3785 2661
rect 3841 2605 3855 2661
rect 3655 2595 3855 2605
rect 3935 2664 4135 2672
rect 3935 2608 3956 2664
rect 4012 2608 4066 2664
rect 4122 2608 4135 2664
rect 3935 2595 4135 2608
rect 4495 2662 4695 2671
rect 5335 2662 5535 2671
rect 4495 2657 4947 2662
rect 4495 2601 4519 2657
rect 4575 2601 4627 2657
rect 4683 2601 4947 2657
rect 4495 2596 4947 2601
rect 2255 2314 2455 2328
rect 2255 2271 2269 2314
rect 1812 2258 2269 2271
rect 2325 2258 2379 2314
rect 2435 2258 2455 2314
rect 1812 2248 2455 2258
rect 2535 2316 2735 2329
rect 2535 2260 2548 2316
rect 2604 2260 2658 2316
rect 2714 2260 2735 2316
rect 2535 2252 2735 2260
rect 2815 2316 3015 2329
rect 2815 2260 2836 2316
rect 2892 2260 2946 2316
rect 3002 2260 3015 2316
rect 2815 2252 3015 2260
rect 3095 2314 3295 2328
rect 3095 2258 3115 2314
rect 3171 2258 3225 2314
rect 3281 2271 3295 2314
rect 3666 2271 3738 2595
rect 4495 2594 4695 2596
rect 4629 2591 4685 2594
rect 4108 2536 4300 2539
rect 4108 2480 4122 2536
rect 4178 2480 4232 2536
rect 4288 2480 4300 2536
rect 4108 2477 4300 2480
rect 4228 2329 4294 2477
rect 4519 2470 4709 2475
rect 4519 2414 4531 2470
rect 4587 2414 4641 2470
rect 4697 2414 4709 2470
rect 4519 2409 4709 2414
rect 3281 2258 3738 2271
rect 2548 2250 2675 2252
rect 1812 2199 2370 2248
rect 855 2009 1055 2019
rect 855 1953 868 2009
rect 924 1953 978 2009
rect 1034 1953 1055 2009
rect 855 1942 1055 1953
rect 1135 2010 1335 2020
rect 1135 1954 1148 2010
rect 1204 1954 1258 2010
rect 1314 1954 1335 2010
rect 1135 1943 1335 1954
rect 2255 2008 2455 2020
rect 2599 2013 2675 2250
rect 2890 2250 3002 2252
rect 2890 2013 2966 2250
rect 3095 2248 3738 2258
rect 4215 2321 4415 2329
rect 4215 2265 4234 2321
rect 4290 2265 4344 2321
rect 4400 2265 4415 2321
rect 4215 2252 4415 2265
rect 4495 2315 4695 2327
rect 4495 2259 4514 2315
rect 4570 2259 4624 2315
rect 4680 2259 4695 2315
rect 4495 2249 4695 2259
rect 3180 2199 3738 2248
rect 2255 1952 2270 2008
rect 2326 1952 2380 2008
rect 2436 1952 2455 2008
rect 1256 1786 1322 1943
rect 2255 1942 2455 1952
rect 2537 2008 2734 2013
rect 2537 1952 2553 2008
rect 2609 1952 2663 2008
rect 2719 1952 2734 2008
rect 2537 1947 2734 1952
rect 2817 2008 3014 2013
rect 2817 1952 2833 2008
rect 2889 1952 2943 2008
rect 2999 1952 3014 2008
rect 2817 1947 3014 1952
rect 3095 2008 3295 2020
rect 3095 1952 3114 2008
rect 3170 1952 3224 2008
rect 3280 1952 3295 2008
rect 3095 1942 3295 1952
rect 4215 2010 4415 2020
rect 4215 1954 4236 2010
rect 4292 1954 4346 2010
rect 4402 1954 4415 2010
rect 4215 1943 4415 1954
rect 4495 2009 4695 2019
rect 4495 1953 4516 2009
rect 4572 1953 4626 2009
rect 4682 1953 4695 2009
rect 2272 1820 2340 1942
rect 1249 1781 1329 1786
rect 1249 1725 1261 1781
rect 1317 1725 1329 1781
rect 1249 1719 1329 1725
rect 1777 1752 2340 1820
rect 3210 1820 3278 1942
rect 3210 1752 3773 1820
rect 4228 1786 4294 1943
rect 4495 1942 4695 1953
rect 1777 1677 1845 1752
rect 3705 1677 3773 1752
rect 4221 1781 4301 1786
rect 4221 1725 4233 1781
rect 4289 1725 4301 1781
rect 4221 1719 4301 1725
rect 855 1667 1055 1677
rect 855 1611 868 1667
rect 924 1611 978 1667
rect 1034 1611 1055 1667
rect 855 1600 1055 1611
rect 1415 1666 1615 1677
rect 1415 1610 1429 1666
rect 1485 1610 1539 1666
rect 1595 1610 1615 1666
rect 1415 1600 1615 1610
rect 1695 1667 1895 1677
rect 1695 1611 1710 1667
rect 1766 1611 1820 1667
rect 1876 1611 1895 1667
rect 1695 1600 1895 1611
rect 3655 1667 3855 1677
rect 3655 1611 3674 1667
rect 3730 1611 3784 1667
rect 3840 1611 3855 1667
rect 3655 1600 3855 1611
rect 3935 1666 4135 1677
rect 3935 1610 3955 1666
rect 4011 1610 4065 1666
rect 4121 1610 4135 1666
rect 3935 1600 4135 1610
rect 4495 1667 4695 1677
rect 4495 1611 4516 1667
rect 4572 1611 4626 1667
rect 4682 1611 4695 1667
rect 4495 1600 4695 1611
rect 1467 1372 1545 1600
rect 857 1364 1054 1369
rect 857 1308 870 1364
rect 926 1308 980 1364
rect 1036 1308 1054 1364
rect 857 1303 1054 1308
rect 1415 1367 1612 1372
rect 1415 1311 1428 1367
rect 1484 1311 1538 1367
rect 1594 1311 1612 1367
rect 1415 1306 1612 1311
rect 2255 1353 2455 1368
rect 2255 1297 2267 1353
rect 2323 1297 2377 1353
rect 2433 1297 2455 1353
rect 2255 1291 2455 1297
rect 3095 1353 3295 1368
rect 3095 1297 3117 1353
rect 3173 1297 3227 1353
rect 3283 1297 3295 1353
rect 3095 1291 3295 1297
rect 2255 1287 2323 1291
rect 3227 1287 3295 1291
rect 2255 1247 2321 1287
rect -519 1183 289 1188
rect -519 1138 105 1183
rect -580 1127 105 1138
rect 161 1127 215 1183
rect 271 1127 289 1183
rect 603 1181 2321 1247
rect 3229 1247 3295 1287
rect 4881 1247 4947 2596
rect 3229 1181 4947 1247
rect 5083 2657 5535 2662
rect 5083 2601 5347 2657
rect 5403 2601 5455 2657
rect 5511 2601 5535 2657
rect 5083 2596 5535 2601
rect 5083 1247 5149 2596
rect 5335 2594 5535 2596
rect 5895 2664 6095 2672
rect 5895 2608 5908 2664
rect 5964 2608 6018 2664
rect 6074 2608 6095 2664
rect 5895 2595 6095 2608
rect 6175 2661 6375 2672
rect 6175 2605 6189 2661
rect 6245 2605 6299 2661
rect 6355 2605 6375 2661
rect 6175 2595 6375 2605
rect 6735 2658 6935 2672
rect 6735 2602 6747 2658
rect 6803 2602 6857 2658
rect 6913 2602 6935 2658
rect 6735 2595 6935 2602
rect 5345 2591 5401 2594
rect 5730 2536 5922 2539
rect 5730 2480 5742 2536
rect 5798 2480 5852 2536
rect 5908 2480 5922 2536
rect 5730 2477 5922 2480
rect 5319 2471 5509 2475
rect 5319 2415 5331 2471
rect 5387 2415 5441 2471
rect 5497 2415 5509 2471
rect 5319 2410 5509 2415
rect 5331 2409 5509 2410
rect 5736 2329 5802 2477
rect 5335 2315 5535 2327
rect 5335 2259 5350 2315
rect 5406 2259 5460 2315
rect 5516 2259 5535 2315
rect 5335 2249 5535 2259
rect 5615 2321 5815 2329
rect 5615 2265 5630 2321
rect 5686 2265 5740 2321
rect 5796 2265 5815 2321
rect 5615 2252 5815 2265
rect 6292 2271 6364 2595
rect 7022 2329 7088 3023
rect 7422 2329 7488 3023
rect 8265 2981 8321 2982
rect 8135 2972 8335 2981
rect 8135 2916 8155 2972
rect 8211 2916 8265 2972
rect 8321 2916 8335 2972
rect 8135 2904 8335 2916
rect 8546 2672 8602 2674
rect 7575 2658 7775 2672
rect 7575 2602 7597 2658
rect 7653 2602 7707 2658
rect 7763 2602 7775 2658
rect 7575 2595 7775 2602
rect 8135 2661 8335 2672
rect 8135 2605 8155 2661
rect 8211 2605 8265 2661
rect 8321 2605 8335 2661
rect 8135 2595 8335 2605
rect 8415 2664 8615 2672
rect 8415 2608 8436 2664
rect 8492 2608 8546 2664
rect 8602 2608 8615 2664
rect 8415 2595 8615 2608
rect 8975 2662 9175 2671
rect 8975 2657 9427 2662
rect 8975 2601 8999 2657
rect 9055 2601 9107 2657
rect 9163 2601 9427 2657
rect 8975 2596 9427 2601
rect 6735 2314 6935 2328
rect 6735 2271 6749 2314
rect 6292 2258 6749 2271
rect 6805 2258 6859 2314
rect 6915 2258 6935 2314
rect 6292 2248 6935 2258
rect 7015 2316 7215 2329
rect 7015 2260 7028 2316
rect 7084 2260 7138 2316
rect 7194 2260 7215 2316
rect 7015 2252 7215 2260
rect 7295 2316 7495 2329
rect 7295 2260 7316 2316
rect 7372 2260 7426 2316
rect 7482 2260 7495 2316
rect 7295 2252 7495 2260
rect 7575 2314 7775 2328
rect 7575 2258 7595 2314
rect 7651 2258 7705 2314
rect 7761 2271 7775 2314
rect 8146 2271 8218 2595
rect 8975 2594 9175 2596
rect 9109 2591 9165 2594
rect 8588 2536 8780 2539
rect 8588 2480 8602 2536
rect 8658 2480 8712 2536
rect 8768 2480 8780 2536
rect 8588 2477 8780 2480
rect 8708 2329 8774 2477
rect 8999 2470 9189 2475
rect 8999 2414 9011 2470
rect 9067 2414 9121 2470
rect 9177 2414 9189 2470
rect 8999 2409 9189 2414
rect 7761 2258 8218 2271
rect 7028 2250 7084 2252
rect 7426 2250 7482 2252
rect 7575 2248 8218 2258
rect 8695 2321 8895 2329
rect 8695 2265 8714 2321
rect 8770 2265 8824 2321
rect 8880 2265 8895 2321
rect 8695 2252 8895 2265
rect 8975 2315 9175 2327
rect 8975 2259 8994 2315
rect 9050 2259 9104 2315
rect 9160 2259 9175 2315
rect 8975 2249 9175 2259
rect 6292 2199 6850 2248
rect 7660 2199 8218 2248
rect 5335 2009 5535 2019
rect 5335 1953 5348 2009
rect 5404 1953 5458 2009
rect 5514 1953 5535 2009
rect 5335 1942 5535 1953
rect 5615 2010 5815 2020
rect 5615 1954 5628 2010
rect 5684 1954 5738 2010
rect 5794 1954 5815 2010
rect 5615 1943 5815 1954
rect 6735 2008 6935 2020
rect 6735 1952 6750 2008
rect 6806 1952 6860 2008
rect 6916 1952 6935 2008
rect 5736 1786 5802 1943
rect 6735 1942 6935 1952
rect 7575 2008 7775 2020
rect 7575 1952 7594 2008
rect 7650 1952 7704 2008
rect 7760 1952 7775 2008
rect 7575 1942 7775 1952
rect 8695 2010 8895 2020
rect 8695 1954 8716 2010
rect 8772 1954 8826 2010
rect 8882 1954 8895 2010
rect 8695 1943 8895 1954
rect 8975 2009 9175 2019
rect 8975 1953 8996 2009
rect 9052 1953 9106 2009
rect 9162 1953 9175 2009
rect 6752 1820 6820 1942
rect 5729 1781 5809 1786
rect 5729 1725 5741 1781
rect 5797 1725 5809 1781
rect 5729 1719 5809 1725
rect 6257 1752 6820 1820
rect 7690 1820 7758 1942
rect 7690 1752 8253 1820
rect 8708 1786 8774 1943
rect 8975 1942 9175 1953
rect 6257 1677 6325 1752
rect 8185 1677 8253 1752
rect 8701 1781 8781 1786
rect 8701 1725 8713 1781
rect 8769 1725 8781 1781
rect 8701 1719 8781 1725
rect 5335 1667 5535 1677
rect 5335 1611 5348 1667
rect 5404 1611 5458 1667
rect 5514 1611 5535 1667
rect 5335 1600 5535 1611
rect 5895 1666 6095 1677
rect 5895 1610 5909 1666
rect 5965 1610 6019 1666
rect 6075 1610 6095 1666
rect 5895 1600 6095 1610
rect 6175 1667 6375 1677
rect 6175 1611 6190 1667
rect 6246 1611 6300 1667
rect 6356 1611 6375 1667
rect 6175 1600 6375 1611
rect 8135 1667 8335 1677
rect 8135 1611 8154 1667
rect 8210 1611 8264 1667
rect 8320 1611 8335 1667
rect 8135 1600 8335 1611
rect 8415 1666 8615 1677
rect 8415 1610 8435 1666
rect 8491 1610 8545 1666
rect 8601 1610 8615 1666
rect 8415 1600 8615 1610
rect 8975 1667 9175 1677
rect 8975 1611 8996 1667
rect 9052 1611 9106 1667
rect 9162 1611 9175 1667
rect 8975 1600 9175 1611
rect 6735 1353 6935 1368
rect 6735 1297 6747 1353
rect 6803 1297 6857 1353
rect 6913 1297 6935 1353
rect 6735 1291 6935 1297
rect 7575 1353 7775 1368
rect 7575 1297 7597 1353
rect 7653 1297 7707 1353
rect 7763 1297 7775 1353
rect 7575 1291 7775 1297
rect 6735 1287 6803 1291
rect 7707 1287 7775 1291
rect 6735 1247 6801 1287
rect 5083 1181 6801 1247
rect 7709 1247 7775 1287
rect 9361 1247 9427 2596
rect 9700 2538 9897 2543
rect 9700 2482 9713 2538
rect 9771 2482 9823 2538
rect 9881 2482 9897 2538
rect 9700 2477 9897 2482
rect 10121 2323 10184 2338
rect 10121 2267 10126 2323
rect 10182 2267 10184 2323
rect 10121 2213 10184 2267
rect 10121 2207 10126 2213
rect 9485 2202 10126 2207
rect 9485 2146 9503 2202
rect 9559 2146 9613 2202
rect 9669 2157 10126 2202
rect 10182 2157 10184 2213
rect 9669 2146 10184 2157
rect 9485 2141 10184 2146
rect 10121 2140 10184 2141
rect 9484 1780 9681 1785
rect 9484 1724 9502 1780
rect 9558 1724 9612 1780
rect 9668 1724 9681 1780
rect 9484 1719 9681 1724
rect 9555 1458 9621 1719
rect 10231 1678 10294 1693
rect 10231 1622 10236 1678
rect 10292 1622 10294 1678
rect 10231 1568 10294 1622
rect 10231 1561 10236 1568
rect 9733 1556 10236 1561
rect 9733 1500 9751 1556
rect 9807 1500 9861 1556
rect 9917 1512 10236 1556
rect 10292 1512 10294 1568
rect 9917 1500 10294 1512
rect 9733 1496 10294 1500
rect 9733 1495 10292 1496
rect 10360 1476 10423 1491
rect 9483 1453 9680 1458
rect 9483 1397 9501 1453
rect 9557 1397 9611 1453
rect 9667 1397 9680 1453
rect 9483 1392 9680 1397
rect 9614 1359 9680 1392
rect 10360 1420 10365 1476
rect 10421 1420 10423 1476
rect 10360 1366 10423 1420
rect 10360 1359 10365 1366
rect 9614 1310 10365 1359
rect 10421 1310 10423 1366
rect 9614 1293 10423 1310
rect 10479 1305 10542 1320
rect 7709 1181 9427 1247
rect 10479 1249 10484 1305
rect 10540 1249 10542 1305
rect 10479 1195 10542 1249
rect 10479 1188 10484 1195
rect 9713 1183 10484 1188
rect -580 1122 289 1127
rect 9713 1127 9731 1183
rect 9787 1127 9841 1183
rect 9897 1139 10484 1183
rect 10540 1139 10542 1195
rect 9897 1127 10542 1139
rect 9713 1123 10542 1127
rect 9713 1122 10540 1123
<< via2 >>
rect 1709 5345 1765 5401
rect 1819 5345 1875 5401
rect 109 4575 165 4631
rect 219 4575 275 4631
rect 101 3929 157 3985
rect 211 3929 267 3985
rect 1428 5037 1484 5093
rect 1538 5037 1594 5093
rect 2267 5031 2323 5087
rect 2377 5031 2433 5087
rect 851 4844 907 4900
rect 961 4844 1017 4900
rect 870 4688 926 4744
rect 980 4688 1036 4744
rect 3675 5345 3731 5401
rect 3785 5345 3841 5401
rect 6189 5345 6245 5401
rect 6299 5345 6355 5401
rect 3117 5031 3173 5087
rect 3227 5031 3283 5087
rect 3956 5037 4012 5093
rect 4066 5037 4122 5093
rect 4531 4843 4587 4899
rect 4641 4843 4697 4899
rect 868 4382 924 4438
rect 978 4382 1034 4438
rect 4514 4688 4570 4744
rect 4624 4688 4680 4744
rect 4516 4382 4572 4438
rect 4626 4382 4682 4438
rect 868 4040 924 4096
rect 978 4040 1034 4096
rect 1429 4039 1485 4095
rect 1539 4039 1595 4095
rect 3955 4039 4011 4095
rect 4065 4039 4121 4095
rect 4516 4040 4572 4096
rect 4626 4040 4682 4096
rect 870 3737 926 3793
rect 980 3737 1036 3793
rect 1428 3739 1484 3795
rect 1538 3739 1594 3795
rect 5908 5037 5964 5093
rect 6018 5037 6074 5093
rect 6747 5031 6803 5087
rect 6857 5031 6913 5087
rect 5331 4844 5387 4900
rect 5441 4844 5497 4900
rect 5350 4688 5406 4744
rect 5460 4688 5516 4744
rect 8155 5345 8211 5401
rect 8265 5345 8321 5401
rect 7597 5031 7653 5087
rect 7707 5031 7763 5087
rect 8436 5037 8492 5093
rect 8546 5037 8602 5093
rect 9011 4843 9067 4899
rect 9121 4843 9177 4899
rect 8994 4688 9050 4744
rect 9104 4688 9160 4744
rect 5348 4382 5404 4438
rect 5458 4382 5514 4438
rect 8996 4382 9052 4438
rect 9106 4382 9162 4438
rect 5348 4040 5404 4096
rect 5458 4040 5514 4096
rect 5909 4039 5965 4095
rect 6019 4039 6075 4095
rect 8435 4039 8491 4095
rect 8545 4039 8601 4095
rect 8996 4040 9052 4096
rect 9106 4040 9162 4096
rect 9713 4911 9769 4967
rect 9823 4911 9879 4967
rect 9751 3929 9807 3985
rect 9861 3929 9917 3985
rect 1709 2916 1765 2972
rect 1819 2916 1875 2972
rect 109 2146 165 2202
rect 219 2146 275 2202
rect 101 1500 157 1556
rect 211 1500 267 1556
rect 1428 2608 1484 2664
rect 1538 2608 1594 2664
rect 2267 2602 2323 2658
rect 2377 2602 2433 2658
rect 851 2415 907 2471
rect 961 2415 1017 2471
rect 870 2259 926 2315
rect 980 2259 1036 2315
rect 3675 2916 3731 2972
rect 3785 2916 3841 2972
rect 6189 2916 6245 2972
rect 6299 2916 6355 2972
rect 3117 2602 3173 2658
rect 3227 2602 3283 2658
rect 3956 2608 4012 2664
rect 4066 2608 4122 2664
rect 4531 2414 4587 2470
rect 4641 2414 4697 2470
rect 868 1953 924 2009
rect 978 1953 1034 2009
rect 4514 2259 4570 2315
rect 4624 2259 4680 2315
rect 4516 1953 4572 2009
rect 4626 1953 4682 2009
rect 868 1611 924 1667
rect 978 1611 1034 1667
rect 1429 1610 1485 1666
rect 1539 1610 1595 1666
rect 3955 1610 4011 1666
rect 4065 1610 4121 1666
rect 4516 1611 4572 1667
rect 4626 1611 4682 1667
rect 870 1308 926 1364
rect 980 1308 1036 1364
rect 1428 1311 1484 1367
rect 1538 1311 1594 1367
rect 5908 2608 5964 2664
rect 6018 2608 6074 2664
rect 6747 2602 6803 2658
rect 6857 2602 6913 2658
rect 5331 2415 5387 2471
rect 5441 2415 5497 2471
rect 5350 2259 5406 2315
rect 5460 2259 5516 2315
rect 8155 2916 8211 2972
rect 8265 2916 8321 2972
rect 7597 2602 7653 2658
rect 7707 2602 7763 2658
rect 8436 2608 8492 2664
rect 8546 2608 8602 2664
rect 9011 2414 9067 2470
rect 9121 2414 9177 2470
rect 8994 2259 9050 2315
rect 9104 2259 9160 2315
rect 5348 1953 5404 2009
rect 5458 1953 5514 2009
rect 8996 1953 9052 2009
rect 9106 1953 9162 2009
rect 5348 1611 5404 1667
rect 5458 1611 5514 1667
rect 5909 1610 5965 1666
rect 6019 1610 6075 1666
rect 8435 1610 8491 1666
rect 8545 1610 8601 1666
rect 8996 1611 9052 1667
rect 9106 1611 9162 1667
rect 9713 2482 9769 2538
rect 9823 2482 9879 2538
rect 9751 1500 9807 1556
rect 9861 1500 9917 1556
<< metal3 >>
rect 1695 5401 1895 5410
rect 1695 5345 1709 5401
rect 1765 5345 1819 5401
rect 1875 5345 1895 5401
rect 1695 5333 1895 5345
rect 3655 5401 3855 5410
rect 3655 5345 3675 5401
rect 3731 5345 3785 5401
rect 3841 5345 3855 5401
rect 3655 5333 3855 5345
rect 6175 5401 6375 5410
rect 6175 5345 6189 5401
rect 6245 5345 6299 5401
rect 6355 5345 6375 5401
rect 6175 5333 6375 5345
rect 8135 5401 8335 5410
rect 8135 5345 8155 5401
rect 8211 5345 8265 5401
rect 8321 5345 8335 5401
rect 8135 5333 8335 5345
rect 1415 5093 1615 5101
rect 1415 5037 1428 5093
rect 1484 5037 1538 5093
rect 1594 5037 1615 5093
rect 1415 5024 1615 5037
rect 1460 4904 1526 5024
rect 713 4900 1526 4904
rect 713 4844 851 4900
rect 907 4844 961 4900
rect 1017 4844 1526 4900
rect 713 4838 1526 4844
rect 855 4744 1055 4756
rect 855 4688 870 4744
rect 926 4688 980 4744
rect 1036 4710 1055 4744
rect 1036 4688 1057 4710
rect 855 4678 1057 4688
rect 932 4668 1057 4678
rect 1708 4668 1772 5333
rect 2255 5087 2455 5101
rect 2255 5031 2267 5087
rect 2323 5031 2377 5087
rect 2433 5031 2455 5087
rect 2255 5024 2455 5031
rect 3095 5087 3295 5101
rect 3095 5031 3117 5087
rect 3173 5031 3227 5087
rect 3283 5031 3295 5087
rect 3095 5024 3295 5031
rect 96 4631 293 4636
rect 96 4575 109 4631
rect 165 4575 219 4631
rect 275 4575 293 4631
rect 96 4570 293 4575
rect 932 4604 1772 4668
rect 160 3990 226 4570
rect 932 4448 1016 4604
rect 855 4438 1055 4448
rect 855 4382 868 4438
rect 924 4382 978 4438
rect 1034 4382 1055 4438
rect 855 4371 1055 4382
rect 982 4286 1055 4371
rect 982 4213 1514 4286
rect 1441 4106 1514 4213
rect 855 4096 1055 4106
rect 855 4040 868 4096
rect 924 4040 978 4096
rect 1034 4040 1055 4096
rect 855 4029 1055 4040
rect 1415 4095 1615 4106
rect 1415 4039 1429 4095
rect 1485 4039 1539 4095
rect 1595 4039 1615 4095
rect 1415 4029 1615 4039
rect 88 3985 285 3990
rect 88 3929 101 3985
rect 157 3929 211 3985
rect 267 3929 285 3985
rect 88 3924 285 3929
rect 954 3973 1055 4029
rect 2352 3973 2418 5024
rect 954 3907 2418 3973
rect 3132 3973 3198 5024
rect 3778 4668 3842 5333
rect 3935 5093 4135 5101
rect 3935 5037 3956 5093
rect 4012 5037 4066 5093
rect 4122 5037 4135 5093
rect 3935 5024 4135 5037
rect 5895 5093 6095 5101
rect 5895 5037 5908 5093
rect 5964 5037 6018 5093
rect 6074 5037 6095 5093
rect 5895 5024 6095 5037
rect 4024 4904 4090 5024
rect 5940 4904 6006 5024
rect 4024 4899 4709 4904
rect 4024 4843 4531 4899
rect 4587 4843 4641 4899
rect 4697 4843 4709 4899
rect 4024 4838 4709 4843
rect 5193 4900 6006 4904
rect 5193 4844 5331 4900
rect 5387 4844 5441 4900
rect 5497 4844 6006 4900
rect 5193 4838 6006 4844
rect 4495 4744 4695 4756
rect 4495 4688 4514 4744
rect 4570 4688 4624 4744
rect 4680 4688 4695 4744
rect 4495 4678 4695 4688
rect 5335 4744 5535 4756
rect 5335 4688 5350 4744
rect 5406 4688 5460 4744
rect 5516 4688 5535 4744
rect 5335 4678 5535 4688
rect 4495 4668 4607 4678
rect 3778 4604 4607 4668
rect 5420 4668 5535 4678
rect 6188 4668 6252 5333
rect 6735 5087 6935 5101
rect 6735 5031 6747 5087
rect 6803 5031 6857 5087
rect 6913 5031 6935 5087
rect 6735 5024 6935 5031
rect 7575 5087 7775 5101
rect 7575 5031 7597 5087
rect 7653 5031 7707 5087
rect 7763 5031 7775 5087
rect 7575 5024 7775 5031
rect 5420 4604 6252 4668
rect 4495 4438 4695 4448
rect 4495 4382 4516 4438
rect 4572 4382 4626 4438
rect 4682 4382 4695 4438
rect 4495 4371 4695 4382
rect 5335 4438 5535 4448
rect 5335 4382 5348 4438
rect 5404 4382 5458 4438
rect 5514 4382 5535 4438
rect 5335 4371 5535 4382
rect 4495 4286 4568 4371
rect 4036 4213 4568 4286
rect 5462 4286 5535 4371
rect 5462 4213 5994 4286
rect 4036 4106 4109 4213
rect 5921 4106 5994 4213
rect 3935 4095 4135 4106
rect 3935 4039 3955 4095
rect 4011 4039 4065 4095
rect 4121 4039 4135 4095
rect 3935 4029 4135 4039
rect 4495 4096 4695 4106
rect 4495 4040 4516 4096
rect 4572 4040 4626 4096
rect 4682 4040 4695 4096
rect 4495 4029 4695 4040
rect 5335 4096 5535 4106
rect 5335 4040 5348 4096
rect 5404 4040 5458 4096
rect 5514 4040 5535 4096
rect 5335 4029 5535 4040
rect 5895 4095 6095 4106
rect 5895 4039 5909 4095
rect 5965 4039 6019 4095
rect 6075 4039 6095 4095
rect 5895 4029 6095 4039
rect 4495 3973 4596 4029
rect 3132 3907 4596 3973
rect 5434 3973 5535 4029
rect 6832 3973 6898 5024
rect 5434 3907 6898 3973
rect 7612 3973 7678 5024
rect 8258 4668 8322 5333
rect 8415 5093 8615 5101
rect 8415 5037 8436 5093
rect 8492 5037 8546 5093
rect 8602 5037 8615 5093
rect 8415 5024 8615 5037
rect 8504 4904 8570 5024
rect 9700 4967 9897 4972
rect 9700 4911 9713 4967
rect 9769 4911 9823 4967
rect 9879 4911 9897 4967
rect 9700 4906 9897 4911
rect 8504 4899 9189 4904
rect 8504 4843 9011 4899
rect 9067 4843 9121 4899
rect 9177 4843 9189 4899
rect 8504 4838 9189 4843
rect 8975 4744 9175 4756
rect 8975 4688 8994 4744
rect 9050 4688 9104 4744
rect 9160 4688 9175 4744
rect 8975 4678 9175 4688
rect 8975 4668 9087 4678
rect 8258 4604 9087 4668
rect 8975 4438 9175 4448
rect 8975 4382 8996 4438
rect 9052 4382 9106 4438
rect 9162 4382 9175 4438
rect 8975 4371 9175 4382
rect 8975 4286 9048 4371
rect 8516 4213 9048 4286
rect 8516 4106 8589 4213
rect 8415 4095 8615 4106
rect 8415 4039 8435 4095
rect 8491 4039 8545 4095
rect 8601 4039 8615 4095
rect 8415 4029 8615 4039
rect 8975 4096 9175 4106
rect 8975 4040 8996 4096
rect 9052 4040 9106 4096
rect 9162 4040 9175 4096
rect 8975 4029 9175 4040
rect 8975 3973 9076 4029
rect 9801 3990 9867 4906
rect 7612 3907 9076 3973
rect 9738 3985 9935 3990
rect 9738 3929 9751 3985
rect 9807 3929 9861 3985
rect 9917 3929 9935 3985
rect 9738 3924 9935 3929
rect 954 3798 1055 3907
rect 857 3793 1055 3798
rect 857 3737 870 3793
rect 926 3737 980 3793
rect 1036 3769 1055 3793
rect 1415 3795 1612 3800
rect 1036 3737 1054 3769
rect 857 3732 1054 3737
rect 1415 3739 1428 3795
rect 1484 3739 1538 3795
rect 1594 3739 1612 3795
rect 1415 3734 1612 3739
rect 1695 2972 1895 2981
rect 1695 2916 1709 2972
rect 1765 2916 1819 2972
rect 1875 2916 1895 2972
rect 1695 2904 1895 2916
rect 3655 2972 3855 2981
rect 3655 2916 3675 2972
rect 3731 2916 3785 2972
rect 3841 2916 3855 2972
rect 3655 2904 3855 2916
rect 6175 2972 6375 2981
rect 6175 2916 6189 2972
rect 6245 2916 6299 2972
rect 6355 2916 6375 2972
rect 6175 2904 6375 2916
rect 8135 2972 8335 2981
rect 8135 2916 8155 2972
rect 8211 2916 8265 2972
rect 8321 2916 8335 2972
rect 8135 2904 8335 2916
rect 1415 2664 1615 2672
rect 1415 2608 1428 2664
rect 1484 2608 1538 2664
rect 1594 2608 1615 2664
rect 1415 2595 1615 2608
rect 1460 2475 1526 2595
rect 713 2471 1526 2475
rect 713 2415 851 2471
rect 907 2415 961 2471
rect 1017 2415 1526 2471
rect 713 2409 1526 2415
rect 855 2315 1055 2327
rect 855 2259 870 2315
rect 926 2259 980 2315
rect 1036 2259 1055 2315
rect 855 2249 1055 2259
rect 924 2239 1055 2249
rect 1708 2239 1772 2904
rect 2255 2658 2455 2672
rect 2255 2602 2267 2658
rect 2323 2602 2377 2658
rect 2433 2602 2455 2658
rect 2255 2595 2455 2602
rect 3095 2658 3295 2672
rect 3095 2602 3117 2658
rect 3173 2602 3227 2658
rect 3283 2602 3295 2658
rect 3095 2595 3295 2602
rect 96 2202 293 2207
rect 96 2146 109 2202
rect 165 2146 219 2202
rect 275 2146 293 2202
rect 924 2175 1772 2239
rect 96 2141 293 2146
rect 160 1561 226 2141
rect 945 2019 1029 2175
rect 855 2009 1055 2019
rect 855 1953 868 2009
rect 924 1953 978 2009
rect 1034 1953 1055 2009
rect 855 1942 1055 1953
rect 982 1857 1055 1942
rect 982 1784 1514 1857
rect 1441 1677 1514 1784
rect 855 1667 1055 1677
rect 855 1611 868 1667
rect 924 1611 978 1667
rect 1034 1611 1055 1667
rect 855 1600 1055 1611
rect 1415 1666 1615 1677
rect 1415 1610 1429 1666
rect 1485 1610 1539 1666
rect 1595 1610 1615 1666
rect 1415 1600 1615 1610
rect 88 1556 285 1561
rect 88 1500 101 1556
rect 157 1500 211 1556
rect 267 1500 285 1556
rect 88 1495 285 1500
rect 954 1544 1055 1600
rect 2352 1544 2418 2595
rect 954 1478 2418 1544
rect 3132 1544 3198 2595
rect 3778 2239 3842 2904
rect 3935 2664 4135 2672
rect 3935 2608 3956 2664
rect 4012 2608 4066 2664
rect 4122 2608 4135 2664
rect 3935 2595 4135 2608
rect 5895 2664 6095 2672
rect 5895 2608 5908 2664
rect 5964 2608 6018 2664
rect 6074 2608 6095 2664
rect 5895 2595 6095 2608
rect 4024 2475 4090 2595
rect 5940 2475 6006 2595
rect 4024 2470 4709 2475
rect 4024 2414 4531 2470
rect 4587 2414 4641 2470
rect 4697 2414 4709 2470
rect 4024 2409 4709 2414
rect 5193 2471 6006 2475
rect 5193 2415 5331 2471
rect 5387 2415 5441 2471
rect 5497 2415 6006 2471
rect 5193 2409 6006 2415
rect 4495 2315 4695 2327
rect 4495 2259 4514 2315
rect 4570 2259 4624 2315
rect 4680 2259 4695 2315
rect 4495 2249 4695 2259
rect 5335 2315 5535 2327
rect 5335 2259 5350 2315
rect 5406 2259 5460 2315
rect 5516 2259 5535 2315
rect 5335 2249 5535 2259
rect 4495 2239 4607 2249
rect 3778 2175 4607 2239
rect 5423 2239 5535 2249
rect 6188 2239 6252 2904
rect 6735 2658 6935 2672
rect 6735 2602 6747 2658
rect 6803 2602 6857 2658
rect 6913 2602 6935 2658
rect 6735 2595 6935 2602
rect 7575 2658 7775 2672
rect 7575 2602 7597 2658
rect 7653 2602 7707 2658
rect 7763 2602 7775 2658
rect 7575 2595 7775 2602
rect 5423 2175 6252 2239
rect 4495 2009 4695 2019
rect 4495 1953 4516 2009
rect 4572 1953 4626 2009
rect 4682 1953 4695 2009
rect 4495 1942 4695 1953
rect 5335 2009 5535 2019
rect 5335 1953 5348 2009
rect 5404 1953 5458 2009
rect 5514 1953 5535 2009
rect 5335 1942 5535 1953
rect 4495 1857 4568 1942
rect 4036 1784 4568 1857
rect 5462 1857 5535 1942
rect 5462 1784 5994 1857
rect 4036 1677 4109 1784
rect 5921 1677 5994 1784
rect 3935 1666 4135 1677
rect 3935 1610 3955 1666
rect 4011 1610 4065 1666
rect 4121 1610 4135 1666
rect 3935 1600 4135 1610
rect 4495 1667 4695 1677
rect 4495 1611 4516 1667
rect 4572 1611 4626 1667
rect 4682 1611 4695 1667
rect 4495 1600 4695 1611
rect 5335 1667 5535 1677
rect 5335 1611 5348 1667
rect 5404 1611 5458 1667
rect 5514 1611 5535 1667
rect 5335 1600 5535 1611
rect 5895 1666 6095 1677
rect 5895 1610 5909 1666
rect 5965 1610 6019 1666
rect 6075 1610 6095 1666
rect 5895 1600 6095 1610
rect 4495 1544 4596 1600
rect 3132 1478 4596 1544
rect 5434 1544 5535 1600
rect 6832 1544 6898 2595
rect 5434 1478 6898 1544
rect 7612 1544 7678 2595
rect 8258 2239 8322 2904
rect 8415 2664 8615 2672
rect 8415 2608 8436 2664
rect 8492 2608 8546 2664
rect 8602 2608 8615 2664
rect 8415 2595 8615 2608
rect 8504 2475 8570 2595
rect 9700 2538 9897 2543
rect 9700 2482 9713 2538
rect 9769 2482 9823 2538
rect 9879 2482 9897 2538
rect 9700 2477 9897 2482
rect 8504 2470 9189 2475
rect 8504 2414 9011 2470
rect 9067 2414 9121 2470
rect 9177 2414 9189 2470
rect 8504 2409 9189 2414
rect 8975 2315 9175 2327
rect 8975 2259 8994 2315
rect 9050 2259 9104 2315
rect 9160 2259 9175 2315
rect 8975 2249 9175 2259
rect 8975 2239 9087 2249
rect 8258 2175 9087 2239
rect 8975 2009 9175 2019
rect 8975 1953 8996 2009
rect 9052 1953 9106 2009
rect 9162 1953 9175 2009
rect 8975 1942 9175 1953
rect 8975 1857 9048 1942
rect 8516 1784 9048 1857
rect 8516 1677 8589 1784
rect 8415 1666 8615 1677
rect 8415 1610 8435 1666
rect 8491 1610 8545 1666
rect 8601 1610 8615 1666
rect 8415 1600 8615 1610
rect 8975 1667 9175 1677
rect 8975 1611 8996 1667
rect 9052 1611 9106 1667
rect 9162 1611 9175 1667
rect 8975 1600 9175 1611
rect 8975 1544 9076 1600
rect 9801 1561 9867 2477
rect 7612 1478 9076 1544
rect 9738 1556 9935 1561
rect 9738 1500 9751 1556
rect 9807 1500 9861 1556
rect 9917 1500 9935 1556
rect 9738 1495 9935 1500
rect 954 1369 1055 1478
rect 857 1364 1055 1369
rect 857 1308 870 1364
rect 926 1308 980 1364
rect 1036 1340 1055 1364
rect 1415 1367 1612 1372
rect 1036 1308 1054 1340
rect 857 1303 1054 1308
rect 1415 1311 1428 1367
rect 1484 1311 1538 1367
rect 1594 1311 1612 1367
rect 1415 1306 1612 1311
<< labels >>
flabel metal2 -186 4177 -186 4177 0 FreeSans 800 0 0 0 E
port 7 nsew
flabel metal2 10122 3943 10122 3943 0 FreeSans 800 0 0 0 D
port 13 nsew
flabel metal2 10113 3748 10113 3748 0 FreeSans 800 0 0 0 F
port 12 nsew
flabel metal2 10126 3578 10126 3578 0 FreeSans 800 0 0 0 H
port 11 nsew
flabel via1 -207 4594 -207 4594 0 FreeSans 800 0 0 0 C
port 9 nsew
flabel metal2 -220 3582 -220 3582 0 FreeSans 800 0 0 0 G
port 5 nsew
flabel metal2 10292 4594 10292 4594 0 FreeSans 800 0 0 0 B
port 3 nsew
flabel metal2 -238 4290 -238 4290 0 FreeSans 800 0 0 0 A
port 0 nsew
flabel metal1 4655 5669 4655 5669 0 FreeSans 1280 0 0 0 VDD
port 15 nsew
<< end >>
