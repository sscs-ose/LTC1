magic
tech gf180mcuC
magscale 1 10
timestamp 1714537808
<< nwell >>
rect 1118 808 2091 1229
<< psubdiff >>
rect 1109 414 2140 430
rect 1109 361 1193 414
rect 1245 361 1354 414
rect 1406 361 1515 414
rect 1567 361 1676 414
rect 1728 361 1837 414
rect 1889 361 1998 414
rect 2050 361 2140 414
rect 1109 348 2140 361
<< nsubdiff >>
rect 1146 1189 1254 1204
rect 1146 1143 1159 1189
rect 1205 1159 1254 1189
rect 1205 1143 1219 1159
rect 1146 1106 1219 1143
<< psubdiffcont >>
rect 1193 361 1245 414
rect 1354 361 1406 414
rect 1515 361 1567 414
rect 1676 361 1728 414
rect 1837 361 1889 414
rect 1998 361 2050 414
<< nsubdiffcont >>
rect 1159 1143 1205 1189
<< polysilicon >>
rect 1325 878 1395 894
rect 1259 876 1395 878
rect 1499 876 1569 894
rect 1673 876 1743 894
rect 1847 876 1917 894
rect 1259 859 1917 876
rect 1259 809 1272 859
rect 1321 809 1917 859
rect 1259 801 1917 809
rect 1259 796 1395 801
rect 1325 761 1395 796
rect 1499 761 1569 801
rect 1673 761 1743 801
rect 1847 761 1917 801
<< polycontact >>
rect 1272 809 1321 859
<< metal1 >>
rect 1017 1250 2227 1332
rect 1017 430 1096 1250
rect 1146 1189 1254 1204
rect 1146 1143 1159 1189
rect 1205 1181 1254 1189
rect 1205 1143 1992 1181
rect 1146 1106 1992 1143
rect 1249 1105 1992 1106
rect 1249 1036 1296 1105
rect 1598 1036 1644 1105
rect 1946 1036 1992 1105
rect 1258 863 1329 866
rect 1154 859 1329 863
rect 1154 809 1272 859
rect 1321 809 1329 859
rect 1154 803 1329 809
rect 1258 798 1329 803
rect 1424 836 1470 940
rect 1772 836 1818 940
rect 1424 790 2004 836
rect 1424 715 1470 790
rect 1772 715 1818 790
rect 1250 430 1296 519
rect 1598 430 1644 521
rect 1946 430 1992 519
rect 2148 430 2227 1250
rect 1017 414 2227 430
rect 1017 361 1193 414
rect 1245 361 1354 414
rect 1406 361 1515 414
rect 1567 361 1676 414
rect 1728 361 1837 414
rect 1889 361 1998 414
rect 2050 361 2227 414
rect 1017 348 2227 361
use nmos_3p3_VDSZE6  nmos_3p3_VDSZE6_0
timestamp 1714126980
transform 1 0 1621 0 1 617
box -408 -168 408 168
use pmos_3p3_HDJZPK  pmos_3p3_HDJZPK_0
timestamp 1714126980
transform 1 0 1621 0 1 988
box -470 -180 470 180
<< labels >>
flabel metal1 1984 810 1984 810 0 FreeSans 640 0 0 0 OUT
port 1 nsew
flabel metal1 1163 825 1163 825 0 FreeSans 640 0 0 0 IN
port 0 nsew
flabel metal1 1270 450 1270 450 0 FreeSans 640 0 0 0 VSS
port 4 nsew
flabel metal1 1621 1140 1621 1140 0 FreeSans 640 0 0 0 VDD
port 3 nsew
<< end >>
