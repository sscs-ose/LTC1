magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2603 -2045 2603 2045
<< psubdiff >>
rect -603 23 603 45
rect -603 -23 -581 23
rect -535 -23 -457 23
rect -411 -23 -333 23
rect -287 -23 -209 23
rect -163 -23 -85 23
rect -39 -23 39 23
rect 85 -23 163 23
rect 209 -23 287 23
rect 333 -23 411 23
rect 457 -23 535 23
rect 581 -23 603 23
rect -603 -45 603 -23
<< psubdiffcont >>
rect -581 -23 -535 23
rect -457 -23 -411 23
rect -333 -23 -287 23
rect -209 -23 -163 23
rect -85 -23 -39 23
rect 39 -23 85 23
rect 163 -23 209 23
rect 287 -23 333 23
rect 411 -23 457 23
rect 535 -23 581 23
<< metal1 >>
rect -592 23 592 34
rect -592 -23 -581 23
rect -535 -23 -457 23
rect -411 -23 -333 23
rect -287 -23 -209 23
rect -163 -23 -85 23
rect -39 -23 39 23
rect 85 -23 163 23
rect 209 -23 287 23
rect 333 -23 411 23
rect 457 -23 535 23
rect 581 -23 592 23
rect -592 -34 592 -23
<< end >>
