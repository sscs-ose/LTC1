magic
tech gf180mcuC
magscale 1 10
timestamp 1691480513
<< error_p >>
rect -314 -23 -303 23
rect 246 -23 257 23
<< nwell >>
rect -402 -159 402 159
<< pmos >>
rect -224 -22 224 22
<< pdiff >>
rect -316 23 -244 36
rect -316 -23 -303 23
rect -257 22 -244 23
rect 244 23 316 36
rect 244 22 257 23
rect -257 -22 -224 22
rect 224 -22 257 22
rect -257 -23 -244 -22
rect -316 -36 -244 -23
rect 244 -23 257 -22
rect 303 -23 316 23
rect 244 -36 316 -23
<< pdiffc >>
rect -303 -23 -257 23
rect 257 -23 303 23
<< polysilicon >>
rect -224 22 224 66
rect -224 -66 224 -22
<< metal1 >>
rect -314 -23 -303 23
rect -257 -23 -246 23
rect 246 -23 257 23
rect 303 -23 314 23
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 0.220 l 2.24 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
