magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -8078 -2278 8078 2278
<< nwell >>
rect -6078 -278 6078 278
<< nsubdiff >>
rect -5995 173 5995 195
rect -5995 -173 -5973 173
rect 5973 -173 5995 173
rect -5995 -195 5995 -173
<< nsubdiffcont >>
rect -5973 -173 5973 173
<< metal1 >>
rect -5984 173 5984 184
rect -5984 -173 -5973 173
rect 5973 -173 5984 173
rect -5984 -184 5984 -173
<< end >>
