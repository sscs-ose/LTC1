** sch_path: /home/shahid/Videos/PGA_DECODER/xschem/pga_parallel_tb.sch
**.subckt pga_parallel_tb
V1 E GND 3
.save i(v1)
V2 VDD GND 3
.save i(v2)
x1 A B C D E F G H VDD pga_res_parallel
V3 H GND 0
.save i(v3)
**** begin user architecture code

.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice res_typical
* .lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice res_statistical



*vp p 0 0
*vm m 0 0
*vb b 0 3.3

.control
save all
*dc vp 0 3.3 0.01
dc v1 0.1 3.3 0.1
let i1 = i(v1)
let r  = maximum(v(A)/i(v1))
plot r
display all
*write res_sch_test.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  pga_res_parallel.sym # of pins=9
** sym_path: /home/shahid/Videos/PGA_DECODER/xschem/pga_res_parallel.sym
** sch_path: /home/shahid/Videos/PGA_DECODER/xschem/pga_res_parallel.sch
.subckt pga_res_parallel A B C D E F G H VDD
*.iopin VDD
*.iopin A
*.iopin B
*.iopin C
*.iopin D
*.iopin E
*.iopin F
*.iopin G
*.iopin H
XR1 net1 A VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR2 net2 net1 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR3 net2 net2 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR4 net2 net2 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR5 net6 net2 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR6 net3 net6 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR7 net4 net3 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR8 net7 net4 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR9 net5 net7 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR10 net78 net5 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR11 net8 net78 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR12 B net8 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR13 net9 B VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR14 net14 net9 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR15 net10 net14 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR16 net11 net10 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR17 net15 net11 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR18 net12 net15 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR19 net13 net12 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR20 C net13 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR25 net16 C VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR26 net22 net16 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR27 net17 net22 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR28 net18 net17 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR29 net23 net18 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR30 net19 net23 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR31 net20 net19 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR32 net24 net20 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR33 net21 net24 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR34 net79 net21 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR35 net25 net79 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR36 D net25 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR37 net26 D VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR38 net32 net26 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR39 net27 net32 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR40 net28 net27 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR41 net33 net28 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR42 net29 net33 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR43 net30 net29 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR44 net34 net30 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR45 net31 net34 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR46 net77 net31 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR47 net35 net77 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR48 net73 net35 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR49 net36 E VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR50 net36 net36 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR51 net37 net36 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR52 net38 net37 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR53 net42 net38 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR54 net39 net42 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR55 net40 net39 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR56 net43 net40 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR57 net41 net43 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR58 net80 net41 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR59 net44 net80 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR60 net70 net44 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR61 net45 F VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR62 net51 net45 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR63 net46 net51 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR64 net47 net46 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR65 net52 net47 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR66 net48 net52 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR67 net49 net48 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR68 net53 net49 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR69 net50 net53 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR70 net81 net50 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR71 net54 net81 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR72 G net54 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR73 G G VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR74 G G VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR75 net55 G VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR76 net56 net55 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR77 net60 net56 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR78 net57 net60 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR79 net58 net57 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR80 net61 net58 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR81 net59 net61 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR82 net82 net59 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR83 net62 net82 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR84 net83 net62 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR85 net63 net83 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR86 net68 net63 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR87 net64 net68 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR88 net65 net64 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR89 net69 net65 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR90 net66 net69 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR91 net67 net66 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR92 H net67 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR99 net71 net70 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR100 net72 net71 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR101 net76 net72 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR105 net74 net73 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR106 net75 net74 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR107 E net75 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR21 VDD VDD VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR22 VDD VDD VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR23 VDD VDD VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR24 VDD VDD VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR93 VDD VDD VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR94 VDD VDD VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR201 F net76 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR202 E E VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR95 net84 A VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR96 net85 net84 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR97 net85 net85 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR98 net85 net85 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR102 net89 net85 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR103 net86 net89 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR104 net87 net86 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR108 net90 net87 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR109 net88 net90 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR110 net161 net88 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR111 net91 net161 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR112 B net91 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR113 net92 B VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR114 net97 net92 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR115 net93 net97 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR116 net94 net93 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR117 net98 net94 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR118 net95 net98 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR119 net96 net95 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR120 C net96 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR121 net99 C VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR122 net105 net99 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR123 net100 net105 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR124 net101 net100 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR125 net106 net101 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR126 net102 net106 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR127 net103 net102 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR128 net107 net103 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR129 net104 net107 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR130 net162 net104 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR131 net108 net162 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR132 D net108 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR133 net109 D VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR134 net115 net109 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR135 net110 net115 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR136 net111 net110 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR137 net116 net111 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR138 net112 net116 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR139 net113 net112 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR140 net117 net113 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR141 net114 net117 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR142 net160 net114 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR143 net118 net160 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR144 net156 net118 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR145 net119 E VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR146 net119 net119 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR147 net120 net119 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR148 net121 net120 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR149 net125 net121 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR150 net122 net125 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR151 net123 net122 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR152 net126 net123 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR153 net124 net126 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR154 net163 net124 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR155 net127 net163 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR156 net153 net127 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR157 net128 F VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR158 net134 net128 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR159 net129 net134 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR160 net130 net129 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR161 net135 net130 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR162 net131 net135 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR163 net132 net131 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR164 net136 net132 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR165 net133 net136 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR166 net164 net133 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR167 net137 net164 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR168 G net137 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR169 G G VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR170 G G VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR171 net138 G VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR172 net139 net138 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR173 net143 net139 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR174 net140 net143 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR175 net141 net140 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR176 net144 net141 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR177 net142 net144 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR178 net165 net142 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR179 net145 net165 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR180 net166 net145 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR181 net146 net166 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR182 net151 net146 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR183 net147 net151 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR184 net148 net147 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR185 net152 net148 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR186 net149 net152 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR187 net150 net149 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR188 H net150 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR189 net154 net153 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR190 net155 net154 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR191 net159 net155 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR192 net157 net156 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR193 net158 net157 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR194 E net158 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR195 VDD VDD VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR196 VDD VDD VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR197 VDD VDD VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR198 VDD VDD VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR199 VDD VDD VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR200 VDD VDD VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR203 F net159 VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
XR204 E E VDD ppolyf_u r_width=1e-6 r_length=1e-6 m=1
.ends

.GLOBAL GND
.end
