magic
tech gf180mcuC
magscale 1 10
timestamp 1692811925
<< error_p >>
rect -34 313 -23 359
rect -34 -359 -23 -313
<< nwell >>
rect -285 -488 285 488
<< pmos >>
rect -35 -280 35 280
<< pdiff >>
rect -123 267 -35 280
rect -123 -267 -110 267
rect -64 -267 -35 267
rect -123 -280 -35 -267
rect 35 267 123 280
rect 35 -267 64 267
rect 110 -267 123 267
rect 35 -280 123 -267
<< pdiffc >>
rect -110 -267 -64 267
rect 64 -267 110 267
<< nsubdiff >>
rect -261 392 261 464
rect -261 348 -189 392
rect -261 -348 -248 348
rect -202 -348 -189 348
rect 189 348 261 392
rect -261 -392 -189 -348
rect 189 -348 202 348
rect 248 -348 261 348
rect 189 -392 261 -348
rect -261 -464 261 -392
<< nsubdiffcont >>
rect -248 -348 -202 348
rect 202 -348 248 348
<< polysilicon >>
rect -36 359 36 372
rect -36 313 -23 359
rect 23 313 36 359
rect -36 300 36 313
rect -35 280 35 300
rect -35 -300 35 -280
rect -36 -313 36 -300
rect -36 -359 -23 -313
rect 23 -359 36 -313
rect -36 -372 36 -359
<< polycontact >>
rect -23 313 23 359
rect -23 -359 23 -313
<< metal1 >>
rect -248 405 248 451
rect -248 348 -202 405
rect -34 313 -23 359
rect 23 313 34 359
rect 202 348 248 405
rect -110 267 -64 278
rect -110 -278 -64 -267
rect 64 267 110 278
rect 64 -278 110 -267
rect -248 -405 -202 -348
rect -34 -359 -23 -313
rect 23 -359 34 -313
rect 202 -405 248 -348
rect -248 -451 248 -405
<< properties >>
string FIXED_BBOX -225 -428 225 428
string gencell pmos_3p3
string library gf180mcu
string parameters w 2.8 l 0.35 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 1 compatible {pmos_3p3 pmos_6p0}
<< end >>
