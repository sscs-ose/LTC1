* NGSPICE file created from PGA_DECODER_magic_flat.ext - technology: gf180mcuC

.subckt pex_PGA_DECODER_magic VDD S6 VSS S4 S3 S5 S2 S1 A B C
X0 a_587_3452# AND_3_magic_3.A.t2 a_439_3441# VSS.t6 nfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
X1 VDD.t65 VDD.t63 VDD.t65 VDD.t64 pfet_03v3 ad=0 pd=0 as=89.8f ps=0.92u w=0.25u l=0.28u
X2 a_1091_5366# AND_3_magic_5.B.t2 a_587_5366# VSS.t0 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X3 a_439_2188# A.t0 a_587_2199# VSS.t52 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X4 a_439_2188# A.t1 VDD.t105 VDD.t13 pfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
X5 a_439_3441# C.t0 VDD.t81 VDD.t80 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X6 a_439_3441# B.t0 VDD.t21 VDD.t20 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X7 AND_3_magic_5.C C.t1 VSS.t34 VSS.t33 nfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X8 VDD a_439_3441# S4.t2 VDD.t115 pfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X9 VSS AND_3_magic_5.C.t2 a_1091_4113# VSS.t53 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X10 VDD B.t1 a_439_4102# VDD.t22 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X11 VDD A.t2 AND_3_magic_3.A VDD.t106 pfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
X12 a_400_841# B.t2 VDD.t26 VDD.t25 pfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
X13 a_252_1525# C.t2 VSS.t36 VSS.t35 nfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X14 S2 a_439_5355# VDD.t140 VDD.t70 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X15 a_252_1525# C.t3 a_400_841# VDD.t30 pfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X16 VDD AND_3_magic_5.C.t3 a_439_6016# VDD.t109 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X17 VDD A.t3 a_1333_1282# VDD.t135 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X18 AND_1.A a_252_1525# VDD.t29 VDD.t27 pfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X19 a_587_2199# A.t4 a_439_2188# VSS.t80 nfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
X20 VDD AND_3_magic_3.A.t3 a_439_3441# VDD.t15 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X21 a_587_4113# B.t3 a_1091_4113# VSS.t9 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X22 a_1091_5366# AND_3_magic_5.B.t3 a_587_5366# VSS.t26 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X23 a_587_5366# AND_3_magic_3.A.t4 a_439_5355# VSS.t5 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X24 S2 a_439_5355# VSS.t89 VSS.t31 nfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X25 VDD.t62 VDD.t61 VDD.t62 VDD.t39 pfet_03v3 ad=0 pd=0 as=89.8f ps=0.92u w=0.25u l=0.28u
X26 VSS B.t4 a_252_1525# VSS.t10 nfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
X27 a_439_4102# AND_3_magic_5.C.t4 VDD.t112 VDD.t34 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X28 VSS A.t5 a_1185_1271# VSS.t81 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X29 a_439_4102# B.t5 VDD.t141 VDD.t84 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X30 a_1091_6027# AND_3_magic_5.C.t5 VSS.t57 VSS.t56 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X31 VDD a_439_4102# S3.t2 VDD.t72 pfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X32 VDD C.t4 AND_3_magic_5.C VDD.t31 pfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
X33 a_1091_4113# B.t6 a_587_4113# VSS.t71 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X34 S1 a_439_6016# VDD.t79 VDD.t78 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X35 a_439_3441# AND_3_magic_3.A.t5 VDD.t14 VDD.t13 pfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
X36 a_439_5355# AND_3_magic_3.A.t6 a_587_5366# VSS.t4 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X37 VDD AND_3_magic_5.B.t4 a_439_5355# VDD.t22 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X38 a_1185_1271# AND_1.A a_1333_1282# VSS.t44 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X39 VDD AND_3_magic_3.A.t7 a_439_4102# VDD.t7 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X40 VSS AND_3_magic_5.C.t6 a_1091_6027# VSS.t58 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X41 VDD.t60 VDD.t58 VDD.t60 VDD.t59 pfet_03v3 ad=0 pd=0 as=89.8f ps=0.92u w=0.25u l=0.28u
X42 S6 a_1333_1282# VDD.t19 VDD.t18 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X43 a_400_841# B.t7 VDD.t142 VDD.t25 pfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
X44 a_587_5366# AND_3_magic_3.A.t8 a_439_5355# VSS.t3 nfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
X45 a_1091_4113# B.t8 a_587_4113# VSS.t72 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X46 a_587_4113# AND_3_magic_3.A.t9 a_439_4102# VSS.t2 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X47 a_1333_1282# AND_1.A a_1185_1271# VSS.t43 nfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
X48 a_439_5355# C.t5 VDD.t35 VDD.t34 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X49 S3 a_439_4102# VSS.t30 VSS.t29 nfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X50 a_439_4102# AND_3_magic_3.A.t10 VDD.t9 VDD.t5 pfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
X51 a_439_5355# AND_3_magic_5.B.t5 VDD.t85 VDD.t84 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X52 a_1185_1271# A.t6 VSS.t85 VSS.t84 nfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X53 VDD AND_3_magic_5.B.t6 a_439_6016# VDD.t86 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X54 VSS AND_3_magic_5.C.t7 a_1091_6027# VSS.t38 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X55 AND_1.A a_252_1525# VDD.t28 VDD.t27 pfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X56 VDD a_439_5355# S2.t1 VDD.t72 pfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X57 a_252_1525# C.t6 a_400_841# VDD.t30 pfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X58 a_439_4102# AND_3_magic_3.A.t11 a_587_4113# VSS.t1 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X59 a_587_6027# AND_3_magic_5.B.t7 a_1091_6027# VSS.t37 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X60 VDD AND_3_magic_3.A.t12 a_439_5355# VDD.t7 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X61 a_1091_3452# C.t7 VSS.t25 VSS.t24 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X62 AND_3_magic_5.B B.t9 VSS.t42 VSS.t41 nfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X63 a_400_841# B.t10 VDD.t96 VDD.t25 pfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
X64 a_439_6016# AND_3_magic_5.C.t8 VDD.t101 VDD.t100 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X65 a_439_6016# AND_3_magic_5.B.t8 VDD.t90 VDD.t89 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X66 AND_3_magic_5.C C.t8 VDD.t37 VDD.t36 pfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X67 VDD.t57 VDD.t56 VDD.t57 VDD.t52 pfet_03v3 ad=0 pd=0 as=89.8f ps=0.92u w=0.25u l=0.28u
X68 a_587_4113# AND_3_magic_3.A.t13 a_439_4102# VSS.t6 nfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
X69 VDD a_439_6016# S1.t1 VDD.t75 pfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X70 a_1091_6027# AND_3_magic_5.B.t9 a_587_6027# VSS.t0 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X71 a_439_5355# AND_3_magic_3.A.t14 VDD.t6 VDD.t5 pfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
X72 VSS C.t9 a_1091_3452# VSS.t68 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X73 VSS.t21 VSS.t19 VSS.t21 VSS.t20 nfet_03v3 ad=0 pd=0 as=0.155p ps=1.64u w=0.25u l=0.28u
X74 VDD AND_3_magic_3.A.t15 a_439_6016# VDD.t2 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X75 VDD AND_3_magic_5.C.t9 a_439_2188# VDD.t102 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X76 a_1091_2199# AND_3_magic_5.C.t10 VSS.t48 VSS.t47 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X77 VDD.t55 VDD.t54 VDD.t55 VDD.t27 pfet_03v3 ad=0 pd=0 as=0.155p ps=1.64u w=0.25u l=0.28u
X78 AND_3_magic_3.A A.t7 VSS.t87 VSS.t86 nfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X79 a_1091_6027# AND_3_magic_5.B.t10 a_587_6027# VSS.t26 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X80 a_252_1525# C.t10 a_400_841# VDD.t30 pfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X81 a_587_6027# AND_3_magic_3.A.t16 a_439_6016# VSS.t5 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X82 VSS C.t11 a_1091_3452# VSS.t53 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X83 a_439_6016# AND_3_magic_3.A.t17 VDD.t1 VDD.t0 pfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
X84 S1 a_439_6016# VSS.t32 VSS.t31 nfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X85 VSS AND_3_magic_5.C.t11 a_1091_2199# VSS.t49 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X86 S6 a_1333_1282# VSS.t8 VSS.t7 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X87 VDD.t53 VDD.t51 VDD.t53 VDD.t52 pfet_03v3 ad=0 pd=0 as=89.8f ps=0.92u w=0.25u l=0.28u
X88 S5 a_439_2188# VDD.t120 VDD.t113 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X89 VSS.t18 VSS.t16 VSS.t18 VSS.t17 nfet_03v3 ad=0 pd=0 as=0.155p ps=1.64u w=0.25u l=0.28u
X90 a_439_6016# AND_3_magic_3.A.t18 a_587_6027# VSS.t4 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X91 a_400_841# B.t11 VDD.t97 VDD.t25 pfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
X92 a_587_3452# B.t12 a_1091_3452# VSS.t9 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X93 a_1333_1282# AND_1.A VDD.t99 VDD.t98 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X94 VDD.t50 VDD.t49 VDD.t50 VDD.t45 pfet_03v3 ad=0 pd=0 as=89.8f ps=0.92u w=0.25u l=0.28u
X95 VDD C.t12 a_439_3441# VDD.t102 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X96 a_1091_5366# C.t13 VSS.t77 VSS.t56 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X97 VSS AND_3_magic_5.C.t12 a_1091_2199# VSS.t64 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X98 a_1091_3452# B.t13 a_587_3452# VSS.t71 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X99 VDD.t48 VDD.t47 VDD.t48 VDD.t42 pfet_03v3 ad=0 pd=0 as=89.8f ps=0.92u w=0.25u l=0.28u
X100 a_587_6027# AND_3_magic_3.A.t19 a_439_6016# VSS.t3 nfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
X101 VDD AND_3_magic_5.B.t11 a_439_2188# VDD.t66 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X102 a_587_2199# AND_3_magic_5.B.t12 a_1091_2199# VSS.t27 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X103 VSS C.t14 a_1091_5366# VSS.t58 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X104 VSS.t15 VSS.t13 VSS.t15 VSS.t14 nfet_03v3 ad=0 pd=0 as=0.155p ps=1.64u w=0.25u l=0.28u
X105 S4 a_439_3441# VDD.t114 VDD.t113 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X106 VDD AND_3_magic_5.C.t13 a_439_4102# VDD.t91 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X107 a_1091_3452# B.t14 a_587_3452# VSS.t72 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X108 AND_3_magic_5.B B.t15 VDD.t129 VDD.t128 pfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X109 AND_1.A a_252_1525# VSS.t23 VSS.t22 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
X110 a_587_3452# AND_3_magic_3.A.t20 a_439_3441# VSS.t2 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X111 a_1091_2199# AND_3_magic_5.B.t13 a_587_2199# VSS.t28 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X112 VDD.t46 VDD.t44 VDD.t46 VDD.t45 pfet_03v3 ad=0 pd=0 as=89.8f ps=0.92u w=0.25u l=0.28u
X113 S4 a_439_3441# VSS.t61 VSS.t29 nfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X114 a_439_2188# AND_3_magic_5.C.t14 VDD.t123 VDD.t80 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X115 a_252_1525# C.t15 a_400_841# VDD.t30 pfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X116 a_439_2188# AND_3_magic_5.B.t14 VDD.t69 VDD.t20 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X117 a_1091_4113# AND_3_magic_5.C.t15 VSS.t67 VSS.t24 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X118 VSS C.t16 a_1091_5366# VSS.t38 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X119 VDD a_439_2188# S5.t1 VDD.t115 pfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X120 VDD.t43 VDD.t41 VDD.t43 VDD.t42 pfet_03v3 ad=0 pd=0 as=89.8f ps=0.92u w=0.25u l=0.28u
X121 S3 a_439_4102# VDD.t71 VDD.t70 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X122 VDD B.t16 AND_3_magic_5.B VDD.t130 pfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
X123 a_439_3441# AND_3_magic_3.A.t21 a_587_3452# VSS.t1 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X124 VDD B.t17 a_439_3441# VDD.t66 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X125 a_1091_2199# AND_3_magic_5.B.t15 a_587_2199# VSS.t90 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X126 a_587_5366# AND_3_magic_5.B.t16 a_1091_5366# VSS.t37 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X127 a_587_2199# A.t8 a_439_2188# VSS.t88 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X128 VDD A.t9 a_439_2188# VDD.t15 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X129 VSS AND_3_magic_5.C.t16 a_1091_4113# VSS.t68 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X130 S5 a_439_2188# VSS.t63 VSS.t62 nfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X131 VDD C.t17 a_439_5355# VDD.t91 pfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X132 AND_3_magic_3.A A.t10 VDD.t127 VDD.t126 pfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X133 VDD.t40 VDD.t38 VDD.t40 VDD.t39 pfet_03v3 ad=0 pd=0 as=89.8f ps=0.92u w=0.25u l=0.28u
R0 AND_3_magic_3.A.n14 AND_3_magic_3.A.t20 33.6616
R1 AND_3_magic_3.A.n10 AND_3_magic_3.A.t9 33.6616
R2 AND_3_magic_3.A.n4 AND_3_magic_3.A.t4 33.6616
R3 AND_3_magic_3.A.n1 AND_3_magic_3.A.t16 33.6616
R4 AND_3_magic_3.A.n9 AND_3_magic_3.A.t7 33.5692
R5 AND_3_magic_3.A.n0 AND_3_magic_3.A.t15 33.5692
R6 AND_3_magic_3.A.n16 AND_3_magic_3.A.t3 33.4389
R7 AND_3_magic_3.A.n6 AND_3_magic_3.A.t12 33.4389
R8 AND_3_magic_3.A.n15 AND_3_magic_3.A.n14 22.7116
R9 AND_3_magic_3.A.n11 AND_3_magic_3.A.n10 22.7116
R10 AND_3_magic_3.A.n5 AND_3_magic_3.A.n4 22.7116
R11 AND_3_magic_3.A.n2 AND_3_magic_3.A.n1 22.7116
R12 AND_3_magic_3.A.n17 AND_3_magic_3.A.n15 16.8166
R13 AND_3_magic_3.A.n12 AND_3_magic_3.A.n11 16.8166
R14 AND_3_magic_3.A.n7 AND_3_magic_3.A.n5 16.8166
R15 AND_3_magic_3.A.n3 AND_3_magic_3.A.n2 16.8166
R16 AND_3_magic_3.A AND_3_magic_3.A.n18 15.6576
R17 AND_3_magic_3.A.n9 AND_3_magic_3.A.t10 11.4719
R18 AND_3_magic_3.A.n0 AND_3_magic_3.A.t17 11.4719
R19 AND_3_magic_3.A.n16 AND_3_magic_3.A.t5 11.3416
R20 AND_3_magic_3.A.n6 AND_3_magic_3.A.t14 11.3416
R21 AND_3_magic_3.A.n14 AND_3_magic_3.A.t21 10.9505
R22 AND_3_magic_3.A.n15 AND_3_magic_3.A.t2 10.9505
R23 AND_3_magic_3.A.n10 AND_3_magic_3.A.t11 10.9505
R24 AND_3_magic_3.A.n11 AND_3_magic_3.A.t13 10.9505
R25 AND_3_magic_3.A.n4 AND_3_magic_3.A.t6 10.9505
R26 AND_3_magic_3.A.n5 AND_3_magic_3.A.t8 10.9505
R27 AND_3_magic_3.A.n1 AND_3_magic_3.A.t18 10.9505
R28 AND_3_magic_3.A.n2 AND_3_magic_3.A.t19 10.9505
R29 AND_3_magic_3.A AND_3_magic_3.A.n17 6.68888
R30 AND_3_magic_3.A AND_3_magic_3.A.n12 6.68888
R31 AND_3_magic_3.A AND_3_magic_3.A.n7 6.68888
R32 AND_3_magic_3.A AND_3_magic_3.A.n3 6.68888
R33 AND_3_magic_3.A.n8 AND_3_magic_3.A 4.6195
R34 AND_3_magic_3.A.n17 AND_3_magic_3.A.n16 4.17193
R35 AND_3_magic_3.A.n7 AND_3_magic_3.A.n6 4.17193
R36 AND_3_magic_3.A.n12 AND_3_magic_3.A.n9 4.04157
R37 AND_3_magic_3.A.n3 AND_3_magic_3.A.n0 4.04157
R38 AND_3_magic_3.A.n18 AND_3_magic_3.A 2.90789
R39 AND_3_magic_3.A.n13 AND_3_magic_3.A 2.90789
R40 AND_3_magic_3.A.n8 AND_3_magic_3.A 2.90789
R41 AND_3_magic_3.A.n18 AND_3_magic_3.A.n13 1.71211
R42 AND_3_magic_3.A.n13 AND_3_magic_3.A.n8 1.29425
R43 VSS.n254 VSS.n253 8568.18
R44 VSS.n163 VSS.n162 8146.86
R45 VSS.n240 VSS.n239 4225.09
R46 VSS.n133 VSS.n132 4223.98
R47 VSS.n134 VSS.n133 3250
R48 VSS.n72 VSS.n71 1846.96
R49 VSS.n120 VSS.n119 1010.97
R50 VSS.n268 VSS.n267 688.559
R51 VSS.n255 VSS.n254 686.29
R52 VSS.n135 VSS.n134 326.76
R53 VSS.n47 VSS.t38 162.014
R54 VSS.n109 VSS.t53 162.014
R55 VSS.n271 VSS.t14 151.483
R56 VSS.n259 VSS.t20 151.483
R57 VSS.n245 VSS.t17 150.632
R58 VSS.n38 VSS.t58 142.572
R59 VSS.n100 VSS.t68 142.572
R60 VSS.n210 VSS.t64 125.677
R61 VSS.n30 VSS.t37 123.132
R62 VSS.n92 VSS.t9 123.132
R63 VSS.n175 VSS.t44 120.65
R64 VSS.n210 VSS.t84 110.597
R65 VSS.n174 VSS.t49 110.597
R66 VSS.n152 VSS.t88 106.668
R67 VSS.n20 VSS.t5 103.689
R68 VSS.n82 VSS.t2 103.689
R69 VSS.n227 VSS.t33 96.3988
R70 VSS.n263 VSS.t41 96.3988
R71 VSS.n249 VSS.t86 95.8572
R72 VSS.n164 VSS.t27 95.5148
R73 VSS.n164 VSS.n163 85.4607
R74 VSS.n17 VSS.t4 84.2478
R75 VSS.n11 VSS.t3 84.2478
R76 VSS.n79 VSS.t1 84.2478
R77 VSS.n73 VSS.t6 84.2478
R78 VSS.n26 VSS.t0 64.8061
R79 VSS.n88 VSS.t71 64.8061
R80 VSS.t35 VSS.t80 63.3338
R81 VSS.n158 VSS.t28 50.2712
R82 VSS.n35 VSS.t26 45.3644
R83 VSS.n97 VSS.t72 45.3644
R84 VSS.n181 VSS.t10 40.0005
R85 VSS.n169 VSS.t90 35.19
R86 VSS.n195 VSS.t22 33.3338
R87 VSS.n44 VSS.t56 25.9227
R88 VSS.n106 VSS.t24 25.9227
R89 VSS.n207 VSS.n206 25.1358
R90 VSS.n143 VSS.t35 23.3338
R91 VSS.n181 VSS.n180 23.3338
R92 VSS.n220 VSS.t7 22.6223
R93 VSS.n207 VSS.t47 20.1088
R94 VSS.n129 VSS.t81 20.1088
R95 VSS.n242 VSS.t16 16.6451
R96 VSS.n235 VSS.t19 16.6451
R97 VSS.n231 VSS.t13 16.6451
R98 VSS.n264 VSS.n262 10.7922
R99 VSS.n262 VSS.n260 10.7922
R100 VSS.n250 VSS.n248 10.7922
R101 VSS.n248 VSS.n246 10.7922
R102 VSS.n167 VSS.n165 10.4059
R103 VSS.n95 VSS.n93 10.2672
R104 VSS.n33 VSS.n31 10.2672
R105 VSS.n192 VSS.n190 10.0121
R106 VSS.n136 VSS.t8 9.13659
R107 VSS.n194 VSS.t23 9.04072
R108 VSS.n241 VSS.t87 6.73354
R109 VSS.n234 VSS.t42 6.73354
R110 VSS.n230 VSS.t34 6.73354
R111 VSS.n191 VSS.t52 6.66717
R112 VSS.n54 VSS.t31 6.48106
R113 VSS.n116 VSS.t29 6.48106
R114 VSS.n226 VSS.n223 5.96355
R115 VSS.n67 VSS.n66 5.6705
R116 VSS.n67 VSS.t61 5.6705
R117 VSS.n69 VSS.n68 5.6705
R118 VSS.n69 VSS.t25 5.6705
R119 VSS.n62 VSS.n61 5.6705
R120 VSS.n62 VSS.t30 5.6705
R121 VSS.n64 VSS.n63 5.6705
R122 VSS.n64 VSS.t67 5.6705
R123 VSS.n140 VSS.n139 5.6705
R124 VSS.n140 VSS.t85 5.6705
R125 VSS.n125 VSS.n124 5.6705
R126 VSS.n125 VSS.t63 5.6705
R127 VSS.n127 VSS.n126 5.6705
R128 VSS.n127 VSS.t48 5.6705
R129 VSS.n178 VSS.n177 5.6705
R130 VSS.n178 VSS.t36 5.6705
R131 VSS.n6 VSS.n5 5.6705
R132 VSS.n6 VSS.t89 5.6705
R133 VSS.n8 VSS.n7 5.6705
R134 VSS.n8 VSS.t77 5.6705
R135 VSS.n1 VSS.n0 5.6705
R136 VSS.n1 VSS.t32 5.6705
R137 VSS.n3 VSS.n2 5.6705
R138 VSS.n3 VSS.t57 5.6705
R139 VSS.n136 VSS.n135 5.30629
R140 VSS.n202 VSS.n176 5.2005
R141 VSS.n138 VSS.n137 5.2005
R142 VSS.n206 VSS.n205 5.2005
R143 VSS.n203 VSS.n175 5.2005
R144 VSS.n217 VSS.t62 5.02757
R145 VSS.n175 VSS.n174 5.02757
R146 VSS.n166 VSS.t43 5.02757
R147 VSS.n244 VSS.n240 4.42558
R148 VSS.n145 VSS.n142 4.38823
R149 VSS.n75 VSS.n72 4.37961
R150 VSS.n13 VSS.n10 4.37961
R151 VSS.n183 VSS.n179 4.36486
R152 VSS.n70 VSS.n69 3.92833
R153 VSS.n65 VSS.n64 3.92833
R154 VSS.n128 VSS.n127 3.92833
R155 VSS.n9 VSS.n8 3.92833
R156 VSS.n4 VSS.n3 3.92833
R157 VSS.n204 VSS.n140 3.46659
R158 VSS.n184 VSS.n178 3.37072
R159 VSS.n70 VSS.n67 3.27094
R160 VSS.n65 VSS.n62 3.27094
R161 VSS.n128 VSS.n125 3.27094
R162 VSS.n9 VSS.n6 3.27094
R163 VSS.n4 VSS.n1 3.27094
R164 VSS.n241 VSS.t18 2.836
R165 VSS.n234 VSS.t21 2.836
R166 VSS.n230 VSS.t15 2.836
R167 VSS.n223 VSS.n222 2.72101
R168 VSS.n123 VSS.n122 2.71312
R169 VSS.n60 VSS.n59 2.70609
R170 VSS.n200 VSS.n199 2.6005
R171 VSS.n199 VSS.n198 2.6005
R172 VSS.n197 VSS.n196 2.6005
R173 VSS.n196 VSS.n195 2.6005
R174 VSS.n193 VSS.n192 2.6005
R175 VSS.n192 VSS.n191 2.6005
R176 VSS.n190 VSS.n188 2.6005
R177 VSS.n190 VSS.n189 2.6005
R178 VSS.n187 VSS.n186 2.6005
R179 VSS.n186 VSS.n185 2.6005
R180 VSS.n182 VSS.n181 2.6005
R181 VSS.n157 VSS.n156 2.6005
R182 VSS.n156 VSS.n155 2.6005
R183 VSS.n154 VSS.n153 2.6005
R184 VSS.n153 VSS.n152 2.6005
R185 VSS.n151 VSS.n150 2.6005
R186 VSS.n150 VSS.n149 2.6005
R187 VSS.n148 VSS.n147 2.6005
R188 VSS.n147 VSS.n146 2.6005
R189 VSS.n144 VSS.n143 2.6005
R190 VSS.n56 VSS.n55 2.6005
R191 VSS.n55 VSS.n54 2.6005
R192 VSS.n52 VSS.n51 2.6005
R193 VSS.n51 VSS.n50 2.6005
R194 VSS.n49 VSS.n48 2.6005
R195 VSS.n48 VSS.n47 2.6005
R196 VSS.n46 VSS.n45 2.6005
R197 VSS.n45 VSS.n44 2.6005
R198 VSS.n43 VSS.n42 2.6005
R199 VSS.n42 VSS.n41 2.6005
R200 VSS.n40 VSS.n39 2.6005
R201 VSS.n39 VSS.n38 2.6005
R202 VSS.n37 VSS.n36 2.6005
R203 VSS.n36 VSS.n35 2.6005
R204 VSS.n34 VSS.n33 2.6005
R205 VSS.n33 VSS.n32 2.6005
R206 VSS.n31 VSS.n29 2.6005
R207 VSS.n31 VSS.n30 2.6005
R208 VSS.n28 VSS.n27 2.6005
R209 VSS.n27 VSS.n26 2.6005
R210 VSS.n25 VSS.n24 2.6005
R211 VSS.n24 VSS.n23 2.6005
R212 VSS.n22 VSS.n21 2.6005
R213 VSS.n21 VSS.n20 2.6005
R214 VSS.n19 VSS.n18 2.6005
R215 VSS.n18 VSS.n17 2.6005
R216 VSS.n16 VSS.n15 2.6005
R217 VSS.n15 VSS.n14 2.6005
R218 VSS.n12 VSS.n11 2.6005
R219 VSS.n59 VSS.n58 2.6005
R220 VSS.n58 VSS.n57 2.6005
R221 VSS.n118 VSS.n117 2.6005
R222 VSS.n117 VSS.n116 2.6005
R223 VSS.n114 VSS.n113 2.6005
R224 VSS.n113 VSS.n112 2.6005
R225 VSS.n111 VSS.n110 2.6005
R226 VSS.n110 VSS.n109 2.6005
R227 VSS.n108 VSS.n107 2.6005
R228 VSS.n107 VSS.n106 2.6005
R229 VSS.n105 VSS.n104 2.6005
R230 VSS.n104 VSS.n103 2.6005
R231 VSS.n102 VSS.n101 2.6005
R232 VSS.n101 VSS.n100 2.6005
R233 VSS.n99 VSS.n98 2.6005
R234 VSS.n98 VSS.n97 2.6005
R235 VSS.n96 VSS.n95 2.6005
R236 VSS.n95 VSS.n94 2.6005
R237 VSS.n93 VSS.n91 2.6005
R238 VSS.n93 VSS.n92 2.6005
R239 VSS.n90 VSS.n89 2.6005
R240 VSS.n89 VSS.n88 2.6005
R241 VSS.n87 VSS.n86 2.6005
R242 VSS.n86 VSS.n85 2.6005
R243 VSS.n84 VSS.n83 2.6005
R244 VSS.n83 VSS.n82 2.6005
R245 VSS.n81 VSS.n80 2.6005
R246 VSS.n80 VSS.n79 2.6005
R247 VSS.n78 VSS.n77 2.6005
R248 VSS.n77 VSS.n76 2.6005
R249 VSS.n74 VSS.n73 2.6005
R250 VSS.n122 VSS.n121 2.6005
R251 VSS.n121 VSS.n120 2.6005
R252 VSS.n219 VSS.n218 2.6005
R253 VSS.n218 VSS.n217 2.6005
R254 VSS.n215 VSS.n214 2.6005
R255 VSS.n214 VSS.n213 2.6005
R256 VSS.n212 VSS.n211 2.6005
R257 VSS.n211 VSS.n210 2.6005
R258 VSS.n209 VSS.n208 2.6005
R259 VSS.n208 VSS.n207 2.6005
R260 VSS.n131 VSS.n130 2.6005
R261 VSS.n130 VSS.n129 2.6005
R262 VSS.n173 VSS.n172 2.6005
R263 VSS.n174 VSS.n173 2.6005
R264 VSS.n171 VSS.n170 2.6005
R265 VSS.n170 VSS.n169 2.6005
R266 VSS.n168 VSS.n167 2.6005
R267 VSS.n167 VSS.n166 2.6005
R268 VSS.n165 VSS.n161 2.6005
R269 VSS.n165 VSS.n164 2.6005
R270 VSS.n160 VSS.n159 2.6005
R271 VSS.n159 VSS.n158 2.6005
R272 VSS.n222 VSS.n221 2.6005
R273 VSS.n221 VSS.n220 2.6005
R274 VSS.n252 VSS.n238 2.6005
R275 VSS.n238 VSS.n237 2.6005
R276 VSS.n251 VSS.n250 2.6005
R277 VSS.n250 VSS.n249 2.6005
R278 VSS.n248 VSS 2.6005
R279 VSS.n248 VSS.n247 2.6005
R280 VSS.n246 VSS.n245 2.6005
R281 VSS.n266 VSS.n233 2.6005
R282 VSS.n233 VSS.n232 2.6005
R283 VSS.n265 VSS.n264 2.6005
R284 VSS.n264 VSS.n263 2.6005
R285 VSS.n262 VSS 2.6005
R286 VSS.n262 VSS.n261 2.6005
R287 VSS.n260 VSS.n258 2.6005
R288 VSS.n260 VSS.n259 2.6005
R289 VSS.n257 VSS.n256 2.6005
R290 VSS.n256 VSS.n255 2.6005
R291 VSS.n226 VSS.n225 2.6005
R292 VSS.n225 VSS.n224 2.6005
R293 VSS.n229 VSS.n228 2.6005
R294 VSS.n228 VSS.n227 2.6005
R295 VSS VSS.n276 2.6005
R296 VSS.n276 VSS.n275 2.6005
R297 VSS.n273 VSS.n272 2.6005
R298 VSS.n272 VSS.n271 2.6005
R299 VSS.n270 VSS.n269 2.6005
R300 VSS.n269 VSS.n268 2.6005
R301 VSS.n123 VSS.n60 2.45364
R302 VSS.n223 VSS.n123 2.44979
R303 VSS.n246 VSS.n244 1.74196
R304 VSS.n145 VSS.n144 1.72392
R305 VSS.n13 VSS.n12 1.7162
R306 VSS.n75 VSS.n74 1.7162
R307 VSS.n183 VSS.n182 1.70135
R308 VSS.n242 VSS.n241 1.70051
R309 VSS.n235 VSS.n234 1.70051
R310 VSS.n231 VSS.n230 1.70051
R311 VSS.n60 VSS 1.09979
R312 VSS.n78 VSS.n75 0.547544
R313 VSS.n16 VSS.n13 0.547544
R314 VSS.n148 VSS.n145 0.544635
R315 VSS.n184 VSS.n183 0.53486
R316 VSS.n257 VSS.n252 0.515798
R317 VSS.n270 VSS.n266 0.505625
R318 VSS.n244 VSS.n243 0.477715
R319 VSS.n201 VSS.n200 0.450204
R320 VSS.n115 VSS.n65 0.32137
R321 VSS.n115 VSS.n70 0.32137
R322 VSS.n216 VSS.n128 0.32137
R323 VSS.n53 VSS.n4 0.32137
R324 VSS.n53 VSS.n9 0.32137
R325 VSS.n202 VSS.n201 0.248691
R326 VSS.n205 VSS.n138 0.1955
R327 VSS.n203 VSS.n202 0.193921
R328 VSS.n252 VSS.n251 0.125375
R329 VSS.n251 VSS 0.125375
R330 VSS.n266 VSS.n265 0.125375
R331 VSS.n265 VSS 0.125375
R332 VSS.n258 VSS.n257 0.125375
R333 VSS.n229 VSS.n226 0.125375
R334 VSS VSS.n229 0.125375
R335 VSS.n273 VSS.n270 0.125375
R336 VSS.n200 VSS.n197 0.0976053
R337 VSS.n188 VSS.n187 0.0976053
R338 VSS.n222 VSS.n219 0.0975588
R339 VSS.n215 VSS.n212 0.0975588
R340 VSS.n212 VSS.n209 0.0975588
R341 VSS.n209 VSS.n131 0.0975588
R342 VSS.n172 VSS.n131 0.0975588
R343 VSS.n172 VSS.n171 0.0975588
R344 VSS.n171 VSS.n168 0.0975588
R345 VSS.n161 VSS.n160 0.0975588
R346 VSS.n160 VSS.n157 0.0975588
R347 VSS.n157 VSS.n154 0.0975588
R348 VSS.n154 VSS.n151 0.0975588
R349 VSS.n151 VSS.n148 0.0975588
R350 VSS.n122 VSS.n118 0.0966165
R351 VSS.n114 VSS.n111 0.0966165
R352 VSS.n111 VSS.n108 0.0966165
R353 VSS.n108 VSS.n105 0.0966165
R354 VSS.n105 VSS.n102 0.0966165
R355 VSS.n102 VSS.n99 0.0966165
R356 VSS.n99 VSS.n96 0.0966165
R357 VSS.n91 VSS.n90 0.0966165
R358 VSS.n90 VSS.n87 0.0966165
R359 VSS.n87 VSS.n84 0.0966165
R360 VSS.n84 VSS.n81 0.0966165
R361 VSS.n81 VSS.n78 0.0966165
R362 VSS.n59 VSS.n56 0.0966165
R363 VSS.n52 VSS.n49 0.0966165
R364 VSS.n49 VSS.n46 0.0966165
R365 VSS.n46 VSS.n43 0.0966165
R366 VSS.n43 VSS.n40 0.0966165
R367 VSS.n40 VSS.n37 0.0966165
R368 VSS.n37 VSS.n34 0.0966165
R369 VSS.n29 VSS.n28 0.0966165
R370 VSS.n28 VSS.n25 0.0966165
R371 VSS.n25 VSS.n22 0.0966165
R372 VSS.n22 VSS.n19 0.0966165
R373 VSS.n19 VSS.n16 0.0966165
R374 VSS.n193 VSS 0.0960263
R375 VSS.n91 VSS 0.0957427
R376 VSS.n29 VSS 0.0957427
R377 VSS VSS.n203 0.0944474
R378 VSS.n243 VSS.n242 0.0905
R379 VSS.n236 VSS.n235 0.0905
R380 VSS.n274 VSS.n231 0.0905
R381 VSS.n243 VSS 0.08825
R382 VSS.n236 VSS 0.08825
R383 VSS VSS.n274 0.08825
R384 VSS.n219 VSS.n216 0.0763824
R385 VSS.n118 VSS.n115 0.0756456
R386 VSS.n56 VSS.n53 0.0756456
R387 VSS.n197 VSS.n194 0.0747105
R388 VSS.n138 VSS.n136 0.0715526
R389 VSS.n204 VSS 0.0676053
R390 VSS.n161 VSS.n141 0.0499118
R391 VSS.n141 VSS 0.0472647
R392 VSS.n258 VSS.n236 0.037625
R393 VSS.n274 VSS.n273 0.037625
R394 VSS.n194 VSS.n193 0.0233947
R395 VSS.n205 VSS.n204 0.0226053
R396 VSS.n187 VSS.n184 0.0218158
R397 VSS.n216 VSS.n215 0.0216765
R398 VSS.n115 VSS.n114 0.0214709
R399 VSS.n53 VSS.n52 0.0214709
R400 VSS.n188 VSS 0.00207895
R401 VSS.n168 VSS 0.00138235
R402 VSS.n96 VSS 0.00137379
R403 VSS.n34 VSS 0.00137379
R404 VDD.t98 VDD.n220 284.437
R405 VDD.n245 VDD.t98 170.881
R406 VDD.n249 VDD.t18 147.625
R407 VDD.n53 VDD.t78 96.0457
R408 VDD.n43 VDD.t109 84.7463
R409 VDD.n258 VDD.t106 75.2467
R410 VDD.n274 VDD.t31 73.5038
R411 VDD.n253 VDD.t130 73.5038
R412 VDD.n33 VDD.t59 73.4468
R413 VDD.n231 VDD.t30 64.9948
R414 VDD.n24 VDD.t89 62.1474
R415 VDD.n127 VDD.t70 55.9829
R416 VDD.n201 VDD.t113 55.9829
R417 VDD.n14 VDD.t0 53.828
R418 VDD.n117 VDD.t91 49.3968
R419 VDD.n191 VDD.t102 49.3968
R420 VDD.n261 VDD.t126 47.8628
R421 VDD.n214 VDD.t36 47.8628
R422 VDD.n269 VDD.t128 47.8628
R423 VDD.n20 VDD.t2 47.0815
R424 VDD.n107 VDD.t39 42.8106
R425 VDD.n181 VDD.t45 42.8106
R426 VDD.n98 VDD.t84 36.2244
R427 VDD.n172 VDD.t20 36.2244
R428 VDD.n30 VDD.t86 35.782
R429 VDD.n88 VDD.t5 32.5123
R430 VDD.n162 VDD.t13 32.5123
R431 VDD.n94 VDD.t7 27.4429
R432 VDD.n168 VDD.t15 27.4429
R433 VDD.n40 VDD.t100 24.4826
R434 VDD.n104 VDD.t22 20.8567
R435 VDD.n178 VDD.t66 20.8567
R436 VDD.n10 VDD.t58 18.4701
R437 VDD.n6 VDD.t63 18.4701
R438 VDD.n74 VDD.t47 18.4701
R439 VDD.n70 VDD.t41 18.4701
R440 VDD.n82 VDD.t38 18.4701
R441 VDD.n78 VDD.t61 18.4701
R442 VDD.n148 VDD.t56 18.4701
R443 VDD.n144 VDD.t51 18.4701
R444 VDD.n156 VDD.t49 18.4701
R445 VDD.n152 VDD.t44 18.4701
R446 VDD.n223 VDD.t54 17.4273
R447 VDD.n228 VDD.t25 16.5878
R448 VDD.n241 VDD.t27 14.3073
R449 VDD.n114 VDD.t34 14.2705
R450 VDD.n188 VDD.t80 14.2705
R451 VDD.n50 VDD.t64 13.1832
R452 VDD.n270 VDD.n268 9.713
R453 VDD.n268 VDD.n254 9.713
R454 VDD.n262 VDD.n260 9.713
R455 VDD.n13 VDD.t1 9.36138
R456 VDD.n62 VDD.n2 9.36138
R457 VDD.n136 VDD.n66 9.36138
R458 VDD.n136 VDD.n65 9.36138
R459 VDD.n87 VDD.t9 9.36138
R460 VDD.n87 VDD.t6 9.36138
R461 VDD.n210 VDD.n140 9.36138
R462 VDD.n210 VDD.n139 9.36138
R463 VDD.n161 VDD.t105 9.36138
R464 VDD.n161 VDD.t14 9.36138
R465 VDD.n221 VDD.t29 9.12573
R466 VDD.n224 VDD.t96 9.12573
R467 VDD.n238 VDD.n236 9.01096
R468 VDD.n221 VDD.t28 8.9005
R469 VDD.n226 VDD.t142 8.9005
R470 VDD.n225 VDD.t26 8.9005
R471 VDD.n224 VDD.t97 8.9005
R472 VDD.n41 VDD.n39 8.88511
R473 VDD.n115 VDD.n113 8.77265
R474 VDD.n189 VDD.n187 8.77265
R475 VDD.n124 VDD.t42 7.68436
R476 VDD.n198 VDD.t52 7.68436
R477 VDD.n246 VDD.t99 6.74137
R478 VDD.n213 VDD.n212 6.49074
R479 VDD.n12 VDD.n11 6.3005
R480 VDD.n12 VDD.t90 6.3005
R481 VDD.n9 VDD.n8 6.3005
R482 VDD.n9 VDD.t60 6.3005
R483 VDD.n7 VDD.t101 6.3005
R484 VDD.n5 VDD.n4 6.3005
R485 VDD.n5 VDD.t65 6.3005
R486 VDD.n3 VDD.t79 6.3005
R487 VDD.n73 VDD.n72 6.3005
R488 VDD.n71 VDD.t48 6.3005
R489 VDD.n71 VDD.t71 6.3005
R490 VDD.n69 VDD.n68 6.3005
R491 VDD.n67 VDD.t43 6.3005
R492 VDD.n67 VDD.t140 6.3005
R493 VDD.n81 VDD.n80 6.3005
R494 VDD.n79 VDD.t40 6.3005
R495 VDD.n79 VDD.t112 6.3005
R496 VDD.n77 VDD.n76 6.3005
R497 VDD.n75 VDD.t62 6.3005
R498 VDD.n75 VDD.t35 6.3005
R499 VDD.n86 VDD.n85 6.3005
R500 VDD.n86 VDD.t141 6.3005
R501 VDD.n84 VDD.n83 6.3005
R502 VDD.n84 VDD.t85 6.3005
R503 VDD.n147 VDD.n146 6.3005
R504 VDD.n147 VDD.t57 6.3005
R505 VDD.n145 VDD.t120 6.3005
R506 VDD.n143 VDD.n142 6.3005
R507 VDD.n141 VDD.t53 6.3005
R508 VDD.n141 VDD.t114 6.3005
R509 VDD.n155 VDD.n154 6.3005
R510 VDD.n153 VDD.t50 6.3005
R511 VDD.n153 VDD.t123 6.3005
R512 VDD.n151 VDD.n150 6.3005
R513 VDD.n149 VDD.t46 6.3005
R514 VDD.n149 VDD.t81 6.3005
R515 VDD.n160 VDD.n159 6.3005
R516 VDD.n160 VDD.t69 6.3005
R517 VDD.n158 VDD.n157 6.3005
R518 VDD.n158 VDD.t21 6.3005
R519 VDD.n256 VDD.n255 6.3005
R520 VDD.n256 VDD.t127 6.3005
R521 VDD.n251 VDD.n250 6.3005
R522 VDD.n251 VDD.t129 6.3005
R523 VDD.n247 VDD.n220 6.3005
R524 VDD.n1 VDD.n0 6.3005
R525 VDD.n1 VDD.t37 6.3005
R526 VDD.n59 VDD.t75 4.86375
R527 VDD.n222 VDD.t55 4.451
R528 VDD.n207 VDD.t115 3.97221
R529 VDD.n133 VDD.t72 3.97219
R530 VDD.n219 VDD.t19 3.6405
R531 VDD.n219 VDD.n218 3.6405
R532 VDD.n61 VDD.n60 3.1505
R533 VDD.n58 VDD.n57 3.1505
R534 VDD.n57 VDD.n56 3.1505
R535 VDD.n55 VDD.n54 3.1505
R536 VDD.n54 VDD.n53 3.1505
R537 VDD.n52 VDD.n51 3.1505
R538 VDD.n51 VDD.n50 3.1505
R539 VDD.n48 VDD.n47 3.1505
R540 VDD.n47 VDD.n46 3.1505
R541 VDD.n45 VDD.n44 3.1505
R542 VDD.n44 VDD.n43 3.1505
R543 VDD.n42 VDD.n41 3.1505
R544 VDD.n41 VDD.n40 3.1505
R545 VDD.n39 VDD.n37 3.1505
R546 VDD.n39 VDD.n38 3.1505
R547 VDD.n35 VDD.n34 3.1505
R548 VDD.n34 VDD.n33 3.1505
R549 VDD.n32 VDD.n31 3.1505
R550 VDD.n31 VDD.n30 3.1505
R551 VDD.n29 VDD.n28 3.1505
R552 VDD.n28 VDD.n27 3.1505
R553 VDD.n26 VDD.n25 3.1505
R554 VDD.n25 VDD.n24 3.1505
R555 VDD.n22 VDD.n21 3.1505
R556 VDD.n21 VDD.n20 3.1505
R557 VDD.n19 VDD.n18 3.1505
R558 VDD.n18 VDD.n17 3.1505
R559 VDD.n16 VDD.n15 3.1505
R560 VDD.n135 VDD.n134 3.1505
R561 VDD.n132 VDD.n131 3.1505
R562 VDD.n131 VDD.n130 3.1505
R563 VDD.n129 VDD.n128 3.1505
R564 VDD.n128 VDD.n127 3.1505
R565 VDD.n126 VDD.n125 3.1505
R566 VDD.n125 VDD.n124 3.1505
R567 VDD.n122 VDD.n121 3.1505
R568 VDD.n121 VDD.n120 3.1505
R569 VDD.n119 VDD.n118 3.1505
R570 VDD.n118 VDD.n117 3.1505
R571 VDD.n116 VDD.n115 3.1505
R572 VDD.n115 VDD.n114 3.1505
R573 VDD.n113 VDD.n111 3.1505
R574 VDD.n113 VDD.n112 3.1505
R575 VDD.n109 VDD.n108 3.1505
R576 VDD.n108 VDD.n107 3.1505
R577 VDD.n106 VDD.n105 3.1505
R578 VDD.n105 VDD.n104 3.1505
R579 VDD.n103 VDD.n102 3.1505
R580 VDD.n102 VDD.n101 3.1505
R581 VDD.n100 VDD.n99 3.1505
R582 VDD.n99 VDD.n98 3.1505
R583 VDD.n96 VDD.n95 3.1505
R584 VDD.n95 VDD.n94 3.1505
R585 VDD.n93 VDD.n92 3.1505
R586 VDD.n92 VDD.n91 3.1505
R587 VDD.n90 VDD.n89 3.1505
R588 VDD.n209 VDD.n208 3.1505
R589 VDD.n206 VDD.n205 3.1505
R590 VDD.n205 VDD.n204 3.1505
R591 VDD.n203 VDD.n202 3.1505
R592 VDD.n202 VDD.n201 3.1505
R593 VDD.n200 VDD.n199 3.1505
R594 VDD.n199 VDD.n198 3.1505
R595 VDD.n196 VDD.n195 3.1505
R596 VDD.n195 VDD.n194 3.1505
R597 VDD.n193 VDD.n192 3.1505
R598 VDD.n192 VDD.n191 3.1505
R599 VDD.n190 VDD.n189 3.1505
R600 VDD.n189 VDD.n188 3.1505
R601 VDD.n187 VDD.n185 3.1505
R602 VDD.n187 VDD.n186 3.1505
R603 VDD.n183 VDD.n182 3.1505
R604 VDD.n182 VDD.n181 3.1505
R605 VDD.n180 VDD.n179 3.1505
R606 VDD.n179 VDD.n178 3.1505
R607 VDD.n177 VDD.n176 3.1505
R608 VDD.n176 VDD.n175 3.1505
R609 VDD.n174 VDD.n173 3.1505
R610 VDD.n173 VDD.n172 3.1505
R611 VDD.n170 VDD.n169 3.1505
R612 VDD.n169 VDD.n168 3.1505
R613 VDD.n167 VDD.n166 3.1505
R614 VDD.n166 VDD.n165 3.1505
R615 VDD.n164 VDD.n163 3.1505
R616 VDD.n263 VDD.n262 3.1505
R617 VDD.n260 VDD.n259 3.1505
R618 VDD.n271 VDD.n270 3.1505
R619 VDD.n268 VDD 3.1505
R620 VDD.n268 VDD.n267 3.1505
R621 VDD.n266 VDD.n254 3.1505
R622 VDD.n243 VDD.n242 3.1505
R623 VDD.n239 VDD.n238 3.1505
R624 VDD.n238 VDD.n237 3.1505
R625 VDD.n236 VDD.n234 3.1505
R626 VDD.n236 VDD.n235 3.1505
R627 VDD.n233 VDD.n232 3.1505
R628 VDD.n232 VDD.n231 3.1505
R629 VDD.n230 VDD.n229 3.1505
R630 VDD.n216 VDD.n215 3.1505
R631 VDD VDD.n279 3.1505
R632 VDD.n279 VDD.n278 3.1505
R633 VDD.n276 VDD.n275 3.1505
R634 VDD.n248 VDD.n219 3.10137
R635 VDD.n23 VDD.n12 3.06138
R636 VDD.n97 VDD.n86 3.06138
R637 VDD.n97 VDD.n84 3.06138
R638 VDD.n171 VDD.n160 3.06138
R639 VDD.n171 VDD.n158 3.06138
R640 VDD.n257 VDD.n256 2.99094
R641 VDD.n252 VDD.n251 2.99094
R642 VDD.n217 VDD.n1 2.99094
R643 VDD.n212 VDD.n211 2.96507
R644 VDD.n138 VDD.n137 2.93063
R645 VDD.n64 VDD.n63 2.9206
R646 VDD.n10 VDD.n9 2.86655
R647 VDD.n10 VDD.n7 2.86655
R648 VDD.n6 VDD.n5 2.86655
R649 VDD.n6 VDD.n3 2.86655
R650 VDD.n74 VDD.n73 2.86655
R651 VDD.n74 VDD.n71 2.86655
R652 VDD.n70 VDD.n69 2.86655
R653 VDD.n70 VDD.n67 2.86655
R654 VDD.n82 VDD.n81 2.86655
R655 VDD.n82 VDD.n79 2.86655
R656 VDD.n78 VDD.n77 2.86655
R657 VDD.n78 VDD.n75 2.86655
R658 VDD.n148 VDD.n147 2.86655
R659 VDD.n148 VDD.n145 2.86655
R660 VDD.n144 VDD.n143 2.86655
R661 VDD.n144 VDD.n141 2.86655
R662 VDD.n156 VDD.n155 2.86655
R663 VDD.n156 VDD.n153 2.86655
R664 VDD.n152 VDD.n151 2.86655
R665 VDD.n152 VDD.n149 2.86655
R666 VDD.n138 VDD.n64 2.46136
R667 VDD.n212 VDD.n138 2.45107
R668 VDD.n260 VDD.n258 1.97857
R669 VDD.n220 VDD.t135 1.78941
R670 VDD.n222 VDD.n221 0.60793
R671 VDD.n245 VDD.n244 0.571942
R672 VDD.n258 VDD 0.53368
R673 VDD.n265 VDD.n264 0.5075
R674 VDD.n273 VDD.n272 0.505625
R675 VDD.n277 VDD.n249 0.451829
R676 VDD.n227 VDD.n226 0.367463
R677 VDD.n225 VDD.n224 0.2316
R678 VDD.n226 VDD.n225 0.22573
R679 VDD.n89 VDD.n88 0.204689
R680 VDD.n208 VDD.n207 0.204689
R681 VDD.n134 VDD.n133 0.20445
R682 VDD.n163 VDD.n162 0.20445
R683 VDD.n242 VDD.n241 0.183695
R684 VDD.n229 VDD.n228 0.183455
R685 VDD.n36 VDD.n10 0.172674
R686 VDD.n49 VDD.n6 0.172674
R687 VDD.n123 VDD.n70 0.172674
R688 VDD.n123 VDD.n74 0.172674
R689 VDD.n110 VDD.n78 0.172674
R690 VDD.n110 VDD.n82 0.172674
R691 VDD.n197 VDD.n144 0.172674
R692 VDD.n197 VDD.n148 0.172674
R693 VDD.n184 VDD.n152 0.172674
R694 VDD.n184 VDD.n156 0.172674
R695 VDD VDD.n246 0.15489
R696 VDD.n60 VDD.n59 0.127116
R697 VDD.n15 VDD.n14 0.126872
R698 VDD.n223 VDD.n222 0.125892
R699 VDD.n264 VDD.n263 0.125375
R700 VDD.n272 VDD.n271 0.125375
R701 VDD VDD.n266 0.125375
R702 VDD.n266 VDD.n265 0.125375
R703 VDD.n216 VDD.n213 0.125375
R704 VDD.n276 VDD.n273 0.125375
R705 VDD.n262 VDD.n261 0.122078
R706 VDD.n254 VDD.n253 0.122078
R707 VDD.n275 VDD.n274 0.122078
R708 VDD.n270 VDD.n269 0.121835
R709 VDD.n215 VDD.n214 0.121835
R710 VDD.n263 VDD.n257 0.118625
R711 VDD.n271 VDD.n252 0.118625
R712 VDD.n217 VDD.n216 0.118625
R713 VDD.n249 VDD.n248 0.116841
R714 VDD.n244 VDD.n243 0.0976053
R715 VDD.n234 VDD.n233 0.0976053
R716 VDD.n233 VDD.n230 0.0976053
R717 VDD.n61 VDD.n58 0.0975588
R718 VDD.n58 VDD.n55 0.0975588
R719 VDD.n55 VDD.n52 0.0975588
R720 VDD.n48 VDD.n45 0.0975588
R721 VDD.n45 VDD.n42 0.0975588
R722 VDD.n35 VDD.n32 0.0975588
R723 VDD.n32 VDD.n29 0.0975588
R724 VDD.n29 VDD.n26 0.0975588
R725 VDD.n22 VDD.n19 0.0975588
R726 VDD.n19 VDD.n16 0.0975588
R727 VDD.n135 VDD.n132 0.0966165
R728 VDD.n132 VDD.n129 0.0966165
R729 VDD.n129 VDD.n126 0.0966165
R730 VDD.n122 VDD.n119 0.0966165
R731 VDD.n119 VDD.n116 0.0966165
R732 VDD.n109 VDD.n106 0.0966165
R733 VDD.n106 VDD.n103 0.0966165
R734 VDD.n103 VDD.n100 0.0966165
R735 VDD.n96 VDD.n93 0.0966165
R736 VDD.n93 VDD.n90 0.0966165
R737 VDD.n209 VDD.n206 0.0966165
R738 VDD.n206 VDD.n203 0.0966165
R739 VDD.n203 VDD.n200 0.0966165
R740 VDD.n196 VDD.n193 0.0966165
R741 VDD.n193 VDD.n190 0.0966165
R742 VDD.n183 VDD.n180 0.0966165
R743 VDD.n180 VDD.n177 0.0966165
R744 VDD.n177 VDD.n174 0.0966165
R745 VDD.n170 VDD.n167 0.0966165
R746 VDD.n167 VDD.n164 0.0966165
R747 VDD.n239 VDD 0.0960263
R748 VDD.n42 VDD 0.0957941
R749 VDD.n116 VDD 0.0948689
R750 VDD.n190 VDD 0.0948689
R751 VDD.n240 VDD.n223 0.0924565
R752 VDD.n49 VDD.n48 0.0913824
R753 VDD.n123 VDD.n122 0.0905
R754 VDD.n197 VDD.n196 0.0905
R755 VDD.n240 VDD.n239 0.0897105
R756 VDD.n62 VDD.n61 0.0737353
R757 VDD.n136 VDD.n135 0.0730243
R758 VDD.n210 VDD.n209 0.0730243
R759 VDD.n277 VDD.n276 0.069125
R760 VDD.n37 VDD.n36 0.0631471
R761 VDD.n111 VDD.n110 0.0625388
R762 VDD.n185 VDD.n184 0.0625388
R763 VDD.n248 VDD.n247 0.0597683
R764 VDD.n64 VDD 0.0596429
R765 VDD.n230 VDD.n227 0.0573421
R766 VDD VDD.n277 0.05675
R767 VDD.n23 VDD.n22 0.0525588
R768 VDD.n97 VDD.n96 0.0520534
R769 VDD.n171 VDD.n170 0.0520534
R770 VDD.n16 VDD.n13 0.0507941
R771 VDD.n90 VDD.n87 0.0503058
R772 VDD.n164 VDD.n161 0.0503058
R773 VDD.n26 VDD.n23 0.0455
R774 VDD.n100 VDD.n97 0.0450631
R775 VDD.n174 VDD.n171 0.0450631
R776 VDD.n36 VDD.n35 0.0349118
R777 VDD.n110 VDD.n109 0.0345777
R778 VDD.n184 VDD.n183 0.0345777
R779 VDD.n63 VDD.n62 0.0243235
R780 VDD.n137 VDD.n136 0.0240922
R781 VDD.n211 VDD.n210 0.0240922
R782 VDD.n247 VDD 0.0209878
R783 VDD.n246 VDD.n245 0.00928049
R784 VDD.n243 VDD.n240 0.00839474
R785 VDD VDD.n257 0.00725
R786 VDD VDD.n252 0.00725
R787 VDD VDD.n217 0.00725
R788 VDD.n52 VDD.n49 0.00667647
R789 VDD.n126 VDD.n123 0.0066165
R790 VDD.n200 VDD.n197 0.0066165
R791 VDD.n37 VDD 0.00226471
R792 VDD.n111 VDD 0.00224757
R793 VDD.n185 VDD 0.00224757
R794 VDD.n234 VDD 0.00207895
R795 AND_3_magic_5.B AND_3_magic_5.B.t14 89.0293
R796 AND_3_magic_5.B AND_3_magic_5.B.t5 89.0293
R797 AND_3_magic_5.B AND_3_magic_5.B.t8 89.0293
R798 AND_3_magic_5.B.n7 AND_3_magic_5.B.t15 35.4088
R799 AND_3_magic_5.B.n3 AND_3_magic_5.B.t3 35.4088
R800 AND_3_magic_5.B.n0 AND_3_magic_5.B.t10 35.4088
R801 AND_3_magic_5.B.t14 AND_3_magic_5.B.n9 34.0527
R802 AND_3_magic_5.B.t5 AND_3_magic_5.B.n5 34.0527
R803 AND_3_magic_5.B.t8 AND_3_magic_5.B.n2 34.0527
R804 AND_3_magic_5.B.n8 AND_3_magic_5.B.n7 25.7624
R805 AND_3_magic_5.B.n4 AND_3_magic_5.B.n3 25.7624
R806 AND_3_magic_5.B.n1 AND_3_magic_5.B.n0 25.7624
R807 AND_3_magic_5.B.n9 AND_3_magic_5.B.n8 22.2916
R808 AND_3_magic_5.B.n5 AND_3_magic_5.B.n4 22.2916
R809 AND_3_magic_5.B.n2 AND_3_magic_5.B.n1 22.2916
R810 AND_3_magic_5.B AND_3_magic_5.B.n10 17.0101
R811 AND_3_magic_5.B.n9 AND_3_magic_5.B.t11 11.3416
R812 AND_3_magic_5.B.n5 AND_3_magic_5.B.t4 11.3416
R813 AND_3_magic_5.B.n2 AND_3_magic_5.B.t6 11.3416
R814 AND_3_magic_5.B.n8 AND_3_magic_5.B.t13 9.64693
R815 AND_3_magic_5.B.n4 AND_3_magic_5.B.t2 9.64693
R816 AND_3_magic_5.B.n1 AND_3_magic_5.B.t9 9.64693
R817 AND_3_magic_5.B.n6 AND_3_magic_5.B 5.99158
R818 AND_3_magic_5.B.n10 AND_3_magic_5.B.n6 3.50889
R819 AND_3_magic_5.B.n10 AND_3_magic_5.B 3.41854
R820 AND_3_magic_5.B.n6 AND_3_magic_5.B 3.41854
R821 AND_3_magic_5.B.n7 AND_3_magic_5.B.t12 3.25943
R822 AND_3_magic_5.B.n3 AND_3_magic_5.B.t16 3.25943
R823 AND_3_magic_5.B.n0 AND_3_magic_5.B.t7 3.25943
R824 A A.t3 75.0339
R825 A.t3 A.n6 40.4981
R826 A.n2 A.t8 33.6616
R827 A.n1 A.t9 33.5692
R828 A.t2 A.n0 31.2628
R829 A.n6 A.t6 30.7213
R830 A.n0 A.t7 27.5059
R831 A.n3 A.n2 22.7116
R832 A A.t2 18.8858
R833 A.n4 A.n3 16.8166
R834 A.n6 A.t5 13.688
R835 A.n1 A.t1 11.4719
R836 A.n2 A.t0 10.9505
R837 A.n3 A.t4 10.9505
R838 A.n0 A.t10 10.2987
R839 A.n7 A 9.28055
R840 A.n5 A 6.85336
R841 A A.n4 6.68888
R842 A.n4 A.n1 4.04157
R843 A A.n7 3.12814
R844 A.n7 A.n5 3.08139
R845 A.n5 A 2.66333
R846 C.t17 C.t5 45.3938
R847 C.t12 C.t0 45.3938
R848 C.t14 C.t17 43.2791
R849 C.t9 C.t12 43.2791
R850 C.n1 C.t16 35.6691
R851 C.n4 C.t11 35.6691
R852 C.t4 C.n0 31.2628
R853 C.n0 C.t1 27.5059
R854 C.n2 C.n1 25.6316
R855 C.n5 C.n4 25.6316
R856 C.n7 C.t2 23.8759
R857 C C.n2 21.1146
R858 C C.n5 21.1146
R859 C C.t4 18.8772
R860 C.t10 C.t15 17.338
R861 C.t15 C.t3 16.9469
R862 C.t6 C.t10 16.9469
R863 C C.n8 12.7448
R864 C.n7 C.t6 11.8831
R865 C.n0 C.t8 10.2987
R866 C.n2 C.t14 10.038
R867 C.n5 C.t9 10.038
R868 C C.n7 4.77137
R869 C.n3 C 3.67093
R870 C.n6 C 3.67093
R871 C.n8 C.n6 3.65675
R872 C.n8 C 3.36767
R873 C.n1 C.t13 3.25943
R874 C.n4 C.t7 3.25943
R875 C.n6 C.n3 3.04121
R876 C.n3 C 1.81336
R877 B B.t5 89.0293
R878 B B.t0 89.0293
R879 B.t10 B.t4 39.3684
R880 B B.t7 36.6468
R881 B.n1 B.t8 35.4088
R882 B.n5 B.t14 35.4088
R883 B.t5 B.n3 34.0527
R884 B.t0 B.n7 34.0527
R885 B.t16 B.n0 31.2628
R886 B.n0 B.t9 27.5059
R887 B.n2 B.n1 25.7624
R888 B.n6 B.n5 25.7624
R889 B.n3 B.n2 22.2916
R890 B.n7 B.n6 22.2916
R891 B.n10 B.t16 18.8525
R892 B.t2 B.t11 17.338
R893 B.t11 B.t10 16.9469
R894 B.t7 B.t2 16.9469
R895 B.n3 B.t1 11.3416
R896 B.n7 B.t17 11.3416
R897 B.n0 B.t15 10.2987
R898 B.n10 B.n9 9.8838
R899 B.n2 B.t6 9.64693
R900 B.n6 B.t13 9.64693
R901 B.n9 B.n8 3.52496
R902 B.n4 B 3.34496
R903 B.n1 B.t3 3.25943
R904 B.n5 B.t12 3.25943
R905 B.n4 B 3.17007
R906 B.n8 B 3.17007
R907 B.n9 B 2.86485
R908 B.n8 B.n4 2.57354
R909 B B.n10 0.00165385
R910 AND_3_magic_5.C.t9 AND_3_magic_5.C.t14 45.3938
R911 AND_3_magic_5.C.t13 AND_3_magic_5.C.t4 45.3938
R912 AND_3_magic_5.C.t3 AND_3_magic_5.C.t8 45.3938
R913 AND_3_magic_5.C.t11 AND_3_magic_5.C.t9 43.2791
R914 AND_3_magic_5.C.t16 AND_3_magic_5.C.t13 43.2791
R915 AND_3_magic_5.C.t6 AND_3_magic_5.C.t3 43.2791
R916 AND_3_magic_5.C.n5 AND_3_magic_5.C.t12 35.6691
R917 AND_3_magic_5.C.n2 AND_3_magic_5.C.t2 35.6691
R918 AND_3_magic_5.C.n0 AND_3_magic_5.C.t7 35.6691
R919 AND_3_magic_5.C.n6 AND_3_magic_5.C.n5 25.6316
R920 AND_3_magic_5.C.n3 AND_3_magic_5.C.n2 25.6316
R921 AND_3_magic_5.C.n1 AND_3_magic_5.C.n0 25.6316
R922 AND_3_magic_5.C AND_3_magic_5.C.n6 21.1146
R923 AND_3_magic_5.C AND_3_magic_5.C.n3 21.1146
R924 AND_3_magic_5.C AND_3_magic_5.C.n1 21.1146
R925 AND_3_magic_5.C AND_3_magic_5.C.n7 18.1627
R926 AND_3_magic_5.C.n6 AND_3_magic_5.C.t11 10.038
R927 AND_3_magic_5.C.n3 AND_3_magic_5.C.t16 10.038
R928 AND_3_magic_5.C.n1 AND_3_magic_5.C.t6 10.038
R929 AND_3_magic_5.C.n4 AND_3_magic_5.C 6.95691
R930 AND_3_magic_5.C.n7 AND_3_magic_5.C 3.91941
R931 AND_3_magic_5.C.n4 AND_3_magic_5.C 3.91941
R932 AND_3_magic_5.C.n5 AND_3_magic_5.C.t10 3.25943
R933 AND_3_magic_5.C.n2 AND_3_magic_5.C.t15 3.25943
R934 AND_3_magic_5.C.n0 AND_3_magic_5.C.t5 3.25943
R935 AND_3_magic_5.C.n7 AND_3_magic_5.C.n4 3.04121
R936 S4.n3 S4.n0 8.96638
R937 S4.n2 S4.n1 6.3005
R938 S4.n2 S4.t2 6.3005
R939 S4.n3 S4.n2 3.22377
R940 S4 S4.n3 0.0768043
R941 S2.n3 S2.n0 8.96638
R942 S2.n2 S2.n1 6.3005
R943 S2.n2 S2.t1 6.3005
R944 S2.n3 S2.n2 3.22377
R945 S2 S2.n3 0.0768043
R946 S3.n3 S3.n2 8.96638
R947 S3.n1 S3.n0 6.3005
R948 S3.n1 S3.t2 6.3005
R949 S3.n3 S3.n1 3.22377
R950 S3 S3.n3 0.0768043
R951 S1.n3 S1.n2 8.96638
R952 S1.n1 S1.n0 6.3005
R953 S1.n1 S1.t1 6.3005
R954 S1.n3 S1.n1 3.22377
R955 S1 S1.n3 0.0768043
R956 S6.n2 S6.n0 9.37773
R957 S6.n2 S6.n1 7.06778
R958 S6 S6.n2 0.0502872
R959 S5.n3 S5.n2 8.96638
R960 S5.n1 S5.n0 6.3005
R961 S5.n1 S5.t1 6.3005
R962 S5.n3 S5.n1 3.22377
R963 S5 S5.n3 0.0768043
C0 AND_3_magic_5.C A 0.177f
C1 VDD a_1333_1282# 0.411f
C2 AND_3_magic_5.B a_439_4102# 5.39e-19
C3 AND_3_magic_5.C a_439_4102# 0.111f
C4 a_439_2188# S5 0.0806f
C5 VDD a_1185_1271# 0.0146f
C6 a_587_3452# A 0.00272f
C7 AND_1.A S6 2.31e-19
C8 AND_3_magic_3.A a_587_4113# 0.0359f
C9 a_587_6027# A 0.00272f
C10 AND_3_magic_5.B a_587_2199# 0.0545f
C11 C S6 1.84e-19
C12 AND_3_magic_5.C a_587_2199# 0.457f
C13 VDD a_252_1525# 0.606f
C14 AND_1.A a_1333_1282# 0.154f
C15 A a_439_2188# 0.199f
C16 C a_1333_1282# 0.00309f
C17 AND_3_magic_3.A a_439_5355# 0.193f
C18 VDD a_1091_2199# 0.00358f
C19 AND_1.A a_1185_1271# 0.134f
C20 B a_1185_1271# 2.28e-20
C21 a_439_5355# S3 1.18e-19
C22 S5 S6 0.00586f
C23 C a_1185_1271# 1.76e-19
C24 a_252_1525# AND_1.A 0.121f
C25 S5 a_1333_1282# 1.73e-19
C26 a_439_2188# a_587_2199# 0.475f
C27 B a_252_1525# 0.022f
C28 C a_252_1525# 0.399f
C29 A S6 0.00142f
C30 AND_3_magic_3.A a_439_6016# 0.193f
C31 a_1091_2199# AND_1.A 3.04e-19
C32 S2 S3 0.00185f
C33 A a_1333_1282# 0.0865f
C34 C a_1091_2199# 7.07e-20
C35 AND_3_magic_3.A VDD 1.59f
C36 VDD S3 0.247f
C37 A a_1185_1271# 0.0448f
C38 S5 a_1091_2199# 0.0134f
C39 a_252_1525# a_400_841# 0.18f
C40 A a_252_1525# 0.0154f
C41 AND_3_magic_3.A AND_1.A 5.81e-20
C42 AND_3_magic_3.A B 3.25f
C43 S1 AND_3_magic_5.B 6.31e-20
C44 S4 S3 0.0092f
C45 A a_1091_2199# 9.99e-19
C46 B S3 6.31e-20
C47 C AND_3_magic_3.A 0.242f
C48 S1 AND_3_magic_5.C 0.00142f
C49 a_587_2199# a_252_1525# 1.36e-19
C50 VDD a_587_4113# 0.00684f
C51 a_439_5355# S2 0.0806f
C52 a_439_6016# a_439_5355# 0.00234f
C53 AND_3_magic_5.B a_439_3441# 5.39e-19
C54 a_587_2199# a_1091_2199# 0.32f
C55 AND_3_magic_5.C a_439_3441# 3.23e-19
C56 a_439_5355# a_1091_5366# 0.285f
C57 VDD a_439_5355# 1.07f
C58 AND_3_magic_5.C a_1091_4113# 0.502f
C59 AND_3_magic_3.A A 3.39f
C60 a_587_3452# a_439_3441# 0.475f
C61 a_439_6016# S2 8.31e-21
C62 B a_587_4113# 0.0549f
C63 C a_587_4113# 7.18e-20
C64 AND_3_magic_3.A a_439_4102# 0.193f
C65 AND_3_magic_5.B a_587_5366# 0.0548f
C66 a_439_4102# S3 0.0806f
C67 a_1091_5366# S2 0.0134f
C68 AND_3_magic_5.C a_587_5366# 5.8e-20
C69 a_439_3441# a_439_2188# 0.00531f
C70 VDD S2 0.247f
C71 a_439_6016# VDD 1.07f
C72 a_439_5355# B 6.46e-19
C73 AND_3_magic_3.A a_587_2199# 1.67e-19
C74 C a_439_5355# 0.111f
C75 VDD a_1091_5366# 0.00358f
C76 AND_3_magic_5.B AND_3_magic_5.C 2.36f
C77 A a_587_4113# 0.00272f
C78 a_439_6016# B 4.08e-19
C79 C S2 0.00142f
C80 C a_439_6016# 2.9e-19
C81 AND_3_magic_5.B a_587_3452# 1.3e-19
C82 a_439_4102# a_587_4113# 0.475f
C83 AND_3_magic_5.C a_587_3452# 5.8e-20
C84 VDD AND_1.A 0.361f
C85 a_587_6027# AND_3_magic_5.B 0.0548f
C86 VDD S4 0.247f
C87 VDD B 3.5f
C88 C a_1091_5366# 0.502f
C89 a_1091_6027# a_439_6016# 0.285f
C90 a_587_6027# AND_3_magic_5.C 0.457f
C91 A a_439_5355# 0.00654f
C92 C VDD 2.12f
C93 AND_3_magic_5.B a_439_2188# 0.0595f
C94 VDD a_1091_3452# 0.00358f
C95 AND_3_magic_5.C a_439_2188# 0.111f
C96 a_439_5355# a_439_4102# 0.00531f
C97 a_1091_6027# VDD 0.00358f
C98 VDD S5 0.248f
C99 B AND_1.A 0.00122f
C100 S4 B 6.31e-20
C101 a_439_6016# A 0.00654f
C102 C AND_1.A 8.36e-19
C103 C S4 0.00142f
C104 C B 1.26f
C105 a_1091_3452# S4 0.0134f
C106 S2 a_439_4102# 1.18e-19
C107 A a_1091_5366# 8.26e-19
C108 a_1091_3452# B 0.0355f
C109 VDD a_400_841# 0.219f
C110 AND_3_magic_5.C S6 6.62e-20
C111 VDD A 2.82f
C112 C a_1091_3452# 0.502f
C113 a_1091_6027# C 1.35e-19
C114 AND_3_magic_5.B a_1333_1282# 2.99e-19
C115 S4 S5 0.00185f
C116 VDD a_439_4102# 1.07f
C117 AND_3_magic_5.C a_1333_1282# 0.00137f
C118 AND_3_magic_5.B a_1185_1271# 3.64e-19
C119 AND_3_magic_5.C a_1185_1271# 4.78e-19
C120 AND_1.A a_400_841# 1.44e-19
C121 VDD a_587_2199# 0.00685f
C122 A AND_1.A 0.0959f
C123 B a_400_841# 0.0203f
C124 A B 0.237f
C125 C a_400_841# 0.0835f
C126 AND_3_magic_3.A a_439_3441# 0.193f
C127 AND_3_magic_5.B a_252_1525# 4.56e-19
C128 C A 1.48f
C129 S3 a_439_3441# 8.31e-21
C130 AND_3_magic_5.C a_252_1525# 4.13e-19
C131 S4 a_439_4102# 8.31e-21
C132 a_1091_3452# A 8.26e-19
C133 B a_439_4102# 0.0597f
C134 a_439_2188# a_1333_1282# 0.00149f
C135 C a_439_4102# 3.71e-19
C136 a_1091_6027# A 8.26e-19
C137 AND_3_magic_5.B a_1091_2199# 0.0349f
C138 S3 a_1091_4113# 0.0134f
C139 AND_3_magic_5.C a_1091_2199# 0.502f
C140 a_587_2199# AND_1.A 6.28e-20
C141 B a_587_2199# 1.58e-19
C142 C a_587_2199# 7.18e-20
C143 AND_3_magic_3.A a_587_5366# 0.0359f
C144 a_439_2188# a_252_1525# 1.04e-19
C145 A a_400_841# 0.00528f
C146 S1 a_439_5355# 8.31e-21
C147 a_1333_1282# S6 0.0742f
C148 a_439_2188# a_1091_2199# 0.285f
C149 A a_439_4102# 0.00654f
C150 a_1185_1271# S6 0.0315f
C151 AND_3_magic_5.B AND_3_magic_3.A 1.61f
C152 AND_3_magic_3.A AND_3_magic_5.C 0.237f
C153 AND_3_magic_5.C S3 0.00142f
C154 a_587_4113# a_1091_4113# 0.32f
C155 a_1185_1271# a_1333_1282# 0.319f
C156 A a_587_2199# 0.0379f
C157 S1 S2 0.0092f
C158 S1 a_439_6016# 0.0806f
C159 a_252_1525# S6 1.77e-20
C160 AND_3_magic_3.A a_587_3452# 0.0359f
C161 a_587_6027# AND_3_magic_3.A 0.0359f
C162 a_252_1525# a_1333_1282# 2.28e-19
C163 S1 VDD 0.247f
C164 AND_3_magic_3.A a_439_2188# 6.02e-19
C165 a_252_1525# a_1185_1271# 0.00119f
C166 a_439_5355# a_587_5366# 0.475f
C167 AND_3_magic_5.B a_587_4113# 1.3e-19
C168 AND_3_magic_5.C a_587_4113# 0.457f
C169 VDD a_439_3441# 1.07f
C170 AND_3_magic_5.B a_439_5355# 0.0596f
C171 VDD a_1091_4113# 0.00358f
C172 AND_3_magic_5.C a_439_5355# 3.23e-19
C173 S1 a_1091_6027# 0.0134f
C174 a_587_5366# a_1091_5366# 0.32f
C175 S4 a_439_3441# 0.0806f
C176 VDD a_587_5366# 0.00684f
C177 B a_439_3441# 0.0597f
C178 C a_439_3441# 0.111f
C179 AND_3_magic_5.B S2 6.31e-20
C180 AND_3_magic_5.B a_439_6016# 0.0596f
C181 a_1091_3452# a_439_3441# 0.285f
C182 B a_1091_4113# 0.0355f
C183 a_439_6016# AND_3_magic_5.C 0.111f
C184 C a_1091_4113# 2.06e-19
C185 AND_3_magic_5.B a_1091_5366# 0.0355f
C186 AND_3_magic_3.A a_252_1525# 0.00115f
C187 AND_3_magic_5.C a_1091_5366# 2.06e-19
C188 AND_3_magic_5.B VDD 2.53f
C189 a_439_3441# S5 1.18e-19
C190 AND_3_magic_5.C VDD 1.19f
C191 a_587_5366# B 1.58e-19
C192 C a_587_5366# 0.457f
C193 a_587_6027# a_439_6016# 0.475f
C194 VDD a_587_3452# 0.00684f
C195 A a_439_3441# 0.00654f
C196 a_587_6027# VDD 0.00684f
C197 AND_3_magic_5.B AND_1.A 0.00266f
C198 AND_3_magic_5.B B 3.51f
C199 AND_3_magic_5.C AND_1.A 8.84e-19
C200 a_439_4102# a_439_3441# 0.00234f
C201 A a_1091_4113# 8.26e-19
C202 AND_3_magic_5.C B 0.125f
C203 C AND_3_magic_5.B 3.18f
C204 VDD a_439_2188# 1.07f
C205 C AND_3_magic_5.C 3.62f
C206 a_439_4102# a_1091_4113# 0.285f
C207 AND_3_magic_5.C a_1091_3452# 2.06e-19
C208 a_1091_6027# AND_3_magic_5.B 0.0355f
C209 a_1091_6027# AND_3_magic_5.C 0.502f
C210 a_587_3452# B 0.0549f
C211 A a_587_5366# 0.00272f
C212 C a_587_3452# 0.457f
C213 AND_3_magic_5.B S5 6.31e-20
C214 a_587_6027# B 1.19e-19
C215 AND_3_magic_5.C S5 0.00142f
C216 a_587_3452# a_1091_3452# 0.32f
C217 a_587_6027# C 7.18e-20
C218 a_439_2188# AND_1.A 6.37e-20
C219 S4 a_439_2188# 1.18e-19
C220 B a_439_2188# 6.46e-19
C221 VDD S6 0.153f
C222 C a_439_2188# 3.88e-19
C223 a_587_6027# a_1091_6027# 0.32f
C224 AND_3_magic_5.B a_400_841# 4.52e-20
C225 AND_3_magic_5.B A 0.278f
C226 S6 VSS 0.482f
C227 a_1333_1282# VSS 0.492f
C228 a_1185_1271# VSS 0.714f
C229 a_400_841# VSS 0.00367f
C230 AND_1.A VSS 0.604f
C231 a_252_1525# VSS 0.627f
C232 a_1091_2199# VSS 0.369f
C233 a_587_2199# VSS 0.084f
C234 S5 VSS 0.368f
C235 a_439_2188# VSS 0.416f
C236 A VSS 4.96f
C237 S4 VSS 0.365f
C238 a_1091_3452# VSS 0.369f
C239 a_587_3452# VSS 0.084f
C240 a_439_3441# VSS 0.415f
C241 a_1091_4113# VSS 0.369f
C242 a_587_4113# VSS 0.084f
C243 S3 VSS 0.365f
C244 a_439_4102# VSS 0.415f
C245 B VSS 5.39f
C246 S2 VSS 0.365f
C247 a_1091_5366# VSS 0.369f
C248 a_587_5366# VSS 0.084f
C249 a_439_5355# VSS 0.415f
C250 C VSS 8.8f
C251 a_1091_6027# VSS 0.369f
C252 a_587_6027# VSS 0.084f
C253 S1 VSS 0.367f
C254 AND_3_magic_5.C VSS 11.9f
C255 a_439_6016# VSS 0.425f
C256 AND_3_magic_3.A VSS 6.7f
C257 AND_3_magic_5.B VSS 7.99f
C258 VDD VSS 26.5f
C259 AND_3_magic_5.C.t5 VSS -0.00196f
C260 AND_3_magic_5.C.t7 VSS 0.0273f
C261 AND_3_magic_5.C.n0 VSS 0.0513f
C262 AND_3_magic_5.C.t8 VSS 0.0368f
C263 AND_3_magic_5.C.t3 VSS 0.0926f
C264 AND_3_magic_5.C.t6 VSS 0.0617f
C265 AND_3_magic_5.C.n1 VSS 0.0745f
C266 AND_3_magic_5.C.t15 VSS -0.00196f
C267 AND_3_magic_5.C.t2 VSS 0.0273f
C268 AND_3_magic_5.C.n2 VSS 0.0513f
C269 AND_3_magic_5.C.t4 VSS 0.0368f
C270 AND_3_magic_5.C.t13 VSS 0.0926f
C271 AND_3_magic_5.C.t16 VSS 0.0617f
C272 AND_3_magic_5.C.n3 VSS 0.0745f
C273 AND_3_magic_5.C.n4 VSS 0.705f
C274 AND_3_magic_5.C.t10 VSS -0.00196f
C275 AND_3_magic_5.C.t12 VSS 0.0273f
C276 AND_3_magic_5.C.n5 VSS 0.0513f
C277 AND_3_magic_5.C.t14 VSS 0.0368f
C278 AND_3_magic_5.C.t9 VSS 0.0926f
C279 AND_3_magic_5.C.t11 VSS 0.0617f
C280 AND_3_magic_5.C.n6 VSS 0.0745f
C281 AND_3_magic_5.C.n7 VSS 1.54f
C282 B.t15 VSS 0.0155f
C283 B.t9 VSS 0.0656f
C284 B.n0 VSS 0.164f
C285 B.t16 VSS 0.15f
C286 B.t1 VSS 0.0186f
C287 B.t3 VSS -0.00493f
C288 B.t8 VSS 0.0673f
C289 B.n1 VSS 0.125f
C290 B.t6 VSS 0.0136f
C291 B.n2 VSS 0.125f
C292 B.n3 VSS 0.15f
C293 B.t5 VSS 0.361f
C294 B.n4 VSS 1.5f
C295 B.t12 VSS -0.00493f
C296 B.t14 VSS 0.0673f
C297 B.n5 VSS 0.125f
C298 B.t13 VSS 0.0136f
C299 B.n6 VSS 0.125f
C300 B.t17 VSS 0.0186f
C301 B.n7 VSS 0.15f
C302 B.t0 VSS 0.361f
C303 B.n8 VSS 1.54f
C304 B.t4 VSS 0.1f
C305 B.t10 VSS 0.164f
C306 B.t11 VSS 0.0997f
C307 B.t2 VSS 0.0997f
C308 B.t7 VSS 0.178f
C309 B.n9 VSS 1.03f
C310 B.n10 VSS 0.785f
C311 C.t8 VSS 0.0113f
C312 C.t1 VSS 0.0478f
C313 C.n0 VSS 0.119f
C314 C.t4 VSS 0.11f
C315 C.t13 VSS -0.00359f
C316 C.t16 VSS 0.0499f
C317 C.n1 VSS 0.094f
C318 C.t5 VSS 0.0674f
C319 C.t17 VSS 0.17f
C320 C.t14 VSS 0.113f
C321 C.n2 VSS 0.136f
C322 C.n3 VSS 0.946f
C323 C.t7 VSS -0.00359f
C324 C.t11 VSS 0.0499f
C325 C.n4 VSS 0.094f
C326 C.t0 VSS 0.0674f
C327 C.t12 VSS 0.17f
C328 C.t9 VSS 0.113f
C329 C.n5 VSS 0.136f
C330 C.n6 VSS 1.26f
C331 C.t2 VSS 0.0413f
C332 C.t3 VSS 0.0254f
C333 C.t15 VSS 0.0727f
C334 C.t10 VSS 0.0727f
C335 C.t6 VSS 0.0636f
C336 C.n7 VSS 0.133f
C337 C.n8 VSS 1.24f
C338 A.t10 VSS 0.0115f
C339 A.t7 VSS 0.0484f
C340 A.n0 VSS 0.121f
C341 A.t2 VSS 0.111f
C342 A.t9 VSS 0.0505f
C343 A.t1 VSS 0.014f
C344 A.n1 VSS 0.073f
C345 A.t8 VSS 0.0491f
C346 A.t0 VSS 0.0129f
C347 A.n2 VSS 0.0914f
C348 A.t4 VSS 0.0129f
C349 A.n3 VSS 0.0798f
C350 A.n4 VSS 0.0817f
C351 A.n5 VSS 1.77f
C352 A.t6 VSS 0.0574f
C353 A.t5 VSS 0.0188f
C354 A.n6 VSS 0.156f
C355 A.t3 VSS 0.221f
C356 A.n7 VSS 0.855f
C357 AND_3_magic_5.B.t6 VSS 0.0162f
C358 AND_3_magic_5.B.t7 VSS -0.00429f
C359 AND_3_magic_5.B.t10 VSS 0.0585f
C360 AND_3_magic_5.B.n0 VSS 0.109f
C361 AND_3_magic_5.B.t9 VSS 0.0119f
C362 AND_3_magic_5.B.n1 VSS 0.109f
C363 AND_3_magic_5.B.n2 VSS 0.13f
C364 AND_3_magic_5.B.t8 VSS 0.314f
C365 AND_3_magic_5.B.t16 VSS -0.00429f
C366 AND_3_magic_5.B.t3 VSS 0.0585f
C367 AND_3_magic_5.B.n3 VSS 0.109f
C368 AND_3_magic_5.B.t2 VSS 0.0119f
C369 AND_3_magic_5.B.n4 VSS 0.109f
C370 AND_3_magic_5.B.t4 VSS 0.0162f
C371 AND_3_magic_5.B.n5 VSS 0.13f
C372 AND_3_magic_5.B.t5 VSS 0.314f
C373 AND_3_magic_5.B.n6 VSS 1.66f
C374 AND_3_magic_5.B.t11 VSS 0.0162f
C375 AND_3_magic_5.B.t12 VSS -0.00429f
C376 AND_3_magic_5.B.t15 VSS 0.0585f
C377 AND_3_magic_5.B.n7 VSS 0.109f
C378 AND_3_magic_5.B.t13 VSS 0.0119f
C379 AND_3_magic_5.B.n8 VSS 0.109f
C380 AND_3_magic_5.B.n9 VSS 0.13f
C381 AND_3_magic_5.B.t14 VSS 0.314f
C382 AND_3_magic_5.B.n10 VSS 3.3f
C383 VDD.t37 VSS 0.00169f
C384 VDD.n0 VSS 0.00169f
C385 VDD.n1 VSS 0.00574f
C386 VDD.n2 VSS 0.00385f
C387 VDD.t79 VSS 0.00169f
C388 VDD.n3 VSS 0.0054f
C389 VDD.t65 VSS 0.00337f
C390 VDD.n4 VSS 0.00169f
C391 VDD.n5 VSS 0.0054f
C392 VDD.t63 VSS 0.00406f
C393 VDD.n6 VSS 0.0353f
C394 VDD.t101 VSS 0.00169f
C395 VDD.n7 VSS 0.0054f
C396 VDD.t60 VSS 0.00337f
C397 VDD.n8 VSS 0.00169f
C398 VDD.n9 VSS 0.0054f
C399 VDD.t58 VSS 0.00406f
C400 VDD.n10 VSS 0.0353f
C401 VDD.t90 VSS 0.00169f
C402 VDD.n11 VSS 0.00169f
C403 VDD.n12 VSS 0.00604f
C404 VDD.t1 VSS 0.00385f
C405 VDD.n13 VSS 0.0921f
C406 VDD.t0 VSS 0.0352f
C407 VDD.n14 VSS 0.0622f
C408 VDD.n15 VSS 0.00966f
C409 VDD.n16 VSS 0.00959f
C410 VDD.n17 VSS 0.0502f
C411 VDD.n18 VSS 0.00966f
C412 VDD.n19 VSS 0.0126f
C413 VDD.t2 VSS 0.0329f
C414 VDD.n20 VSS 0.0404f
C415 VDD.n21 VSS 0.00966f
C416 VDD.n22 VSS 0.00971f
C417 VDD.n23 VSS 0.0199f
C418 VDD.t89 VSS 0.0329f
C419 VDD.n24 VSS 0.0428f
C420 VDD.n25 VSS 0.00966f
C421 VDD.n26 VSS 0.00925f
C422 VDD.n27 VSS 0.0502f
C423 VDD.n28 VSS 0.00966f
C424 VDD.n29 VSS 0.0126f
C425 VDD.t86 VSS 0.0329f
C426 VDD.n30 VSS 0.0386f
C427 VDD.n31 VSS 0.00966f
C428 VDD.n32 VSS 0.0126f
C429 VDD.t59 VSS 0.0329f
C430 VDD.n33 VSS 0.0446f
C431 VDD.n34 VSS 0.00966f
C432 VDD.n35 VSS 0.00856f
C433 VDD.n36 VSS 0.0086f
C434 VDD.n37 VSS 0.00419f
C435 VDD.n38 VSS 0.0502f
C436 VDD.n39 VSS 0.00966f
C437 VDD.t100 VSS 0.0329f
C438 VDD.n40 VSS 0.0368f
C439 VDD.n41 VSS 0.00966f
C440 VDD.n42 VSS 0.0125f
C441 VDD.t109 VSS 0.0329f
C442 VDD.n43 VSS 0.0464f
C443 VDD.n44 VSS 0.00966f
C444 VDD.n45 VSS 0.0126f
C445 VDD.n46 VSS 0.0502f
C446 VDD.n47 VSS 0.00966f
C447 VDD.n48 VSS 0.0122f
C448 VDD.n49 VSS 0.0086f
C449 VDD.t64 VSS 0.0329f
C450 VDD.n50 VSS 0.035f
C451 VDD.n51 VSS 0.00966f
C452 VDD.n52 VSS 0.00672f
C453 VDD.t78 VSS 0.0329f
C454 VDD.n53 VSS 0.0481f
C455 VDD.n54 VSS 0.00966f
C456 VDD.n55 VSS 0.0126f
C457 VDD.n56 VSS 0.0502f
C458 VDD.n57 VSS 0.00966f
C459 VDD.n58 VSS 0.0126f
C460 VDD.t75 VSS 0.0541f
C461 VDD.n59 VSS 0.0402f
C462 VDD.n60 VSS 0.00966f
C463 VDD.n61 VSS 0.0111f
C464 VDD.n62 VSS 0.0244f
C465 VDD.n63 VSS 0.104f
C466 VDD.n64 VSS 0.0824f
C467 VDD.n65 VSS 0.00385f
C468 VDD.n66 VSS 0.00385f
C469 VDD.t140 VSS 0.00169f
C470 VDD.t43 VSS 0.00337f
C471 VDD.n67 VSS 0.0054f
C472 VDD.n68 VSS 0.00169f
C473 VDD.n69 VSS 0.0054f
C474 VDD.t41 VSS 0.00406f
C475 VDD.n70 VSS 0.0353f
C476 VDD.t71 VSS 0.00169f
C477 VDD.t48 VSS 0.00337f
C478 VDD.n71 VSS 0.0054f
C479 VDD.n72 VSS 0.00169f
C480 VDD.n73 VSS 0.0054f
C481 VDD.t47 VSS 0.00406f
C482 VDD.n74 VSS 0.0353f
C483 VDD.t35 VSS 0.00169f
C484 VDD.t62 VSS 0.00337f
C485 VDD.n75 VSS 0.0054f
C486 VDD.n76 VSS 0.00169f
C487 VDD.n77 VSS 0.0054f
C488 VDD.t61 VSS 0.00406f
C489 VDD.n78 VSS 0.0353f
C490 VDD.t112 VSS 0.00169f
C491 VDD.t40 VSS 0.00337f
C492 VDD.n79 VSS 0.0054f
C493 VDD.n80 VSS 0.00169f
C494 VDD.n81 VSS 0.0054f
C495 VDD.t38 VSS 0.00406f
C496 VDD.n82 VSS 0.0353f
C497 VDD.t85 VSS 0.00169f
C498 VDD.n83 VSS 0.00169f
C499 VDD.n84 VSS 0.00604f
C500 VDD.t141 VSS 0.00169f
C501 VDD.n85 VSS 0.00169f
C502 VDD.n86 VSS 0.00604f
C503 VDD.t6 VSS 0.00385f
C504 VDD.t9 VSS 0.00385f
C505 VDD.n87 VSS 0.146f
C506 VDD.t5 VSS 0.0629f
C507 VDD.n88 VSS 0.105f
C508 VDD.n89 VSS 0.00979f
C509 VDD.n90 VSS 0.00969f
C510 VDD.n91 VSS 0.0862f
C511 VDD.n92 VSS 0.00979f
C512 VDD.n93 VSS 0.0128f
C513 VDD.t7 VSS 0.0564f
C514 VDD.n94 VSS 0.0693f
C515 VDD.n95 VSS 0.00979f
C516 VDD.n96 VSS 0.0098f
C517 VDD.n97 VSS 0.0336f
C518 VDD.t84 VSS 0.0564f
C519 VDD.n98 VSS 0.0734f
C520 VDD.n99 VSS 0.00979f
C521 VDD.n100 VSS 0.00934f
C522 VDD.n101 VSS 0.0862f
C523 VDD.n102 VSS 0.00979f
C524 VDD.n103 VSS 0.0128f
C525 VDD.t22 VSS 0.0564f
C526 VDD.n104 VSS 0.0662f
C527 VDD.n105 VSS 0.00979f
C528 VDD.n106 VSS 0.0128f
C529 VDD.t39 VSS 0.0564f
C530 VDD.n107 VSS 0.0764f
C531 VDD.n108 VSS 0.00979f
C532 VDD.n109 VSS 0.00864f
C533 VDD.n110 VSS 0.0109f
C534 VDD.n111 VSS 0.00423f
C535 VDD.n112 VSS 0.0862f
C536 VDD.n113 VSS 0.00979f
C537 VDD.t34 VSS 0.0564f
C538 VDD.n114 VSS 0.0631f
C539 VDD.n115 VSS 0.00979f
C540 VDD.n116 VSS 0.0126f
C541 VDD.t91 VSS 0.0564f
C542 VDD.n117 VSS 0.0795f
C543 VDD.n118 VSS 0.00979f
C544 VDD.n119 VSS 0.0128f
C545 VDD.n120 VSS 0.0862f
C546 VDD.n121 VSS 0.00979f
C547 VDD.n122 VSS 0.0124f
C548 VDD.n123 VSS 0.0109f
C549 VDD.t42 VSS 0.0564f
C550 VDD.n124 VSS 0.06f
C551 VDD.n125 VSS 0.00979f
C552 VDD.n126 VSS 0.00679f
C553 VDD.t70 VSS 0.0564f
C554 VDD.n127 VSS 0.0826f
C555 VDD.n128 VSS 0.00979f
C556 VDD.n129 VSS 0.0128f
C557 VDD.n130 VSS 0.0862f
C558 VDD.n131 VSS 0.00979f
C559 VDD.n132 VSS 0.0128f
C560 VDD.t72 VSS 0.1f
C561 VDD.n133 VSS 0.062f
C562 VDD.n134 VSS 0.00979f
C563 VDD.n135 VSS 0.0112f
C564 VDD.n136 VSS 0.0425f
C565 VDD.n137 VSS 0.148f
C566 VDD.n138 VSS 0.156f
C567 VDD.n139 VSS 0.00385f
C568 VDD.n140 VSS 0.00385f
C569 VDD.t114 VSS 0.00169f
C570 VDD.t53 VSS 0.00337f
C571 VDD.n141 VSS 0.0054f
C572 VDD.n142 VSS 0.00169f
C573 VDD.n143 VSS 0.0054f
C574 VDD.t51 VSS 0.00406f
C575 VDD.n144 VSS 0.0353f
C576 VDD.t120 VSS 0.00169f
C577 VDD.n145 VSS 0.0054f
C578 VDD.t57 VSS 0.00337f
C579 VDD.n146 VSS 0.00169f
C580 VDD.n147 VSS 0.0054f
C581 VDD.t56 VSS 0.00406f
C582 VDD.n148 VSS 0.0353f
C583 VDD.t81 VSS 0.00169f
C584 VDD.t46 VSS 0.00337f
C585 VDD.n149 VSS 0.0054f
C586 VDD.n150 VSS 0.00169f
C587 VDD.n151 VSS 0.0054f
C588 VDD.t44 VSS 0.00406f
C589 VDD.n152 VSS 0.0353f
C590 VDD.t123 VSS 0.00169f
C591 VDD.t50 VSS 0.00337f
C592 VDD.n153 VSS 0.0054f
C593 VDD.n154 VSS 0.00169f
C594 VDD.n155 VSS 0.0054f
C595 VDD.t49 VSS 0.00406f
C596 VDD.n156 VSS 0.0353f
C597 VDD.t21 VSS 0.00169f
C598 VDD.n157 VSS 0.00169f
C599 VDD.n158 VSS 0.00604f
C600 VDD.t69 VSS 0.00169f
C601 VDD.n159 VSS 0.00169f
C602 VDD.n160 VSS 0.00604f
C603 VDD.t14 VSS 0.00385f
C604 VDD.t105 VSS 0.00385f
C605 VDD.n161 VSS 0.146f
C606 VDD.t13 VSS 0.0629f
C607 VDD.n162 VSS 0.105f
C608 VDD.n163 VSS 0.00979f
C609 VDD.n164 VSS 0.00969f
C610 VDD.n165 VSS 0.0862f
C611 VDD.n166 VSS 0.00979f
C612 VDD.n167 VSS 0.0128f
C613 VDD.t15 VSS 0.0564f
C614 VDD.n168 VSS 0.0693f
C615 VDD.n169 VSS 0.00979f
C616 VDD.n170 VSS 0.0098f
C617 VDD.n171 VSS 0.0336f
C618 VDD.t20 VSS 0.0564f
C619 VDD.n172 VSS 0.0734f
C620 VDD.n173 VSS 0.00979f
C621 VDD.n174 VSS 0.00934f
C622 VDD.n175 VSS 0.0862f
C623 VDD.n176 VSS 0.00979f
C624 VDD.n177 VSS 0.0128f
C625 VDD.t66 VSS 0.0564f
C626 VDD.n178 VSS 0.0662f
C627 VDD.n179 VSS 0.00979f
C628 VDD.n180 VSS 0.0128f
C629 VDD.t45 VSS 0.0564f
C630 VDD.n181 VSS 0.0764f
C631 VDD.n182 VSS 0.00979f
C632 VDD.n183 VSS 0.00864f
C633 VDD.n184 VSS 0.0109f
C634 VDD.n185 VSS 0.00423f
C635 VDD.n186 VSS 0.0862f
C636 VDD.n187 VSS 0.00979f
C637 VDD.t80 VSS 0.0564f
C638 VDD.n188 VSS 0.0631f
C639 VDD.n189 VSS 0.00979f
C640 VDD.n190 VSS 0.0126f
C641 VDD.t102 VSS 0.0564f
C642 VDD.n191 VSS 0.0795f
C643 VDD.n192 VSS 0.00979f
C644 VDD.n193 VSS 0.0128f
C645 VDD.n194 VSS 0.0862f
C646 VDD.n195 VSS 0.00979f
C647 VDD.n196 VSS 0.0124f
C648 VDD.n197 VSS 0.0109f
C649 VDD.t52 VSS 0.0564f
C650 VDD.n198 VSS 0.06f
C651 VDD.n199 VSS 0.00979f
C652 VDD.n200 VSS 0.00679f
C653 VDD.t113 VSS 0.0564f
C654 VDD.n201 VSS 0.0826f
C655 VDD.n202 VSS 0.00979f
C656 VDD.n203 VSS 0.0128f
C657 VDD.n204 VSS 0.0862f
C658 VDD.n205 VSS 0.00979f
C659 VDD.n206 VSS 0.0128f
C660 VDD.t115 VSS 0.1f
C661 VDD.n207 VSS 0.062f
C662 VDD.n208 VSS 0.00979f
C663 VDD.n209 VSS 0.0112f
C664 VDD.n210 VSS 0.0425f
C665 VDD.n211 VSS 0.146f
C666 VDD.n212 VSS 0.199f
C667 VDD.n213 VSS 0.103f
C668 VDD.t36 VSS 0.0315f
C669 VDD.n214 VSS 0.0528f
C670 VDD.n215 VSS 0.009f
C671 VDD.n216 VSS 0.00973f
C672 VDD.n217 VSS 0.017f
C673 VDD.t18 VSS 0.0799f
C674 VDD.t19 VSS 0.00293f
C675 VDD.n218 VSS 0.00293f
C676 VDD.n219 VSS 0.00733f
C677 VDD.t135 VSS 0.0507f
C678 VDD.n220 VSS 0.057f
C679 VDD.t99 VSS 0.00682f
C680 VDD.t98 VSS 0.0829f
C681 VDD.t29 VSS 0.00346f
C682 VDD.t28 VSS 0.00323f
C683 VDD.n221 VSS 0.0276f
C684 VDD.t55 VSS 0.00676f
C685 VDD.n222 VSS 0.0133f
C686 VDD.t54 VSS 0.00387f
C687 VDD.n223 VSS 0.0308f
C688 VDD.t96 VSS 0.00346f
C689 VDD.t97 VSS 0.00323f
C690 VDD.n224 VSS 0.0209f
C691 VDD.t26 VSS 0.00323f
C692 VDD.n225 VSS 0.0117f
C693 VDD.t142 VSS 0.00323f
C694 VDD.n226 VSS 0.0134f
C695 VDD.n227 VSS 0.123f
C696 VDD.t25 VSS 0.0729f
C697 VDD.n228 VSS 0.0957f
C698 VDD.n229 VSS 0.0119f
C699 VDD.n230 VSS 0.0125f
C700 VDD.t30 VSS 0.0608f
C701 VDD.n231 VSS 0.083f
C702 VDD.n232 VSS 0.0119f
C703 VDD.n233 VSS 0.0158f
C704 VDD.n234 VSS 0.00803f
C705 VDD.n235 VSS 0.0934f
C706 VDD.n236 VSS 0.0119f
C707 VDD.n237 VSS 0.117f
C708 VDD.n238 VSS 0.0119f
C709 VDD.n239 VSS 0.015f
C710 VDD.n240 VSS 0.00911f
C711 VDD.t27 VSS 0.0747f
C712 VDD.n241 VSS 0.0932f
C713 VDD.n242 VSS 0.0119f
C714 VDD.n243 VSS 0.00854f
C715 VDD.n244 VSS 0.125f
C716 VDD.n245 VSS 0.129f
C717 VDD.n246 VSS 0.0343f
C718 VDD.n247 VSS 0.0142f
C719 VDD.n248 VSS 0.0309f
C720 VDD.n249 VSS 0.151f
C721 VDD.t129 VSS 0.00169f
C722 VDD.n250 VSS 0.00169f
C723 VDD.n251 VSS 0.00574f
C724 VDD.n252 VSS 0.017f
C725 VDD.t130 VSS 0.0308f
C726 VDD.n253 VSS 0.0546f
C727 VDD.n254 VSS 0.009f
C728 VDD.t127 VSS 0.00169f
C729 VDD.n255 VSS 0.00169f
C730 VDD.n256 VSS 0.00574f
C731 VDD.n257 VSS 0.017f
C732 VDD.t106 VSS 0.0324f
C733 VDD.n258 VSS 0.066f
C734 VDD.n259 VSS 0.0443f
C735 VDD.n260 VSS 0.00902f
C736 VDD.t126 VSS 0.0315f
C737 VDD.n261 VSS 0.0528f
C738 VDD.n262 VSS 0.009f
C739 VDD.n263 VSS 0.00973f
C740 VDD.n264 VSS 0.072f
C741 VDD.n265 VSS 0.0661f
C742 VDD.n266 VSS 0.01f
C743 VDD.n267 VSS 0.0443f
C744 VDD.n268 VSS 0.009f
C745 VDD.t128 VSS 0.0315f
C746 VDD.n269 VSS 0.0528f
C747 VDD.n270 VSS 0.009f
C748 VDD.n271 VSS 0.00973f
C749 VDD.n272 VSS 0.072f
C750 VDD.n273 VSS 0.0661f
C751 VDD.t31 VSS 0.0308f
C752 VDD.n274 VSS 0.0546f
C753 VDD.n275 VSS 0.009f
C754 VDD.n276 VSS 0.00775f
C755 VDD.n277 VSS 0.02f
C756 VDD.n278 VSS 0.0443f
C757 VDD.n279 VSS 0.009f
C758 AND_3_magic_3.A.t15 VSS 0.0399f
C759 AND_3_magic_3.A.t17 VSS 0.0111f
C760 AND_3_magic_3.A.n0 VSS 0.0576f
C761 AND_3_magic_3.A.t16 VSS 0.0388f
C762 AND_3_magic_3.A.t18 VSS 0.0102f
C763 AND_3_magic_3.A.n1 VSS 0.0722f
C764 AND_3_magic_3.A.t19 VSS 0.0102f
C765 AND_3_magic_3.A.n2 VSS 0.063f
C766 AND_3_magic_3.A.n3 VSS 0.0645f
C767 AND_3_magic_3.A.t4 VSS 0.0388f
C768 AND_3_magic_3.A.t6 VSS 0.0102f
C769 AND_3_magic_3.A.n4 VSS 0.0722f
C770 AND_3_magic_3.A.t8 VSS 0.0102f
C771 AND_3_magic_3.A.n5 VSS 0.063f
C772 AND_3_magic_3.A.t12 VSS 0.0399f
C773 AND_3_magic_3.A.t14 VSS 0.0108f
C774 AND_3_magic_3.A.n6 VSS 0.0576f
C775 AND_3_magic_3.A.n7 VSS 0.0648f
C776 AND_3_magic_3.A.n8 VSS 0.519f
C777 AND_3_magic_3.A.t7 VSS 0.0399f
C778 AND_3_magic_3.A.t10 VSS 0.0111f
C779 AND_3_magic_3.A.n9 VSS 0.0576f
C780 AND_3_magic_3.A.t9 VSS 0.0388f
C781 AND_3_magic_3.A.t11 VSS 0.0102f
C782 AND_3_magic_3.A.n10 VSS 0.0722f
C783 AND_3_magic_3.A.t13 VSS 0.0102f
C784 AND_3_magic_3.A.n11 VSS 0.063f
C785 AND_3_magic_3.A.n12 VSS 0.0645f
C786 AND_3_magic_3.A.n13 VSS 0.459f
C787 AND_3_magic_3.A.t20 VSS 0.0388f
C788 AND_3_magic_3.A.t21 VSS 0.0102f
C789 AND_3_magic_3.A.n14 VSS 0.0722f
C790 AND_3_magic_3.A.t2 VSS 0.0102f
C791 AND_3_magic_3.A.n15 VSS 0.063f
C792 AND_3_magic_3.A.t3 VSS 0.0399f
C793 AND_3_magic_3.A.t5 VSS 0.0108f
C794 AND_3_magic_3.A.n16 VSS 0.0576f
C795 AND_3_magic_3.A.n17 VSS 0.0648f
C796 AND_3_magic_3.A.n18 VSS 1.84f
.ends

