* NGSPICE file created from LF_mag_flat.ext - technology: gf180mcuC

.subckt LF_mag_flat VSS VDD VCNTL
X0 cap80p_mag_0.P VSS.t64 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X1 cap80p_mag_0.P VSS.t63 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X2 cap80p_mag_0.P VSS.t62 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X3 cap80p_mag_0.P VSS.t61 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X4 cap80p_mag_0.P VSS.t60 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X5 cap80p_mag_0.P VSS.t59 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X6 a_45980_43837# a_45740_41735# VDD.t9 ppolyf_u r_width=0.8u r_length=10u
X7 cap80p_mag_0.P VSS.t58 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X8 cap80p_mag_0.P VSS.t57 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X9 cap80p_mag_0.P VSS.t56 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X10 a_45980_43837# a_46220_41735# VDD.t4 ppolyf_u r_width=0.8u r_length=10u
X11 cap80p_mag_0.P VSS.t55 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X12 a_46460_43837# a_46700_41735# VDD.t1 ppolyf_u r_width=0.8u r_length=10u
X13 cap80p_mag_0.P VSS.t54 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X14 cap80p_mag_0.P VSS.t53 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X15 VCNTL.t0 a_45740_41735# VDD.t0 ppolyf_u r_width=0.8u r_length=10u
X16 cap80p_mag_0.P VSS.t52 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X17 cap80p_mag_0.P VSS.t51 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X18 cap80p_mag_0.P VSS.t50 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X19 cap80p_mag_0.P VSS.t49 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X20 cap80p_mag_0.P VSS.t48 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X21 cap80p_mag_0.P VSS.t47 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X22 cap80p_mag_0.P VSS.t46 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X23 cap80p_mag_0.P VSS.t45 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X24 cap80p_mag_0.P VSS.t44 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X25 cap80p_mag_0.P VSS.t43 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X26 cap80p_mag_0.P VSS.t42 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X27 cap80p_mag_0.P VSS.t41 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X28 cap80p_mag_0.P VSS.t40 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X29 VCNTL.t1 VSS.t0 cap_mim_2f0_m4m5_noshield c_width=42.5u c_length=42.5u
X30 cap80p_mag_0.P VSS.t39 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X31 cap80p_mag_0.P VSS.t38 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X32 cap80p_mag_0.P VSS.t37 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X33 cap80p_mag_0.P VSS.t36 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X34 cap80p_mag_0.P VSS.t35 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X35 cap80p_mag_0.P VSS.t34 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X36 cap80p_mag_0.P VSS.t33 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X37 cap80p_mag_0.P VSS.t32 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X38 cap80p_mag_0.P VSS.t31 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X39 cap80p_mag_0.P VSS.t30 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X40 cap80p_mag_0.P VSS.t29 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X41 cap80p_mag_0.P VSS.t28 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X42 cap80p_mag_0.P VSS.t27 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X43 cap80p_mag_0.P VSS.t26 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X44 cap80p_mag_0.P VSS.t25 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X45 cap80p_mag_0.P VSS.t24 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X46 cap80p_mag_0.P VSS.t23 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X47 a_46940_43837# a_47180_41735# VDD.t5 ppolyf_u r_width=0.8u r_length=10u
X48 cap80p_mag_0.P VSS.t22 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X49 cap80p_mag_0.P VSS.t21 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X50 cap80p_mag_0.P VSS.t20 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X51 cap80p_mag_0.P VSS.t19 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X52 a_47420_43837# a_47660_41735# VDD.t3 ppolyf_u r_width=0.8u r_length=10u
X53 cap80p_mag_0.P VSS.t18 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X54 cap80p_mag_0.P VSS.t17 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X55 cap80p_mag_0.P VSS.t16 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X56 cap80p_mag_0.P VSS.t15 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X57 cap80p_mag_0.P VSS.t14 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X58 cap80p_mag_0.P VSS.t13 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X59 cap80p_mag_0.P VSS.t12 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X60 cap80p_mag_0.P VSS.t11 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X61 cap80p_mag_0.P VSS.t10 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X62 cap80p_mag_0.P VSS.t9 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X63 a_47420_43837# a_47180_41735# VDD.t6 ppolyf_u r_width=0.8u r_length=10u
X64 cap80p_mag_0.P VSS.t8 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X65 cap80p_mag_0.P a_47660_41735# VDD.t8 ppolyf_u r_width=0.8u r_length=10u
X66 cap80p_mag_0.P VSS.t7 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X67 cap80p_mag_0.P VSS.t6 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X68 cap80p_mag_0.P VSS.t5 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X69 a_46460_43837# a_46220_41735# VDD.t7 ppolyf_u r_width=0.8u r_length=10u
X70 cap80p_mag_0.P VSS.t4 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X71 cap80p_mag_0.P VSS.t3 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X72 cap80p_mag_0.P VSS.t2 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X73 cap80p_mag_0.P VSS.t1 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X74 a_46940_43837# a_46700_41735# VDD.t2 ppolyf_u r_width=0.8u r_length=10u
R0 VSS.n74 VSS 13.3173
R1 VSS.n67 VSS.n0 4.53825
R2 VSS.n72 VSS.n2 4.52915
R3 VSS.n73 VSS.n0 4.52872
R4 VSS VSS.n2 4.52418
R5 VSS.n71 VSS.n70 4.5005
R6 VSS.n73 VSS.n1 4.5005
R7 VSS.n74 VSS.t0 4.37478
R8 VSS VSS.n73 4.32389
R9 VSS.n24 VSS.t49 3.26618
R10 VSS.n17 VSS.t22 3.26618
R11 VSS.n10 VSS.t43 3.26618
R12 VSS.n3 VSS.t50 3.26618
R13 VSS.n34 VSS.t48 3.26618
R14 VSS.n41 VSS.t44 3.26618
R15 VSS.n48 VSS.t26 3.26618
R16 VSS.n55 VSS.t52 3.26618
R17 VSS.n24 VSS.t41 2.25486
R18 VSS.n25 VSS.t12 2.25486
R19 VSS.n26 VSS.t63 2.25486
R20 VSS.n27 VSS.t28 2.25486
R21 VSS.n28 VSS.t32 2.25486
R22 VSS.n29 VSS.t7 2.25486
R23 VSS.n30 VSS.t14 2.25486
R24 VSS.n17 VSS.t11 2.25486
R25 VSS.n18 VSS.t47 2.25486
R26 VSS.n19 VSS.t39 2.25486
R27 VSS.n20 VSS.t56 2.25486
R28 VSS.n21 VSS.t61 2.25486
R29 VSS.n22 VSS.t31 2.25486
R30 VSS.n23 VSS.t38 2.25486
R31 VSS.n10 VSS.t35 2.25486
R32 VSS.n11 VSS.t3 2.25486
R33 VSS.n12 VSS.t53 2.25486
R34 VSS.n13 VSS.t20 2.25486
R35 VSS.n14 VSS.t24 2.25486
R36 VSS.n15 VSS.t8 2.25486
R37 VSS.n16 VSS.t15 2.25486
R38 VSS.n3 VSS.t42 2.25486
R39 VSS.n4 VSS.t13 2.25486
R40 VSS.n5 VSS.t64 2.25486
R41 VSS.n6 VSS.t29 2.25486
R42 VSS.n7 VSS.t33 2.25486
R43 VSS.n8 VSS.t57 2.25486
R44 VSS.n9 VSS.t5 2.25486
R45 VSS.n34 VSS.t40 2.25486
R46 VSS.n35 VSS.t10 2.25486
R47 VSS.n36 VSS.t58 2.25486
R48 VSS.n37 VSS.t27 2.25486
R49 VSS.n38 VSS.t30 2.25486
R50 VSS.n39 VSS.t16 2.25486
R51 VSS.n40 VSS.t23 2.25486
R52 VSS.n41 VSS.t36 2.25486
R53 VSS.n42 VSS.t4 2.25486
R54 VSS.n43 VSS.t54 2.25486
R55 VSS.n44 VSS.t21 2.25486
R56 VSS.n45 VSS.t25 2.25486
R57 VSS.n46 VSS.t60 2.25486
R58 VSS.n47 VSS.t6 2.25486
R59 VSS.n48 VSS.t17 2.25486
R60 VSS.n49 VSS.t51 2.25486
R61 VSS.n50 VSS.t45 2.25486
R62 VSS.n51 VSS.t62 2.25486
R63 VSS.n52 VSS.t1 2.25486
R64 VSS.n53 VSS.t9 2.25486
R65 VSS.n54 VSS.t19 2.25486
R66 VSS.n55 VSS.t46 2.25486
R67 VSS.n56 VSS.t18 2.25486
R68 VSS.n57 VSS.t2 2.25486
R69 VSS.n58 VSS.t34 2.25486
R70 VSS.n59 VSS.t37 2.25486
R71 VSS.n60 VSS.t55 2.25486
R72 VSS.n61 VSS.t59 2.25486
R73 VSS.n31 VSS.n30 1.63171
R74 VSS.n62 VSS.n61 1.6308
R75 VSS.n69 VSS.n68 1.5005
R76 VSS.n73 VSS.n72 1.1247
R77 VSS.n33 VSS.n32 1.07514
R78 VSS.n64 VSS.n63 1.07514
R79 VSS.n32 VSS.n31 1.07476
R80 VSS.n63 VSS.n62 1.07438
R81 VSS.n25 VSS.n24 1.01182
R82 VSS.n26 VSS.n25 1.01182
R83 VSS.n27 VSS.n26 1.01182
R84 VSS.n28 VSS.n27 1.01182
R85 VSS.n29 VSS.n28 1.01182
R86 VSS.n30 VSS.n29 1.01182
R87 VSS.n18 VSS.n17 1.01182
R88 VSS.n19 VSS.n18 1.01182
R89 VSS.n20 VSS.n19 1.01182
R90 VSS.n21 VSS.n20 1.01182
R91 VSS.n22 VSS.n21 1.01182
R92 VSS.n23 VSS.n22 1.01182
R93 VSS.n11 VSS.n10 1.01182
R94 VSS.n12 VSS.n11 1.01182
R95 VSS.n13 VSS.n12 1.01182
R96 VSS.n14 VSS.n13 1.01182
R97 VSS.n15 VSS.n14 1.01182
R98 VSS.n16 VSS.n15 1.01182
R99 VSS.n4 VSS.n3 1.01182
R100 VSS.n5 VSS.n4 1.01182
R101 VSS.n6 VSS.n5 1.01182
R102 VSS.n7 VSS.n6 1.01182
R103 VSS.n8 VSS.n7 1.01182
R104 VSS.n9 VSS.n8 1.01182
R105 VSS.n35 VSS.n34 1.01182
R106 VSS.n36 VSS.n35 1.01182
R107 VSS.n37 VSS.n36 1.01182
R108 VSS.n38 VSS.n37 1.01182
R109 VSS.n39 VSS.n38 1.01182
R110 VSS.n40 VSS.n39 1.01182
R111 VSS.n42 VSS.n41 1.01182
R112 VSS.n43 VSS.n42 1.01182
R113 VSS.n44 VSS.n43 1.01182
R114 VSS.n45 VSS.n44 1.01182
R115 VSS.n46 VSS.n45 1.01182
R116 VSS.n47 VSS.n46 1.01182
R117 VSS.n49 VSS.n48 1.01182
R118 VSS.n50 VSS.n49 1.01182
R119 VSS.n51 VSS.n50 1.01182
R120 VSS.n52 VSS.n51 1.01182
R121 VSS.n53 VSS.n52 1.01182
R122 VSS.n54 VSS.n53 1.01182
R123 VSS.n56 VSS.n55 1.01182
R124 VSS.n57 VSS.n56 1.01182
R125 VSS.n58 VSS.n57 1.01182
R126 VSS.n59 VSS.n58 1.01182
R127 VSS.n60 VSS.n59 1.01182
R128 VSS.n61 VSS.n60 1.01182
R129 VSS.n67 VSS.n66 0.898925
R130 VSS.n66 VSS.n65 0.71213
R131 VSS.n31 VSS.n23 0.556878
R132 VSS.n32 VSS.n16 0.556878
R133 VSS.n33 VSS.n9 0.556878
R134 VSS.n64 VSS.n40 0.556878
R135 VSS.n63 VSS.n47 0.556878
R136 VSS.n62 VSS.n54 0.556878
R137 VSS.n65 VSS.n33 0.539639
R138 VSS.n65 VSS.n64 0.53562
R139 VSS.n70 VSS.n2 0.0357703
R140 VSS.n68 VSS.n0 0.0267703
R141 VSS.n69 VSS.n67 0.008809
R142 VSS.n72 VSS.n71 0.00798833
R143 VSS.n70 VSS.n69 0.00463514
R144 VSS.n71 VSS.n1 0.00268919
R145 VSS.n68 VSS.n1 0.00244595
R146 VSS.n66 VSS 0.000932432
R147 VSS VSS.n74 0.000613314
R148 VDD.t3 VDD.t8 87.2098
R149 VDD.t6 VDD.t3 87.2098
R150 VDD.t5 VDD.t6 87.2098
R151 VDD.t2 VDD.t5 87.2098
R152 VDD.t1 VDD.t7 87.2098
R153 VDD.t7 VDD.t4 87.2098
R154 VDD.t4 VDD.t9 87.2098
R155 VDD.t9 VDD.t0 87.2098
R156 VDD.n0 VDD.t1 66.4976
R157 VDD.n0 VDD.t2 20.7127
R158 VDD VDD.n0 6.30057
R159 VCNTL.n0 VCNTL 9.51376
R160 VCNTL VCNTL.t0 7.11604
R161 VCNTL.n0 VCNTL.t1 2.35318
R162 VCNTL VCNTL.n0 0.000668776
C0 cap80p_mag_0.P a_47420_43837# 0.113f
C1 VDD a_45740_41735# 0.368f
C2 VSS a_46220_41735# 4.56e-19
C3 a_46220_41735# a_46700_41735# 0.0759f
C4 VDD cap80p_mag_0.P 0.208f
C5 a_47660_41735# a_47180_41735# 0.0754f
C6 VCNTL VDD 0.473f
C7 cap80p_mag_0.P a_45740_41735# 1.73e-19
C8 a_46460_43837# a_45980_43837# 0.0759f
C9 VDD a_47180_41735# 0.358f
C10 VCNTL a_45740_41735# 0.016f
C11 VDD a_45980_43837# 0.248f
C12 VSS VDD 0.0874f
C13 VDD a_46220_41735# 0.358f
C14 VDD a_46700_41735# 0.358f
C15 VCNTL cap80p_mag_0.P 0.113f
C16 VSS a_45740_41735# 0.00374f
C17 a_46220_41735# a_45740_41735# 0.0759f
C18 VDD a_47420_43837# 0.248f
C19 VSS cap80p_mag_0.P 0.295p
C20 VCNTL a_45980_43837# 0.0767f
C21 a_47420_43837# a_46940_43837# 0.0759f
C22 VDD a_47660_41735# 0.367f
C23 VSS VCNTL 4.18f
C24 VDD a_46460_43837# 0.248f
C25 a_46940_43837# a_46460_43837# 0.0759f
C26 VSS a_45980_43837# 0.00217f
C27 VDD a_46940_43837# 0.248f
C28 a_47180_41735# a_46700_41735# 0.0759f
C29 VSS VSUBS 0.176p
C30 VCNTL VSUBS 23.9f
C31 VDD VSUBS 22.7f
C32 cap80p_mag_0.P VSUBS 0.378p
C33 a_47660_41735# VSUBS 0.18f
C34 a_47420_43837# VSUBS 0.205f
C35 a_47180_41735# VSUBS 0.159f
C36 a_46940_43837# VSUBS 0.224f
C37 a_46700_41735# VSUBS 0.159f
C38 a_46460_43837# VSUBS 0.224f
C39 a_46220_41735# VSUBS 0.159f
C40 a_45980_43837# VSUBS 0.224f
C41 a_45740_41735# VSUBS 0.169f
C42 VCNTL.t0 VSUBS 3.45e-19
C43 VCNTL.t1 VSUBS 2.16f
C44 VCNTL.n0 VSUBS 1.94f
C45 VSS.t0 VSUBS 5.32f
C46 VSS.n0 VSUBS 0.0586f
C47 VSS.n1 VSUBS 0.00257f
C48 VSS.n2 VSUBS 0.044f
C49 VSS.t50 VSUBS 3.32f
C50 VSS.t42 VSUBS 3.03f
C51 VSS.n3 VSUBS 1.57f
C52 VSS.t13 VSUBS 3.03f
C53 VSS.n4 VSUBS 0.929f
C54 VSS.t64 VSUBS 3.03f
C55 VSS.n5 VSUBS 0.929f
C56 VSS.t29 VSUBS 3.03f
C57 VSS.n6 VSUBS 0.929f
C58 VSS.t33 VSUBS 3.03f
C59 VSS.n7 VSUBS 0.929f
C60 VSS.t57 VSUBS 3.03f
C61 VSS.n8 VSUBS 0.929f
C62 VSS.t5 VSUBS 3.03f
C63 VSS.n9 VSUBS 0.721f
C64 VSS.t43 VSUBS 3.32f
C65 VSS.t35 VSUBS 3.03f
C66 VSS.n10 VSUBS 1.57f
C67 VSS.t3 VSUBS 3.02f
C68 VSS.n11 VSUBS 0.929f
C69 VSS.t53 VSUBS 3.03f
C70 VSS.n12 VSUBS 0.929f
C71 VSS.t20 VSUBS 3.03f
C72 VSS.n13 VSUBS 0.929f
C73 VSS.t24 VSUBS 3.03f
C74 VSS.n14 VSUBS 0.929f
C75 VSS.t8 VSUBS 3.03f
C76 VSS.n15 VSUBS 0.929f
C77 VSS.t15 VSUBS 3.03f
C78 VSS.n16 VSUBS 0.721f
C79 VSS.t22 VSUBS 3.32f
C80 VSS.t11 VSUBS 3.03f
C81 VSS.n17 VSUBS 1.57f
C82 VSS.t47 VSUBS 3.02f
C83 VSS.n18 VSUBS 0.929f
C84 VSS.t39 VSUBS 3.03f
C85 VSS.n19 VSUBS 0.929f
C86 VSS.t56 VSUBS 3.03f
C87 VSS.n20 VSUBS 0.929f
C88 VSS.t61 VSUBS 3.03f
C89 VSS.n21 VSUBS 0.929f
C90 VSS.t31 VSUBS 3.03f
C91 VSS.n22 VSUBS 0.929f
C92 VSS.t38 VSUBS 3.03f
C93 VSS.n23 VSUBS 0.721f
C94 VSS.t49 VSUBS 3.32f
C95 VSS.t41 VSUBS 3.03f
C96 VSS.n24 VSUBS 1.57f
C97 VSS.t12 VSUBS 3.02f
C98 VSS.n25 VSUBS 0.929f
C99 VSS.t63 VSUBS 3.03f
C100 VSS.n26 VSUBS 0.929f
C101 VSS.t28 VSUBS 3.03f
C102 VSS.n27 VSUBS 0.929f
C103 VSS.t32 VSUBS 3.03f
C104 VSS.n28 VSUBS 0.929f
C105 VSS.t7 VSUBS 3.03f
C106 VSS.n29 VSUBS 0.929f
C107 VSS.t14 VSUBS 3.03f
C108 VSS.n30 VSUBS 1.22f
C109 VSS.n31 VSUBS 1.47f
C110 VSS.n32 VSUBS 1.21f
C111 VSS.n33 VSUBS 0.973f
C112 VSS.t48 VSUBS 3.32f
C113 VSS.t40 VSUBS 3.03f
C114 VSS.n34 VSUBS 1.57f
C115 VSS.t10 VSUBS 3.03f
C116 VSS.n35 VSUBS 0.929f
C117 VSS.t58 VSUBS 3.03f
C118 VSS.n36 VSUBS 0.929f
C119 VSS.t27 VSUBS 3.03f
C120 VSS.n37 VSUBS 0.929f
C121 VSS.t30 VSUBS 3.03f
C122 VSS.n38 VSUBS 0.929f
C123 VSS.t16 VSUBS 3.03f
C124 VSS.n39 VSUBS 0.929f
C125 VSS.t23 VSUBS 3.03f
C126 VSS.n40 VSUBS 0.721f
C127 VSS.t44 VSUBS 3.32f
C128 VSS.t36 VSUBS 3.03f
C129 VSS.n41 VSUBS 1.57f
C130 VSS.t4 VSUBS 3.03f
C131 VSS.n42 VSUBS 0.929f
C132 VSS.t54 VSUBS 3.03f
C133 VSS.n43 VSUBS 0.929f
C134 VSS.t21 VSUBS 3.03f
C135 VSS.n44 VSUBS 0.929f
C136 VSS.t25 VSUBS 3.03f
C137 VSS.n45 VSUBS 0.929f
C138 VSS.t60 VSUBS 3.03f
C139 VSS.n46 VSUBS 0.929f
C140 VSS.t6 VSUBS 3.03f
C141 VSS.n47 VSUBS 0.721f
C142 VSS.t26 VSUBS 3.32f
C143 VSS.t17 VSUBS 3.03f
C144 VSS.n48 VSUBS 1.57f
C145 VSS.t51 VSUBS 3.03f
C146 VSS.n49 VSUBS 0.929f
C147 VSS.t45 VSUBS 3.03f
C148 VSS.n50 VSUBS 0.929f
C149 VSS.t62 VSUBS 3.03f
C150 VSS.n51 VSUBS 0.929f
C151 VSS.t1 VSUBS 3.03f
C152 VSS.n52 VSUBS 0.929f
C153 VSS.t9 VSUBS 3.03f
C154 VSS.n53 VSUBS 0.929f
C155 VSS.t19 VSUBS 3.03f
C156 VSS.n54 VSUBS 0.721f
C157 VSS.t52 VSUBS 3.32f
C158 VSS.t46 VSUBS 3.03f
C159 VSS.n55 VSUBS 1.57f
C160 VSS.t18 VSUBS 3.03f
C161 VSS.n56 VSUBS 0.929f
C162 VSS.t2 VSUBS 3.03f
C163 VSS.n57 VSUBS 0.929f
C164 VSS.t34 VSUBS 3.03f
C165 VSS.n58 VSUBS 0.929f
C166 VSS.t37 VSUBS 3.03f
C167 VSS.n59 VSUBS 0.929f
C168 VSS.t55 VSUBS 3.03f
C169 VSS.n60 VSUBS 0.929f
C170 VSS.t59 VSUBS 3.03f
C171 VSS.n61 VSUBS 1.22f
C172 VSS.n62 VSUBS 1.47f
C173 VSS.n63 VSUBS 1.21f
C174 VSS.n64 VSUBS 0.971f
C175 VSS.n65 VSUBS 2.82f
C176 VSS.n66 VSUBS 1.79f
C177 VSS.n67 VSUBS 0.0536f
C178 VSS.n68 VSUBS 0.0175f
C179 VSS.n69 VSUBS 0.0233f
C180 VSS.n70 VSUBS 0.0245f
C181 VSS.n71 VSUBS 0.0189f
C182 VSS.n72 VSUBS 0.0482f
C183 VSS.n73 VSUBS 1.59f
C184 VSS.n74 VSUBS 4.55f
.ends

