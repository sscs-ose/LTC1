** sch_path: /home/shahid/GF180Projects/Top_test/Decoder_muxes/Xschem/2x1_mux_PEX_TB_ibr..sym
**.subckt 2x1_mux_PEX_TB_ibr.
V1 VDD VSS 3.3
.save i(v1)
V2 VSS GND 0
.save i(v2)
V4 S0 VSS pulse(3.3 0 0 100p 100p 350n 700n)
.save i(v4)
V6 I0 VSS pulse(0 3.3 0 100p 100p 200n 400n)3.3
.save i(v6)
V7 I1 VSS pulse(0 3.3 0 100p 100p 100n 200n)
.save i(v7)
x1 VSS S0 OUT I0 I1 VDD pex_mux_2x1_ibr
**** begin user architecture code

.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical



.include pex_mux_2x1_ibr.spice
.control
save all
tran 50p 800n
plot v(S0)  v(I0)+5 v(I1)+10 v(OUT)+15


*write test_nfet_03v3.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
