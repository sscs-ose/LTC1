magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2216 -2216 2416 2416
<< nwell >>
rect -216 -216 416 416
<< mvnsubdiff >>
rect -168 355 368 368
rect -168 309 -155 355
rect -109 309 -39 355
rect 7 309 77 355
rect 123 309 193 355
rect 239 309 309 355
rect 355 309 368 355
rect -168 296 368 309
rect -168 239 -96 296
rect -168 193 -155 239
rect -109 193 -96 239
rect 296 239 368 296
rect -168 123 -96 193
rect -168 77 -155 123
rect -109 77 -96 123
rect -168 7 -96 77
rect -168 -39 -155 7
rect -109 -39 -96 7
rect 296 193 309 239
rect 355 193 368 239
rect 296 123 368 193
rect 296 77 309 123
rect 355 77 368 123
rect 296 7 368 77
rect -168 -96 -96 -39
rect 296 -39 309 7
rect 355 -39 368 7
rect 296 -96 368 -39
rect -168 -109 368 -96
rect -168 -155 -155 -109
rect -109 -155 -39 -109
rect 7 -155 77 -109
rect 123 -155 193 -109
rect 239 -155 309 -109
rect 355 -155 368 -109
rect -168 -168 368 -155
<< mvnsubdiffcont >>
rect -155 309 -109 355
rect -39 309 7 355
rect 77 309 123 355
rect 193 309 239 355
rect 309 309 355 355
rect -155 193 -109 239
rect -155 77 -109 123
rect -155 -39 -109 7
rect 309 193 355 239
rect 309 77 355 123
rect 309 -39 355 7
rect -155 -155 -109 -109
rect -39 -155 7 -109
rect 77 -155 123 -109
rect 193 -155 239 -109
rect 309 -155 355 -109
<< mvpdiode >>
rect 0 187 200 200
rect 0 141 13 187
rect 59 141 141 187
rect 187 141 200 187
rect 0 59 200 141
rect 0 13 13 59
rect 59 13 141 59
rect 187 13 200 59
rect 0 0 200 13
<< mvpdiodec >>
rect 13 141 59 187
rect 141 141 187 187
rect 13 13 59 59
rect 141 13 187 59
<< metal1 >>
rect -168 355 368 368
rect -168 309 -155 355
rect -109 309 -39 355
rect 7 309 77 355
rect 123 309 193 355
rect 239 309 309 355
rect 355 309 368 355
rect -168 296 368 309
rect -168 239 -96 296
rect -168 193 -155 239
rect -109 193 -96 239
rect 296 239 368 296
rect -168 123 -96 193
rect -168 77 -155 123
rect -109 77 -96 123
rect -168 7 -96 77
rect -168 -39 -155 7
rect -109 -39 -96 7
rect 0 187 200 200
rect 0 141 13 187
rect 59 141 141 187
rect 187 141 200 187
rect 0 59 200 141
rect 0 13 13 59
rect 59 13 141 59
rect 187 13 200 59
rect 0 0 200 13
rect 296 193 309 239
rect 355 193 368 239
rect 296 123 368 193
rect 296 77 309 123
rect 355 77 368 123
rect 296 7 368 77
rect -168 -96 -96 -39
rect 296 -39 309 7
rect 355 -39 368 7
rect 296 -96 368 -39
rect -168 -109 368 -96
rect -168 -155 -155 -109
rect -109 -155 -39 -109
rect 7 -155 77 -109
rect 123 -155 193 -109
rect 239 -155 309 -109
rect 355 -155 368 -109
rect -168 -168 368 -155
<< labels >>
rlabel mvnsubdiffcont 100 -132 100 -132 4 MINUS
rlabel mvnsubdiffcont 100 332 100 332 4 MINUS
rlabel mvnsubdiffcont 332 100 332 100 4 MINUS
rlabel mvnsubdiffcont -132 100 -132 100 4 MINUS
rlabel metal1 100 100 100 100 4 PLUS
<< end >>
