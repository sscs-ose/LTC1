magic
tech gf180mcuC
magscale 1 10
timestamp 1693836168
<< psubdiff >>
rect 28514 10224 28561 10279
<< metal1 >>
rect 17927 14293 18154 14470
rect 17890 14268 18200 14293
rect 17890 14216 17931 14268
rect 17983 14216 18035 14268
rect 18087 14216 18139 14268
rect 18191 14216 18200 14268
rect 17890 14164 18200 14216
rect 17890 14112 17931 14164
rect 17983 14112 18035 14164
rect 18087 14112 18139 14164
rect 18191 14112 18200 14164
rect 17890 14060 18200 14112
rect 18742 14067 18894 14153
rect 19403 14109 19597 14176
rect 19390 14095 19702 14109
rect 17890 14008 17931 14060
rect 17983 14008 18035 14060
rect 18087 14008 18139 14060
rect 18191 14008 18200 14060
rect 17890 13943 18200 14008
rect 17890 13891 17919 13943
rect 17971 13891 18023 13943
rect 18075 13891 18127 13943
rect 18179 13891 18200 13943
rect 17890 13839 18200 13891
rect 17890 13787 17919 13839
rect 17971 13787 18023 13839
rect 18075 13787 18127 13839
rect 18179 13787 18200 13839
rect 17890 13735 18200 13787
rect 17890 13683 17919 13735
rect 17971 13683 18023 13735
rect 18075 13683 18127 13735
rect 18179 13683 18200 13735
rect 17890 13631 18200 13683
rect 17890 13579 17919 13631
rect 17971 13579 18023 13631
rect 18075 13579 18127 13631
rect 18179 13579 18200 13631
rect 17890 13527 18200 13579
rect 17890 13475 17919 13527
rect 17971 13475 18023 13527
rect 18075 13475 18127 13527
rect 18179 13475 18200 13527
rect 17890 13423 18200 13475
rect 17890 13371 17919 13423
rect 17971 13371 18023 13423
rect 18075 13371 18127 13423
rect 18179 13371 18200 13423
rect 17890 13319 18200 13371
rect 17890 13267 17919 13319
rect 17971 13267 18023 13319
rect 18075 13267 18127 13319
rect 18179 13267 18200 13319
rect 17890 13215 18200 13267
rect 17890 13163 17919 13215
rect 17971 13163 18023 13215
rect 18075 13163 18127 13215
rect 18179 13163 18200 13215
rect 18712 14013 18924 14067
rect 18712 13961 18736 14013
rect 18788 13961 18840 14013
rect 18892 13961 18924 14013
rect 18712 13909 18924 13961
rect 18712 13857 18736 13909
rect 18788 13857 18840 13909
rect 18892 13857 18924 13909
rect 18712 13805 18924 13857
rect 18712 13753 18736 13805
rect 18788 13753 18840 13805
rect 18892 13753 18924 13805
rect 18712 13701 18924 13753
rect 18712 13649 18736 13701
rect 18788 13649 18840 13701
rect 18892 13649 18924 13701
rect 18712 13597 18924 13649
rect 18712 13545 18736 13597
rect 18788 13545 18840 13597
rect 18892 13545 18924 13597
rect 18712 13493 18924 13545
rect 18712 13441 18736 13493
rect 18788 13441 18840 13493
rect 18892 13441 18924 13493
rect 18712 13389 18924 13441
rect 18712 13337 18736 13389
rect 18788 13337 18840 13389
rect 18892 13337 18924 13389
rect 18712 13285 18924 13337
rect 18712 13233 18736 13285
rect 18788 13233 18840 13285
rect 18892 13233 18924 13285
rect 18712 13212 18924 13233
rect 19367 14057 19702 14095
rect 22087 14087 23144 14135
rect 19367 14005 19390 14057
rect 19442 14005 19494 14057
rect 19546 14005 19598 14057
rect 19650 14005 19702 14057
rect 19367 13953 19702 14005
rect 19367 13901 19390 13953
rect 19442 13901 19494 13953
rect 19546 13901 19598 13953
rect 19650 13901 19702 13953
rect 21918 13926 22114 14087
rect 22275 14086 22915 14087
rect 22275 13927 22497 14086
rect 22656 13927 22915 14086
rect 22275 13926 22915 13927
rect 23076 13926 23144 14087
rect 22087 13904 23144 13926
rect 28009 13917 45862 14382
rect 19367 13849 19702 13901
rect 19367 13797 19390 13849
rect 19442 13797 19494 13849
rect 19546 13797 19598 13849
rect 19650 13797 19702 13849
rect 19367 13745 19702 13797
rect 19367 13693 19390 13745
rect 19442 13693 19494 13745
rect 19546 13693 19598 13745
rect 19650 13693 19702 13745
rect 19367 13641 19702 13693
rect 19367 13589 19390 13641
rect 19442 13589 19494 13641
rect 19546 13589 19598 13641
rect 19650 13589 19702 13641
rect 19367 13537 19702 13589
rect 19367 13485 19390 13537
rect 19442 13485 19494 13537
rect 19546 13485 19598 13537
rect 19650 13485 19702 13537
rect 21938 13528 22849 13570
rect 19367 13433 19702 13485
rect 19367 13381 19390 13433
rect 19442 13381 19494 13433
rect 19546 13381 19598 13433
rect 19650 13381 19702 13433
rect 21833 13392 21964 13528
rect 22100 13527 22678 13528
rect 22100 13393 22388 13527
rect 22522 13393 22678 13527
rect 22100 13392 22678 13393
rect 22814 13392 22849 13528
rect 19367 13329 19702 13381
rect 21938 13367 22849 13392
rect 19367 13277 19390 13329
rect 19442 13277 19494 13329
rect 19546 13277 19598 13329
rect 19650 13277 19702 13329
rect 19367 13225 19702 13277
rect 17890 13111 18200 13163
rect 19367 13173 19390 13225
rect 19442 13173 19494 13225
rect 19546 13173 19598 13225
rect 19650 13173 19702 13225
rect 19367 13155 19656 13173
rect 17890 13059 17919 13111
rect 17971 13059 18023 13111
rect 18075 13059 18127 13111
rect 18179 13059 18200 13111
rect 17890 13028 18200 13059
rect 21781 13104 22530 13132
rect 21781 13002 21813 13104
rect 21915 13103 22385 13104
rect 21915 13003 22053 13103
rect 22153 13003 22385 13103
rect 21915 13002 22385 13003
rect 22487 13002 22530 13104
rect 21781 12982 22530 13002
rect 28009 12882 28474 13917
rect 29503 13648 30444 13693
rect 29388 13471 29511 13648
rect 29688 13647 30247 13648
rect 29688 13472 29857 13647
rect 30032 13472 30247 13647
rect 29688 13471 30247 13472
rect 30424 13471 30444 13648
rect 29503 13439 30444 13471
rect 25831 12651 30284 12882
rect 18916 12491 24077 12615
rect 25831 12525 30285 12651
rect 19381 12486 19601 12491
rect 22275 12489 24077 12491
rect 22275 12487 23800 12489
rect 22275 12486 23246 12487
rect 18770 11989 18860 12015
rect 18770 11928 18788 11989
rect 18849 11928 18860 11989
rect 22410 11980 22490 12486
rect 22823 12412 22947 12486
rect 23122 12412 23246 12486
rect 23406 12412 23530 12487
rect 23676 12412 23800 12487
rect 23953 12412 24077 12489
rect 25830 12504 30285 12525
rect 25830 12503 30284 12504
rect 24624 12412 24967 12413
rect 25540 12412 25770 12413
rect 25830 12412 26744 12503
rect 22793 12410 26744 12412
rect 22793 11960 26566 12410
rect 18770 11853 18860 11928
rect 18770 11790 18787 11853
rect 18850 11790 18860 11853
rect 18770 11721 18860 11790
rect 19772 11835 19858 11845
rect 19772 11762 19795 11835
rect 19849 11762 19858 11835
rect 18770 11720 18949 11721
rect 18770 11659 18788 11720
rect 18849 11659 18949 11720
rect 18770 11658 18949 11659
rect 18770 11647 18860 11658
rect 19772 11620 19858 11762
rect 22312 11238 22390 11860
rect 26630 11857 26747 11897
rect 26630 11794 26657 11857
rect 26720 11794 26747 11857
rect 26630 11738 26747 11794
rect 26630 11737 26774 11738
rect 26630 11676 26657 11737
rect 26718 11676 26774 11737
rect 26630 11675 26774 11676
rect 26630 11664 26747 11675
rect 30430 11557 30771 11566
rect 30430 11556 30577 11557
rect 30430 11504 30442 11556
rect 30494 11505 30577 11556
rect 30629 11543 30771 11557
rect 30629 11505 30703 11543
rect 30494 11504 30703 11505
rect 30430 11491 30703 11504
rect 30755 11491 30771 11543
rect 30430 11455 30771 11491
rect 30430 11448 30663 11455
rect 30430 11396 30443 11448
rect 30495 11447 30663 11448
rect 30495 11396 30560 11447
rect 30430 11395 30560 11396
rect 30612 11395 30663 11447
rect 30430 11381 30663 11395
rect 30861 11355 31027 13592
rect 31886 11708 32351 13917
rect 33469 13170 34585 13216
rect 33327 12964 33480 13170
rect 33686 13169 34367 13170
rect 33686 12965 33963 13169
rect 34167 12965 34367 13169
rect 33686 12964 34367 12965
rect 34573 12964 34585 13170
rect 44097 13128 44562 13917
rect 45397 13128 45862 13917
rect 47868 13160 52184 13374
rect 33469 12930 34585 12964
rect 41677 12670 41885 12734
rect 41677 12547 41720 12670
rect 41843 12547 41885 12670
rect 41677 12421 41885 12547
rect 41677 12296 41719 12421
rect 41844 12296 41885 12421
rect 41677 12214 41885 12296
rect 41677 12196 42058 12214
rect 41677 12073 41720 12196
rect 41843 12073 42058 12196
rect 41677 12061 42058 12073
rect 30796 11319 31027 11355
rect 30796 11251 31001 11319
rect 22312 11079 22783 11238
rect 30893 11205 31001 11251
rect 30893 11146 30909 11205
rect 30894 11133 30909 11146
rect 30981 11133 31001 11205
rect 22312 10710 22390 11079
rect 30894 11056 31001 11133
rect 30894 10986 30903 11056
rect 30973 10986 31001 11056
rect 30894 10967 31001 10986
rect 19749 10620 19858 10644
rect 19749 10563 19768 10620
rect 19838 10563 19858 10620
rect 19749 10408 19858 10563
rect 22383 10516 22415 10522
rect 16721 10041 19619 10338
rect 29638 10333 30181 10361
rect 27356 10322 28991 10329
rect 29062 10322 29497 10329
rect 27356 10300 29497 10322
rect 27356 10209 29617 10300
rect 27356 10203 29480 10209
rect 29638 10181 29655 10333
rect 29807 10332 30181 10333
rect 29807 10182 30014 10332
rect 30164 10182 30181 10332
rect 29807 10181 30181 10182
rect 29638 10167 30181 10181
rect 16721 4908 17018 10041
rect 19780 9902 19892 10120
rect 30649 10018 31431 10169
rect 22320 9505 22424 9707
rect 22320 9472 22743 9505
rect 22320 9390 22985 9472
rect 22320 9358 22743 9390
rect 18785 8751 18894 8764
rect 18785 8690 18809 8751
rect 18870 8750 18894 8751
rect 18870 8690 18955 8750
rect 18785 8687 18955 8690
rect 18785 8637 18894 8687
rect 18785 8574 18808 8637
rect 18871 8574 18894 8637
rect 18785 8517 18894 8574
rect 19791 8646 19863 8717
rect 19791 8573 19803 8646
rect 19857 8573 19863 8646
rect 19791 8558 19863 8573
rect 22320 8553 22424 9358
rect 30649 9096 30800 10018
rect 30898 9879 31296 9909
rect 30898 9875 31077 9879
rect 30898 9823 30905 9875
rect 30957 9827 31077 9875
rect 31129 9827 31296 9879
rect 30957 9823 31296 9827
rect 30898 9803 31296 9823
rect 33817 9606 34300 9721
rect 34174 9565 34300 9606
rect 34174 9541 34877 9565
rect 34174 9540 34455 9541
rect 34174 9427 34184 9540
rect 34297 9427 34455 9540
rect 34174 9426 34455 9427
rect 34570 9540 34877 9541
rect 34570 9427 34743 9540
rect 34856 9427 34877 9540
rect 34570 9426 34877 9427
rect 34174 9411 34877 9426
rect 34566 9410 34877 9411
rect 31950 9211 32102 9410
rect 31203 9198 32130 9211
rect 31203 9197 31614 9198
rect 30530 8898 31075 9096
rect 31203 9047 31221 9197
rect 31371 9047 31614 9197
rect 31203 9046 31614 9047
rect 31766 9197 32130 9198
rect 31766 9047 31951 9197
rect 32101 9047 32130 9197
rect 31766 9046 32130 9047
rect 31203 9030 32130 9046
rect 26726 8764 26927 8827
rect 26726 8737 26844 8764
rect 26726 8676 26752 8737
rect 26813 8676 26844 8737
rect 26726 8621 26844 8676
rect 18785 8456 18809 8517
rect 18870 8456 18894 8517
rect 18785 8424 18894 8456
rect 26351 8450 26561 8578
rect 26726 8558 26751 8621
rect 26814 8558 26844 8621
rect 26726 8535 26844 8558
rect 22865 7922 22989 8384
rect 23323 7922 23447 8384
rect 24418 7922 24542 8396
rect 25281 7922 25405 8393
rect 25975 7922 26099 8413
rect 26224 8326 26561 8450
rect 26343 8324 26561 8326
rect 26351 7922 26561 8324
rect 22340 7916 26561 7922
rect 30436 7916 30437 7921
rect 22340 7798 30444 7916
rect 26351 7706 30444 7798
rect 17724 6842 18965 6957
rect 17619 6679 17758 6842
rect 17921 6841 18758 6842
rect 17921 6680 18215 6841
rect 18376 6680 18758 6841
rect 17921 6679 18758 6680
rect 18921 6679 18965 6842
rect 22085 6822 22546 6850
rect 21988 6705 22102 6822
rect 22219 6821 22546 6822
rect 22219 6706 22399 6821
rect 22514 6706 22546 6821
rect 22219 6705 22546 6706
rect 22085 6683 22546 6705
rect 17724 6618 18965 6679
rect 18925 6328 19703 6349
rect 18855 6194 18960 6328
rect 19094 6327 19554 6328
rect 19094 6195 19250 6327
rect 19382 6195 19554 6327
rect 19094 6194 19554 6195
rect 19688 6194 19703 6328
rect 18925 6169 19703 6194
rect 27190 5845 27445 7706
rect 30849 6635 31075 8898
rect 27177 5817 27780 5845
rect 27177 5816 27596 5817
rect 27177 5658 27194 5816
rect 27352 5658 27596 5816
rect 27177 5657 27596 5658
rect 27756 5657 27780 5817
rect 27177 5568 27780 5657
rect 27177 5408 27211 5568
rect 27371 5567 27780 5568
rect 27371 5409 27597 5567
rect 27755 5409 27780 5567
rect 27371 5408 27780 5409
rect 27177 5392 27780 5408
rect 32225 5373 32329 5795
rect 33295 5113 33729 9309
rect 47868 8256 48082 13160
rect 47615 8242 48082 8256
rect 47615 8241 47935 8242
rect 47615 8163 47780 8241
rect 47858 8163 47935 8241
rect 47615 8162 47935 8163
rect 48015 8162 48082 8242
rect 47615 8150 48082 8162
rect 43227 7112 43321 7123
rect 46171 7119 46241 7209
rect 46432 7119 46521 7206
rect 46706 7119 46795 7208
rect 46908 7119 46997 7216
rect 43227 7111 43449 7112
rect 43820 7111 43992 7112
rect 43227 6941 43278 7111
rect 43448 6941 43821 7111
rect 43991 7110 44714 7111
rect 43991 6942 44532 7110
rect 44700 6942 44714 7110
rect 46136 7091 47059 7119
rect 46136 7086 46925 7091
rect 46136 7008 46183 7086
rect 46259 7083 46925 7086
rect 46259 7081 46709 7083
rect 46259 7008 46429 7081
rect 46136 7003 46429 7008
rect 46505 7005 46709 7081
rect 46785 7013 46925 7083
rect 47001 7013 47059 7091
rect 46785 7005 47059 7013
rect 46505 7003 47059 7005
rect 46136 6961 47059 7003
rect 43991 6941 44714 6942
rect 43227 6940 43449 6941
rect 43820 6940 43992 6941
rect 43227 6919 43321 6940
rect 43759 6087 44718 6127
rect 43759 6009 43813 6087
rect 43889 6074 44718 6087
rect 43889 6009 44062 6074
rect 43759 5996 44062 6009
rect 44138 6073 44718 6074
rect 44138 6069 44518 6073
rect 44138 5996 44296 6069
rect 43759 5991 44296 5996
rect 44372 5995 44518 6069
rect 44594 5995 44718 6073
rect 44372 5991 44718 5995
rect 43759 5971 44718 5991
rect 40140 4953 42232 5122
rect 16721 4611 24352 4908
rect 30400 4524 30604 4659
rect 27094 4444 27485 4463
rect 27094 4443 27342 4444
rect 27094 4315 27111 4443
rect 27239 4315 27342 4443
rect 27094 4314 27342 4315
rect 27472 4314 27485 4444
rect 27094 4248 27485 4314
rect 30400 4399 30434 4524
rect 30559 4399 30604 4524
rect 30400 4263 30604 4399
rect 27094 4118 27107 4248
rect 27237 4247 27485 4248
rect 27237 4119 27343 4247
rect 27471 4119 27485 4247
rect 30300 4262 30604 4263
rect 30300 4139 30435 4262
rect 30558 4139 30604 4262
rect 42800 4230 42910 4490
rect 43290 4210 43400 4470
rect 30300 4138 30604 4139
rect 30400 4129 30604 4138
rect 27237 4118 27485 4119
rect 27094 4108 27485 4118
rect 27110 3940 27240 4108
rect 44729 2789 45104 4670
rect 48134 1877 48214 2325
rect 47978 1179 48050 1247
rect 47970 1164 48050 1179
rect 47978 864 48050 1164
rect 47432 -795 54511 -568
<< via1 >>
rect 17931 14216 17983 14268
rect 18035 14216 18087 14268
rect 18139 14216 18191 14268
rect 17931 14112 17983 14164
rect 18035 14112 18087 14164
rect 18139 14112 18191 14164
rect 17931 14008 17983 14060
rect 18035 14008 18087 14060
rect 18139 14008 18191 14060
rect 17919 13891 17971 13943
rect 18023 13891 18075 13943
rect 18127 13891 18179 13943
rect 17919 13787 17971 13839
rect 18023 13787 18075 13839
rect 18127 13787 18179 13839
rect 17919 13683 17971 13735
rect 18023 13683 18075 13735
rect 18127 13683 18179 13735
rect 17919 13579 17971 13631
rect 18023 13579 18075 13631
rect 18127 13579 18179 13631
rect 17919 13475 17971 13527
rect 18023 13475 18075 13527
rect 18127 13475 18179 13527
rect 17919 13371 17971 13423
rect 18023 13371 18075 13423
rect 18127 13371 18179 13423
rect 17919 13267 17971 13319
rect 18023 13267 18075 13319
rect 18127 13267 18179 13319
rect 17919 13163 17971 13215
rect 18023 13163 18075 13215
rect 18127 13163 18179 13215
rect 18736 13961 18788 14013
rect 18840 13961 18892 14013
rect 18736 13857 18788 13909
rect 18840 13857 18892 13909
rect 18736 13753 18788 13805
rect 18840 13753 18892 13805
rect 18736 13649 18788 13701
rect 18840 13649 18892 13701
rect 18736 13545 18788 13597
rect 18840 13545 18892 13597
rect 18736 13441 18788 13493
rect 18840 13441 18892 13493
rect 18736 13337 18788 13389
rect 18840 13337 18892 13389
rect 18736 13233 18788 13285
rect 18840 13233 18892 13285
rect 19390 14005 19442 14057
rect 19494 14005 19546 14057
rect 19598 14005 19650 14057
rect 19390 13901 19442 13953
rect 19494 13901 19546 13953
rect 19598 13901 19650 13953
rect 22114 13926 22275 14087
rect 22497 13927 22656 14086
rect 22915 13926 23076 14087
rect 19390 13797 19442 13849
rect 19494 13797 19546 13849
rect 19598 13797 19650 13849
rect 19390 13693 19442 13745
rect 19494 13693 19546 13745
rect 19598 13693 19650 13745
rect 19390 13589 19442 13641
rect 19494 13589 19546 13641
rect 19598 13589 19650 13641
rect 19390 13485 19442 13537
rect 19494 13485 19546 13537
rect 19598 13485 19650 13537
rect 19390 13381 19442 13433
rect 19494 13381 19546 13433
rect 19598 13381 19650 13433
rect 21964 13392 22100 13528
rect 22388 13393 22522 13527
rect 22678 13392 22814 13528
rect 19390 13277 19442 13329
rect 19494 13277 19546 13329
rect 19598 13277 19650 13329
rect 19390 13173 19442 13225
rect 19494 13173 19546 13225
rect 19598 13173 19650 13225
rect 17919 13059 17971 13111
rect 18023 13059 18075 13111
rect 18127 13059 18179 13111
rect 21813 13002 21915 13104
rect 22053 13003 22153 13103
rect 22385 13002 22487 13104
rect 29511 13471 29688 13648
rect 29857 13472 30032 13647
rect 30247 13471 30424 13648
rect 18788 11928 18849 11989
rect 18787 11790 18850 11853
rect 19795 11762 19849 11835
rect 18788 11659 18849 11720
rect 26657 11794 26720 11857
rect 26657 11676 26718 11737
rect 30442 11504 30494 11556
rect 30577 11505 30629 11557
rect 30703 11491 30755 11543
rect 30443 11396 30495 11448
rect 30560 11395 30612 11447
rect 33480 12964 33686 13170
rect 33963 12965 34167 13169
rect 34367 12964 34573 13170
rect 41720 12547 41843 12670
rect 41719 12296 41844 12421
rect 41720 12073 41843 12196
rect 30909 11133 30981 11205
rect 30903 10986 30973 11056
rect 19768 10563 19838 10620
rect 29655 10181 29807 10333
rect 30014 10182 30164 10332
rect 18809 8690 18870 8751
rect 18808 8574 18871 8637
rect 19803 8573 19857 8646
rect 30905 9823 30957 9875
rect 31077 9827 31129 9879
rect 34184 9427 34297 9540
rect 34455 9426 34570 9541
rect 34743 9427 34856 9540
rect 31221 9047 31371 9197
rect 31614 9046 31766 9198
rect 31951 9047 32101 9197
rect 26752 8676 26813 8737
rect 18809 8456 18870 8517
rect 26751 8558 26814 8621
rect 17758 6679 17921 6842
rect 18215 6680 18376 6841
rect 18758 6679 18921 6842
rect 22102 6705 22219 6822
rect 22399 6706 22514 6821
rect 18960 6194 19094 6328
rect 19250 6195 19382 6327
rect 19554 6194 19688 6328
rect 27194 5658 27352 5816
rect 27596 5657 27756 5817
rect 27211 5408 27371 5568
rect 27597 5409 27755 5567
rect 47780 8163 47858 8241
rect 47935 8162 48015 8242
rect 43278 6941 43448 7111
rect 43821 6941 43991 7111
rect 44532 6942 44700 7110
rect 46183 7008 46259 7086
rect 46429 7003 46505 7081
rect 46709 7005 46785 7083
rect 46925 7013 47001 7091
rect 43813 6009 43889 6087
rect 44062 5996 44138 6074
rect 44296 5991 44372 6069
rect 44518 5995 44594 6073
rect 27111 4315 27239 4443
rect 27342 4314 27472 4444
rect 30434 4399 30559 4524
rect 27107 4118 27237 4248
rect 27343 4119 27471 4247
rect 30435 4139 30558 4262
<< metal2 >>
rect 41677 16508 44499 16716
rect 17890 14268 18200 14293
rect 17890 14216 17931 14268
rect 17983 14216 18035 14268
rect 18087 14216 18139 14268
rect 18191 14216 18200 14268
rect 17890 14164 18200 14216
rect 17890 14112 17931 14164
rect 17983 14112 18035 14164
rect 18087 14112 18139 14164
rect 18191 14112 18200 14164
rect 17890 14060 18200 14112
rect 19390 14095 19702 14109
rect 17890 14008 17931 14060
rect 17983 14008 18035 14060
rect 18087 14008 18139 14060
rect 18191 14008 18200 14060
rect 17890 13943 18200 14008
rect 17890 13891 17919 13943
rect 17971 13891 18023 13943
rect 18075 13891 18127 13943
rect 18179 13891 18200 13943
rect 17890 13839 18200 13891
rect 17890 13787 17919 13839
rect 17971 13787 18023 13839
rect 18075 13787 18127 13839
rect 18179 13787 18200 13839
rect 17890 13735 18200 13787
rect 17890 13683 17919 13735
rect 17971 13683 18023 13735
rect 18075 13683 18127 13735
rect 18179 13683 18200 13735
rect 17890 13631 18200 13683
rect 17890 13579 17919 13631
rect 17971 13579 18023 13631
rect 18075 13579 18127 13631
rect 18179 13579 18200 13631
rect 17890 13527 18200 13579
rect 17890 13475 17919 13527
rect 17971 13475 18023 13527
rect 18075 13475 18127 13527
rect 18179 13475 18200 13527
rect 17890 13423 18200 13475
rect 17890 13371 17919 13423
rect 17971 13371 18023 13423
rect 18075 13371 18127 13423
rect 18179 13371 18200 13423
rect 17890 13319 18200 13371
rect 17890 13267 17919 13319
rect 17971 13267 18023 13319
rect 18075 13267 18127 13319
rect 18179 13267 18200 13319
rect 17890 13215 18200 13267
rect 17890 13163 17919 13215
rect 17971 13163 18023 13215
rect 18075 13163 18127 13215
rect 18179 13163 18200 13215
rect 18712 14013 18924 14067
rect 18712 13961 18736 14013
rect 18788 13961 18840 14013
rect 18892 13961 18924 14013
rect 18712 13909 18924 13961
rect 18712 13857 18736 13909
rect 18788 13857 18840 13909
rect 18892 13857 18924 13909
rect 18712 13805 18924 13857
rect 18712 13753 18736 13805
rect 18788 13753 18840 13805
rect 18892 13753 18924 13805
rect 18712 13701 18924 13753
rect 18712 13649 18736 13701
rect 18788 13649 18840 13701
rect 18892 13649 18924 13701
rect 18712 13597 18924 13649
rect 18712 13545 18736 13597
rect 18788 13545 18840 13597
rect 18892 13545 18924 13597
rect 18712 13493 18924 13545
rect 18712 13441 18736 13493
rect 18788 13441 18840 13493
rect 18892 13441 18924 13493
rect 18712 13389 18924 13441
rect 18712 13337 18736 13389
rect 18788 13337 18840 13389
rect 18892 13337 18924 13389
rect 18712 13285 18924 13337
rect 18712 13233 18736 13285
rect 18788 13233 18840 13285
rect 18892 13233 18924 13285
rect 18712 13212 18924 13233
rect 19367 14057 19702 14095
rect 19367 14005 19390 14057
rect 19442 14005 19494 14057
rect 19546 14005 19598 14057
rect 19650 14005 19702 14057
rect 19367 13953 19702 14005
rect 19367 13901 19390 13953
rect 19442 13901 19494 13953
rect 19546 13901 19598 13953
rect 19650 13901 19702 13953
rect 22087 14087 23144 14135
rect 26184 14087 27185 14111
rect 22087 13926 22114 14087
rect 22275 14086 22915 14087
rect 22275 13927 22497 14086
rect 22656 13927 22915 14086
rect 22275 13926 22915 13927
rect 23076 13926 26211 14087
rect 26372 13926 26578 14087
rect 26739 13926 26997 14087
rect 27158 13926 27185 14087
rect 22087 13904 23144 13926
rect 19367 13849 19702 13901
rect 26184 13889 27185 13926
rect 19367 13797 19390 13849
rect 19442 13797 19494 13849
rect 19546 13797 19598 13849
rect 19650 13797 19702 13849
rect 19367 13745 19702 13797
rect 19367 13693 19390 13745
rect 19442 13693 19494 13745
rect 19546 13693 19598 13745
rect 19650 13693 19702 13745
rect 19367 13641 19702 13693
rect 29503 13648 30444 13693
rect 19367 13589 19390 13641
rect 19442 13589 19494 13641
rect 19546 13589 19598 13641
rect 19650 13589 19702 13641
rect 19367 13537 19702 13589
rect 19367 13485 19390 13537
rect 19442 13485 19494 13537
rect 19546 13485 19598 13537
rect 19650 13485 19702 13537
rect 19367 13433 19702 13485
rect 19367 13381 19390 13433
rect 19442 13381 19494 13433
rect 19546 13381 19598 13433
rect 19650 13381 19702 13433
rect 19367 13329 19702 13381
rect 21938 13528 22849 13570
rect 25430 13528 26138 13541
rect 21938 13392 21964 13528
rect 22100 13527 22678 13528
rect 22100 13393 22388 13527
rect 22522 13393 22678 13527
rect 22100 13392 22678 13393
rect 22814 13512 26138 13528
rect 22814 13408 25496 13512
rect 25600 13408 25684 13512
rect 25788 13408 25879 13512
rect 25983 13408 26138 13512
rect 29502 13471 29511 13648
rect 29688 13647 30247 13648
rect 29688 13472 29857 13647
rect 30032 13472 30247 13647
rect 29688 13471 30247 13472
rect 30424 13471 30444 13648
rect 29503 13439 30444 13471
rect 22814 13392 26138 13408
rect 21938 13367 22849 13392
rect 25430 13374 26138 13392
rect 25430 13373 26015 13374
rect 19367 13277 19390 13329
rect 19442 13277 19494 13329
rect 19546 13277 19598 13329
rect 19650 13277 19702 13329
rect 19367 13225 19702 13277
rect 17890 13111 18200 13163
rect 17890 13059 17919 13111
rect 17971 13059 18023 13111
rect 18075 13059 18127 13111
rect 18179 13059 18200 13111
rect 17890 13028 18200 13059
rect 17927 10567 18154 13028
rect 18742 11989 18894 13212
rect 19367 13173 19390 13225
rect 19442 13173 19494 13225
rect 19546 13173 19598 13225
rect 19650 13173 19702 13225
rect 30247 13313 30424 13439
rect 19367 13155 19656 13173
rect 19403 12673 19597 13155
rect 30247 13136 30786 13313
rect 21799 13104 22548 13132
rect 21799 13002 21813 13104
rect 21915 13103 22385 13104
rect 21915 13003 22053 13103
rect 22153 13003 22385 13103
rect 21915 13002 22385 13003
rect 22487 13002 25242 13104
rect 21799 12982 22548 13002
rect 18742 11942 18788 11989
rect 18741 11928 18788 11942
rect 18849 11928 18894 11989
rect 18741 11853 18894 11928
rect 18741 11790 18787 11853
rect 18850 11790 18894 11853
rect 18741 11720 18894 11790
rect 18741 11659 18788 11720
rect 18849 11659 18894 11720
rect 18741 11646 18894 11659
rect 19460 11721 19597 12673
rect 25140 12604 25242 13002
rect 25140 12502 26739 12604
rect 26637 11906 26739 12502
rect 26630 11857 26747 11906
rect 19772 11835 19858 11845
rect 19772 11762 19795 11835
rect 19849 11762 19858 11835
rect 19772 11721 19858 11762
rect 19460 11620 19858 11721
rect 26630 11794 26657 11857
rect 26720 11794 26747 11857
rect 26630 11737 26747 11794
rect 26630 11676 26657 11737
rect 26718 11676 26747 11737
rect 26630 11673 26747 11676
rect 27323 11637 27684 11723
rect 19460 11573 19597 11620
rect 27323 11613 27409 11637
rect 26556 11527 27409 11613
rect 30609 11564 30786 13136
rect 33469 13170 34585 13216
rect 33469 12964 33480 13170
rect 33686 13169 34367 13170
rect 33686 12965 33963 13169
rect 34167 12965 34367 13169
rect 33686 12964 34367 12965
rect 34573 12964 34585 13170
rect 33469 12930 34585 12964
rect 30433 11557 30786 11564
rect 30433 11556 30577 11557
rect 30433 11504 30442 11556
rect 30494 11505 30577 11556
rect 30629 11543 30786 11557
rect 30629 11505 30703 11543
rect 30494 11504 30703 11505
rect 30433 11491 30703 11504
rect 30755 11491 30786 11543
rect 30433 11448 30786 11491
rect 30433 11396 30443 11448
rect 30495 11447 30786 11448
rect 30495 11396 30560 11447
rect 30433 11395 30560 11396
rect 30612 11395 30786 11447
rect 30433 11387 30786 11395
rect 19749 10629 19858 10644
rect 19749 10620 19860 10629
rect 19749 10567 19768 10620
rect 17927 10563 19768 10567
rect 19838 10567 19860 10620
rect 19838 10563 19866 10567
rect 17927 10340 19866 10563
rect 26981 10494 27288 10523
rect 26981 10493 27122 10494
rect 26981 10433 26998 10493
rect 27058 10434 27122 10493
rect 27182 10434 27288 10494
rect 27058 10433 27288 10434
rect 26981 10417 27288 10433
rect 29638 10333 30181 10361
rect 28991 10280 29059 10289
rect 28987 10263 29059 10280
rect 28891 10157 29059 10263
rect 29638 10181 29655 10333
rect 29807 10181 30013 10333
rect 30165 10181 30181 10333
rect 29638 10167 30181 10181
rect 27209 10052 27449 10088
rect 27209 10051 27358 10052
rect 27209 9991 27234 10051
rect 27294 9992 27358 10051
rect 27418 9992 27449 10052
rect 27294 9991 27449 9992
rect 27209 9965 27449 9991
rect 30609 9936 30786 11387
rect 30894 11340 31001 11353
rect 30894 11268 31103 11340
rect 30894 11205 31001 11268
rect 30894 11133 30909 11205
rect 30981 11133 31001 11205
rect 30894 11056 31001 11133
rect 30894 10986 30903 11056
rect 30973 10986 31001 11056
rect 30894 10967 31001 10986
rect 34367 9963 34573 12930
rect 41677 12670 41885 16508
rect 41677 12547 41720 12670
rect 41843 12547 41885 12670
rect 41677 12421 41885 12547
rect 41677 12296 41719 12421
rect 41844 12296 41885 12421
rect 41677 12214 41885 12296
rect 41677 12196 42058 12214
rect 41677 12073 41720 12196
rect 41843 12073 42058 12196
rect 41677 12061 42058 12073
rect 30609 9909 31266 9936
rect 34201 9932 34573 9963
rect 30609 9879 31296 9909
rect 30609 9875 31077 9879
rect 30609 9823 30905 9875
rect 30957 9827 31077 9875
rect 31129 9827 31296 9879
rect 30957 9823 31296 9827
rect 30609 9803 31296 9823
rect 30609 9759 31266 9803
rect 33725 9795 34573 9932
rect 33725 9789 34200 9795
rect 34055 9721 34212 9724
rect 33817 9715 34212 9721
rect 33764 9698 34212 9715
rect 33764 9606 34213 9698
rect 33764 9605 33840 9606
rect 34036 9581 34213 9606
rect 34036 9541 48092 9581
rect 34036 9540 34455 9541
rect 34036 9427 34184 9540
rect 34297 9427 34455 9540
rect 34036 9426 34455 9427
rect 34570 9540 48092 9541
rect 34570 9427 34743 9540
rect 34856 9427 48092 9540
rect 34570 9426 48092 9427
rect 34036 9386 48092 9426
rect 31203 9198 32130 9211
rect 31203 9046 31220 9198
rect 31372 9046 31614 9198
rect 31766 9046 31950 9198
rect 32102 9046 32130 9198
rect 31203 9030 32130 9046
rect 26597 8889 27507 9025
rect 27371 8886 27507 8889
rect 19554 8788 19688 8804
rect 19788 8788 19865 8844
rect 18757 8751 18921 8769
rect 18757 8690 18809 8751
rect 18870 8690 18921 8751
rect 18757 8637 18921 8690
rect 18757 8574 18808 8637
rect 18871 8574 18921 8637
rect 18757 8517 18921 8574
rect 18757 8456 18809 8517
rect 18870 8456 18921 8517
rect 18757 8298 18921 8456
rect 18758 6957 18921 8298
rect 19554 8719 19865 8788
rect 26726 8737 26844 8827
rect 27371 8750 27837 8886
rect 19554 8687 19863 8719
rect 17724 6842 18965 6957
rect 17724 6679 17758 6842
rect 17921 6841 18758 6842
rect 17921 6680 18215 6841
rect 18376 6680 18758 6841
rect 17921 6679 18758 6680
rect 18921 6679 18965 6842
rect 17724 6618 18965 6679
rect 19554 6349 19688 8687
rect 19788 8646 19863 8687
rect 19788 8573 19803 8646
rect 19857 8573 19863 8646
rect 19788 8558 19863 8573
rect 26726 8676 26752 8737
rect 26813 8676 26844 8737
rect 26726 8621 26844 8676
rect 26726 8558 26751 8621
rect 26814 8558 26844 8621
rect 47897 8560 48092 9386
rect 26726 8535 26844 8558
rect 26726 8425 26843 8535
rect 26684 6907 26884 8425
rect 47867 8256 48122 8560
rect 47615 8242 48122 8256
rect 47615 8241 47935 8242
rect 47615 8163 47780 8241
rect 47858 8163 47935 8241
rect 47615 8162 47935 8163
rect 48015 8162 48122 8242
rect 47615 8150 48122 8162
rect 44110 7124 44460 7130
rect 43227 7111 44715 7124
rect 43227 6941 43278 7111
rect 43448 6941 43821 7111
rect 43991 6941 44531 7111
rect 44701 6941 44715 7111
rect 46136 7091 47059 7119
rect 46136 7086 46925 7091
rect 46136 7008 46183 7086
rect 46259 7083 46925 7086
rect 46259 7081 46709 7083
rect 46259 7008 46429 7081
rect 46136 7003 46429 7008
rect 46505 7005 46709 7081
rect 46785 7013 46925 7083
rect 47001 7013 47059 7091
rect 46785 7005 47059 7013
rect 46505 7003 47059 7005
rect 46136 6961 47059 7003
rect 43227 6919 44715 6941
rect 22083 6822 26884 6907
rect 22083 6707 22102 6822
rect 22085 6705 22102 6707
rect 22219 6821 26884 6822
rect 22219 6706 22399 6821
rect 22514 6707 26884 6821
rect 44110 6850 44480 6919
rect 44110 6810 44460 6850
rect 22514 6706 26843 6707
rect 22219 6705 26843 6706
rect 22085 6683 22546 6705
rect 18925 6328 19703 6349
rect 18925 6194 18960 6328
rect 19094 6327 19554 6328
rect 19094 6195 19250 6327
rect 19382 6195 19554 6327
rect 19094 6194 19554 6195
rect 19688 6194 19703 6328
rect 18925 6169 19703 6194
rect 43759 6087 44718 6127
rect 43759 6009 43813 6087
rect 43889 6074 44718 6087
rect 43889 6009 44062 6074
rect 43759 5996 44062 6009
rect 44138 6073 44718 6074
rect 44138 6069 44518 6073
rect 44138 5996 44296 6069
rect 43759 5991 44296 5996
rect 44372 5995 44518 6069
rect 44594 5995 44718 6073
rect 44372 5991 44718 5995
rect 43759 5971 44718 5991
rect 27177 5817 27780 5845
rect 27177 5657 27193 5817
rect 27353 5657 27596 5817
rect 27756 5657 27780 5817
rect 27177 5568 27780 5657
rect 27177 5408 27211 5568
rect 27371 5408 27596 5568
rect 27756 5408 27780 5568
rect 27177 5392 27780 5408
rect 30400 4524 30604 4659
rect 47867 4534 48122 8150
rect 27094 4444 27485 4463
rect 27094 4314 27110 4444
rect 27240 4314 27342 4444
rect 27472 4314 27485 4444
rect 27094 4248 27485 4314
rect 27094 4118 27107 4248
rect 27237 4118 27342 4248
rect 27472 4118 27485 4248
rect 30400 4399 30434 4524
rect 30559 4399 30604 4524
rect 30400 4263 30604 4399
rect 46238 4279 48122 4534
rect 30400 4138 30434 4263
rect 30559 4138 30604 4263
rect 30400 4129 30604 4138
rect 27094 4108 27485 4118
<< via2 >>
rect 26211 13926 26372 14087
rect 26578 13926 26739 14087
rect 26997 13926 27158 14087
rect 25496 13408 25600 13512
rect 25684 13408 25788 13512
rect 25879 13408 25983 13512
rect 26998 10433 27058 10493
rect 27122 10434 27182 10494
rect 29655 10181 29807 10333
rect 30013 10332 30165 10333
rect 30013 10182 30014 10332
rect 30014 10182 30164 10332
rect 30164 10182 30165 10332
rect 30013 10181 30165 10182
rect 27234 9991 27294 10051
rect 27358 9992 27418 10052
rect 31220 9197 31372 9198
rect 31220 9047 31221 9197
rect 31221 9047 31371 9197
rect 31371 9047 31372 9197
rect 31220 9046 31372 9047
rect 31614 9046 31766 9198
rect 31950 9197 32102 9198
rect 31950 9047 31951 9197
rect 31951 9047 32101 9197
rect 32101 9047 32102 9197
rect 31950 9046 32102 9047
rect 43278 6941 43448 7111
rect 43821 6941 43991 7111
rect 44531 7110 44701 7111
rect 44531 6942 44532 7110
rect 44532 6942 44700 7110
rect 44700 6942 44701 7110
rect 44531 6941 44701 6942
rect 46183 7008 46259 7086
rect 46429 7003 46505 7081
rect 46709 7005 46785 7083
rect 46925 7013 47001 7091
rect 43813 6009 43889 6087
rect 44062 5996 44138 6074
rect 44296 5991 44372 6069
rect 44518 5995 44594 6073
rect 27193 5816 27353 5817
rect 27193 5658 27194 5816
rect 27194 5658 27352 5816
rect 27352 5658 27353 5816
rect 27193 5657 27353 5658
rect 27596 5657 27756 5817
rect 27211 5408 27371 5568
rect 27596 5567 27756 5568
rect 27596 5409 27597 5567
rect 27597 5409 27755 5567
rect 27755 5409 27756 5567
rect 27596 5408 27756 5409
rect 27110 4443 27240 4444
rect 27110 4315 27111 4443
rect 27111 4315 27239 4443
rect 27239 4315 27240 4443
rect 27110 4314 27240 4315
rect 27342 4314 27472 4444
rect 27107 4118 27237 4248
rect 27342 4247 27472 4248
rect 27342 4119 27343 4247
rect 27343 4119 27471 4247
rect 27471 4119 27472 4247
rect 27342 4118 27472 4119
rect 30434 4399 30559 4524
rect 30434 4262 30559 4263
rect 30434 4139 30435 4262
rect 30435 4139 30558 4262
rect 30558 4139 30559 4262
rect 30434 4138 30559 4139
<< metal3 >>
rect 26184 14087 27185 14111
rect 26184 13926 26211 14087
rect 26372 13926 26578 14087
rect 26739 13926 26997 14087
rect 27158 13926 27185 14087
rect 26184 13889 27185 13926
rect 26035 13541 26139 13542
rect 25430 13512 26139 13541
rect 25430 13408 25496 13512
rect 25600 13408 25684 13512
rect 25788 13408 25879 13512
rect 25983 13408 26139 13512
rect 25430 13373 26139 13408
rect 26035 10281 26139 13373
rect 26992 12944 27163 13889
rect 27022 10510 27132 12944
rect 26983 10494 27202 10510
rect 26983 10493 27122 10494
rect 26983 10433 26998 10493
rect 27058 10434 27122 10493
rect 27182 10434 27202 10494
rect 27058 10433 27202 10434
rect 26983 10417 27202 10433
rect 29638 10333 30181 10361
rect 26035 10177 27374 10281
rect 27258 10068 27374 10177
rect 29638 10181 29655 10333
rect 29807 10181 30013 10333
rect 30165 10181 30600 10333
rect 29638 10167 30181 10181
rect 27219 10052 27438 10068
rect 27219 10051 27358 10052
rect 27219 9991 27234 10051
rect 27294 9992 27358 10051
rect 27418 9992 27438 10052
rect 27294 9991 27438 9992
rect 27219 9975 27438 9991
rect 30448 9198 30600 10181
rect 31203 9198 32130 9211
rect 30448 9046 31220 9198
rect 31372 9046 31614 9198
rect 31766 9046 31950 9198
rect 32102 9046 32130 9198
rect 31203 9030 32130 9046
rect 30400 7124 43272 7125
rect 44110 7124 44460 7130
rect 30400 7111 44715 7124
rect 30400 6941 43278 7111
rect 43448 6941 43821 7111
rect 43991 6941 44531 7111
rect 44701 6941 44715 7111
rect 46136 7091 47059 7119
rect 46136 7086 46925 7091
rect 46136 7008 46183 7086
rect 46259 7083 46925 7086
rect 46259 7081 46709 7083
rect 46259 7008 46429 7081
rect 46136 7003 46429 7008
rect 46505 7005 46709 7081
rect 46785 7013 46925 7083
rect 47001 7013 47059 7091
rect 46785 7005 47059 7013
rect 46505 7003 47059 7005
rect 46136 6961 47059 7003
rect 30400 6919 44715 6941
rect 27177 5817 27780 5845
rect 27177 5657 27193 5817
rect 27353 5657 27596 5817
rect 27756 5657 27780 5817
rect 27177 5568 27780 5657
rect 27177 5408 27211 5568
rect 27371 5408 27596 5568
rect 27756 5408 27780 5568
rect 27177 5392 27780 5408
rect 27211 4463 27371 5392
rect 30400 4524 30606 6919
rect 44110 6850 44480 6919
rect 44110 6810 44460 6850
rect 46593 6130 46752 6961
rect 43759 6087 46752 6130
rect 43759 6009 43813 6087
rect 43889 6074 46752 6087
rect 43889 6009 44062 6074
rect 43759 5996 44062 6009
rect 44138 6073 46752 6074
rect 44138 6069 44518 6073
rect 44138 5996 44296 6069
rect 43759 5991 44296 5996
rect 44372 5995 44518 6069
rect 44594 5995 46752 6073
rect 44372 5991 46752 5995
rect 43759 5971 46752 5991
rect 27094 4444 27485 4463
rect 27094 4314 27110 4444
rect 27240 4314 27342 4444
rect 27472 4314 27485 4444
rect 27094 4248 27485 4314
rect 27094 4118 27107 4248
rect 27237 4118 27342 4248
rect 27472 4118 27485 4248
rect 30400 4399 30434 4524
rect 30559 4399 30606 4524
rect 30400 4263 30606 4399
rect 30400 4138 30434 4263
rect 30559 4138 30606 4263
rect 30400 4129 30606 4138
rect 27094 4108 27485 4118
<< metal5 >>
rect 94588 92926 98134 93436
rect 97358 483 98134 92926
rect 67761 -293 98134 483
use A_MUX  A_MUX_0 ~/GF180Projects/Layout/Magic/VCO1/A_MUx
timestamp 1693500185
transform 1 0 42495 0 1 4782
box -285 -452 3979 2227
use cap_11p  cap_11p_0 ~/GF180Projects/Layout/Magic/ATIF/CP
timestamp 1693309357
transform 1 0 74717 0 1 12873
box -26450 -13708 -6739 632
use cap_240p  cap_240p_0 ~/GF180Projects/Layout/Magic/ATIF/CP
timestamp 1693315383
transform 1 0 89584 0 -1 24489
box -68140 -68970 6839 8429
use CP_1  CP_1_0 ~/GF180Projects/Layout/Magic/ATIF/CP
timestamp 1691774029
transform 1 0 32106 0 1 10461
box -1319 -1188 2101 1378
use mux_magic  mux_magic_0 ~/GF180Projects/Layout/Magic/ATIF/mux_magic
timestamp 1693836065
transform 1 0 28348 0 1 11078
box -1637 -890 2187 1549
use mux_magic  mux_magic_1
timestamp 1693836065
transform 1 0 28501 0 -1 9424
box -1637 -890 2187 1549
use mux_magic  mux_magic_2
timestamp 1693836065
transform 1 0 20523 0 1 11061
box -1637 -890 2187 1549
use mux_magic  mux_magic_3
timestamp 1693836065
transform 1 0 20529 0 -1 9347
box -1637 -890 2187 1549
use PFD_T2  PFD_T2_0 ~/GF180Projects/Layout/Magic/ATIF/PFD_2
timestamp 1693469249
transform 1 0 22661 0 1 8437
box -28 -113 4062 3793
use RES_74k  RES_74k_1 ~/GF180Projects/Layout/Magic/ATIF/Res/RES_p
timestamp 1692794530
transform -1 0 51462 0 -1 12102
box 3672 -1094 9598 4966
use VCO_DFF_C  VCO_DFF_C_0 ~/GF180Projects/Layout/Magic/VCO1/VCO_DFF_C
timestamp 1693141881
transform 1 0 24282 0 1 -1600
box 0 -27 23932 7170
<< labels >>
flabel metal1 30954 13379 30954 13379 0 FreeSans 1280 0 0 0 ITAIL
port 14 nsew
flabel metal1 21788 13047 21788 13047 0 FreeSans 1600 0 0 0 S2
port 20 nsew
flabel metal1 22036 6756 22036 6756 0 FreeSans 1600 0 0 0 S3
port 19 nsew
flabel metal1 18804 14117 18804 14117 0 FreeSans 1600 0 0 0 S1
port 23 nsew
flabel metal1 17670 6747 17670 6747 0 FreeSans 1600 0 0 0 S6
port 24 nsew
flabel metal1 21995 13993 21995 13993 0 FreeSans 1600 0 0 0 UP_INPUT
port 25 nsew
flabel metal1 21858 13460 21858 13460 0 FreeSans 1600 0 0 0 DN_INPUT
port 26 nsew
flabel metal1 19504 14129 19504 14129 0 FreeSans 800 0 0 0 PRE_SCALAR
port 28 nsew
flabel metal1 18022 14399 18022 14399 0 FreeSans 1600 0 0 0 F_IN
port 29 nsew
flabel metal1 18872 6250 18872 6250 0 FreeSans 1600 0 0 0 DIV_OUT
port 30 nsew
flabel metal1 29437 13558 29437 13558 0 FreeSans 1600 0 0 0 UP
port 31 nsew
flabel metal1 30955 6730 30955 6730 0 FreeSans 1600 0 0 0 DN
port 32 nsew
flabel metal1 33398 13080 33398 13080 0 FreeSans 1600 0 0 0 ITAIL1
port 33 nsew
flabel metal1 48168 1912 48168 1912 0 FreeSans 1600 0 0 0 OUTB
port 37 nsew
flabel metal1 48004 888 48004 888 0 FreeSans 1600 0 0 0 OUT
port 38 nsew
flabel metal1 32279 5743 32279 5743 0 FreeSans 1600 0 0 0 VCTRL2
port 39 nsew
flabel metal1 33470 8331 33470 8331 0 FreeSans 1600 0 0 0 VSS
port 40 nsew
flabel metal1 30024 14122 30024 14122 0 FreeSans 1600 0 0 0 VDD
port 41 nsew
flabel metal1 42870 4240 42870 4240 0 FreeSans 1600 0 0 0 VCTRL_IN
port 42 nsew
flabel metal1 43370 4280 43370 4280 0 FreeSans 1600 0 0 0 S4
port 43 nsew
<< end >>
