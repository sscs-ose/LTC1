magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1453 -1732 1453 1732
<< metal2 >>
rect -453 727 453 732
rect -453 699 -448 727
rect -420 699 -386 727
rect -358 699 -324 727
rect -296 699 -262 727
rect -234 699 -200 727
rect -172 699 -138 727
rect -110 699 -76 727
rect -48 699 -14 727
rect 14 699 48 727
rect 76 699 110 727
rect 138 699 172 727
rect 200 699 234 727
rect 262 699 296 727
rect 324 699 358 727
rect 386 699 420 727
rect 448 699 453 727
rect -453 665 453 699
rect -453 637 -448 665
rect -420 637 -386 665
rect -358 637 -324 665
rect -296 637 -262 665
rect -234 637 -200 665
rect -172 637 -138 665
rect -110 637 -76 665
rect -48 637 -14 665
rect 14 637 48 665
rect 76 637 110 665
rect 138 637 172 665
rect 200 637 234 665
rect 262 637 296 665
rect 324 637 358 665
rect 386 637 420 665
rect 448 637 453 665
rect -453 603 453 637
rect -453 575 -448 603
rect -420 575 -386 603
rect -358 575 -324 603
rect -296 575 -262 603
rect -234 575 -200 603
rect -172 575 -138 603
rect -110 575 -76 603
rect -48 575 -14 603
rect 14 575 48 603
rect 76 575 110 603
rect 138 575 172 603
rect 200 575 234 603
rect 262 575 296 603
rect 324 575 358 603
rect 386 575 420 603
rect 448 575 453 603
rect -453 541 453 575
rect -453 513 -448 541
rect -420 513 -386 541
rect -358 513 -324 541
rect -296 513 -262 541
rect -234 513 -200 541
rect -172 513 -138 541
rect -110 513 -76 541
rect -48 513 -14 541
rect 14 513 48 541
rect 76 513 110 541
rect 138 513 172 541
rect 200 513 234 541
rect 262 513 296 541
rect 324 513 358 541
rect 386 513 420 541
rect 448 513 453 541
rect -453 479 453 513
rect -453 451 -448 479
rect -420 451 -386 479
rect -358 451 -324 479
rect -296 451 -262 479
rect -234 451 -200 479
rect -172 451 -138 479
rect -110 451 -76 479
rect -48 451 -14 479
rect 14 451 48 479
rect 76 451 110 479
rect 138 451 172 479
rect 200 451 234 479
rect 262 451 296 479
rect 324 451 358 479
rect 386 451 420 479
rect 448 451 453 479
rect -453 417 453 451
rect -453 389 -448 417
rect -420 389 -386 417
rect -358 389 -324 417
rect -296 389 -262 417
rect -234 389 -200 417
rect -172 389 -138 417
rect -110 389 -76 417
rect -48 389 -14 417
rect 14 389 48 417
rect 76 389 110 417
rect 138 389 172 417
rect 200 389 234 417
rect 262 389 296 417
rect 324 389 358 417
rect 386 389 420 417
rect 448 389 453 417
rect -453 355 453 389
rect -453 327 -448 355
rect -420 327 -386 355
rect -358 327 -324 355
rect -296 327 -262 355
rect -234 327 -200 355
rect -172 327 -138 355
rect -110 327 -76 355
rect -48 327 -14 355
rect 14 327 48 355
rect 76 327 110 355
rect 138 327 172 355
rect 200 327 234 355
rect 262 327 296 355
rect 324 327 358 355
rect 386 327 420 355
rect 448 327 453 355
rect -453 293 453 327
rect -453 265 -448 293
rect -420 265 -386 293
rect -358 265 -324 293
rect -296 265 -262 293
rect -234 265 -200 293
rect -172 265 -138 293
rect -110 265 -76 293
rect -48 265 -14 293
rect 14 265 48 293
rect 76 265 110 293
rect 138 265 172 293
rect 200 265 234 293
rect 262 265 296 293
rect 324 265 358 293
rect 386 265 420 293
rect 448 265 453 293
rect -453 231 453 265
rect -453 203 -448 231
rect -420 203 -386 231
rect -358 203 -324 231
rect -296 203 -262 231
rect -234 203 -200 231
rect -172 203 -138 231
rect -110 203 -76 231
rect -48 203 -14 231
rect 14 203 48 231
rect 76 203 110 231
rect 138 203 172 231
rect 200 203 234 231
rect 262 203 296 231
rect 324 203 358 231
rect 386 203 420 231
rect 448 203 453 231
rect -453 169 453 203
rect -453 141 -448 169
rect -420 141 -386 169
rect -358 141 -324 169
rect -296 141 -262 169
rect -234 141 -200 169
rect -172 141 -138 169
rect -110 141 -76 169
rect -48 141 -14 169
rect 14 141 48 169
rect 76 141 110 169
rect 138 141 172 169
rect 200 141 234 169
rect 262 141 296 169
rect 324 141 358 169
rect 386 141 420 169
rect 448 141 453 169
rect -453 107 453 141
rect -453 79 -448 107
rect -420 79 -386 107
rect -358 79 -324 107
rect -296 79 -262 107
rect -234 79 -200 107
rect -172 79 -138 107
rect -110 79 -76 107
rect -48 79 -14 107
rect 14 79 48 107
rect 76 79 110 107
rect 138 79 172 107
rect 200 79 234 107
rect 262 79 296 107
rect 324 79 358 107
rect 386 79 420 107
rect 448 79 453 107
rect -453 45 453 79
rect -453 17 -448 45
rect -420 17 -386 45
rect -358 17 -324 45
rect -296 17 -262 45
rect -234 17 -200 45
rect -172 17 -138 45
rect -110 17 -76 45
rect -48 17 -14 45
rect 14 17 48 45
rect 76 17 110 45
rect 138 17 172 45
rect 200 17 234 45
rect 262 17 296 45
rect 324 17 358 45
rect 386 17 420 45
rect 448 17 453 45
rect -453 -17 453 17
rect -453 -45 -448 -17
rect -420 -45 -386 -17
rect -358 -45 -324 -17
rect -296 -45 -262 -17
rect -234 -45 -200 -17
rect -172 -45 -138 -17
rect -110 -45 -76 -17
rect -48 -45 -14 -17
rect 14 -45 48 -17
rect 76 -45 110 -17
rect 138 -45 172 -17
rect 200 -45 234 -17
rect 262 -45 296 -17
rect 324 -45 358 -17
rect 386 -45 420 -17
rect 448 -45 453 -17
rect -453 -79 453 -45
rect -453 -107 -448 -79
rect -420 -107 -386 -79
rect -358 -107 -324 -79
rect -296 -107 -262 -79
rect -234 -107 -200 -79
rect -172 -107 -138 -79
rect -110 -107 -76 -79
rect -48 -107 -14 -79
rect 14 -107 48 -79
rect 76 -107 110 -79
rect 138 -107 172 -79
rect 200 -107 234 -79
rect 262 -107 296 -79
rect 324 -107 358 -79
rect 386 -107 420 -79
rect 448 -107 453 -79
rect -453 -141 453 -107
rect -453 -169 -448 -141
rect -420 -169 -386 -141
rect -358 -169 -324 -141
rect -296 -169 -262 -141
rect -234 -169 -200 -141
rect -172 -169 -138 -141
rect -110 -169 -76 -141
rect -48 -169 -14 -141
rect 14 -169 48 -141
rect 76 -169 110 -141
rect 138 -169 172 -141
rect 200 -169 234 -141
rect 262 -169 296 -141
rect 324 -169 358 -141
rect 386 -169 420 -141
rect 448 -169 453 -141
rect -453 -203 453 -169
rect -453 -231 -448 -203
rect -420 -231 -386 -203
rect -358 -231 -324 -203
rect -296 -231 -262 -203
rect -234 -231 -200 -203
rect -172 -231 -138 -203
rect -110 -231 -76 -203
rect -48 -231 -14 -203
rect 14 -231 48 -203
rect 76 -231 110 -203
rect 138 -231 172 -203
rect 200 -231 234 -203
rect 262 -231 296 -203
rect 324 -231 358 -203
rect 386 -231 420 -203
rect 448 -231 453 -203
rect -453 -265 453 -231
rect -453 -293 -448 -265
rect -420 -293 -386 -265
rect -358 -293 -324 -265
rect -296 -293 -262 -265
rect -234 -293 -200 -265
rect -172 -293 -138 -265
rect -110 -293 -76 -265
rect -48 -293 -14 -265
rect 14 -293 48 -265
rect 76 -293 110 -265
rect 138 -293 172 -265
rect 200 -293 234 -265
rect 262 -293 296 -265
rect 324 -293 358 -265
rect 386 -293 420 -265
rect 448 -293 453 -265
rect -453 -327 453 -293
rect -453 -355 -448 -327
rect -420 -355 -386 -327
rect -358 -355 -324 -327
rect -296 -355 -262 -327
rect -234 -355 -200 -327
rect -172 -355 -138 -327
rect -110 -355 -76 -327
rect -48 -355 -14 -327
rect 14 -355 48 -327
rect 76 -355 110 -327
rect 138 -355 172 -327
rect 200 -355 234 -327
rect 262 -355 296 -327
rect 324 -355 358 -327
rect 386 -355 420 -327
rect 448 -355 453 -327
rect -453 -389 453 -355
rect -453 -417 -448 -389
rect -420 -417 -386 -389
rect -358 -417 -324 -389
rect -296 -417 -262 -389
rect -234 -417 -200 -389
rect -172 -417 -138 -389
rect -110 -417 -76 -389
rect -48 -417 -14 -389
rect 14 -417 48 -389
rect 76 -417 110 -389
rect 138 -417 172 -389
rect 200 -417 234 -389
rect 262 -417 296 -389
rect 324 -417 358 -389
rect 386 -417 420 -389
rect 448 -417 453 -389
rect -453 -451 453 -417
rect -453 -479 -448 -451
rect -420 -479 -386 -451
rect -358 -479 -324 -451
rect -296 -479 -262 -451
rect -234 -479 -200 -451
rect -172 -479 -138 -451
rect -110 -479 -76 -451
rect -48 -479 -14 -451
rect 14 -479 48 -451
rect 76 -479 110 -451
rect 138 -479 172 -451
rect 200 -479 234 -451
rect 262 -479 296 -451
rect 324 -479 358 -451
rect 386 -479 420 -451
rect 448 -479 453 -451
rect -453 -513 453 -479
rect -453 -541 -448 -513
rect -420 -541 -386 -513
rect -358 -541 -324 -513
rect -296 -541 -262 -513
rect -234 -541 -200 -513
rect -172 -541 -138 -513
rect -110 -541 -76 -513
rect -48 -541 -14 -513
rect 14 -541 48 -513
rect 76 -541 110 -513
rect 138 -541 172 -513
rect 200 -541 234 -513
rect 262 -541 296 -513
rect 324 -541 358 -513
rect 386 -541 420 -513
rect 448 -541 453 -513
rect -453 -575 453 -541
rect -453 -603 -448 -575
rect -420 -603 -386 -575
rect -358 -603 -324 -575
rect -296 -603 -262 -575
rect -234 -603 -200 -575
rect -172 -603 -138 -575
rect -110 -603 -76 -575
rect -48 -603 -14 -575
rect 14 -603 48 -575
rect 76 -603 110 -575
rect 138 -603 172 -575
rect 200 -603 234 -575
rect 262 -603 296 -575
rect 324 -603 358 -575
rect 386 -603 420 -575
rect 448 -603 453 -575
rect -453 -637 453 -603
rect -453 -665 -448 -637
rect -420 -665 -386 -637
rect -358 -665 -324 -637
rect -296 -665 -262 -637
rect -234 -665 -200 -637
rect -172 -665 -138 -637
rect -110 -665 -76 -637
rect -48 -665 -14 -637
rect 14 -665 48 -637
rect 76 -665 110 -637
rect 138 -665 172 -637
rect 200 -665 234 -637
rect 262 -665 296 -637
rect 324 -665 358 -637
rect 386 -665 420 -637
rect 448 -665 453 -637
rect -453 -699 453 -665
rect -453 -727 -448 -699
rect -420 -727 -386 -699
rect -358 -727 -324 -699
rect -296 -727 -262 -699
rect -234 -727 -200 -699
rect -172 -727 -138 -699
rect -110 -727 -76 -699
rect -48 -727 -14 -699
rect 14 -727 48 -699
rect 76 -727 110 -699
rect 138 -727 172 -699
rect 200 -727 234 -699
rect 262 -727 296 -699
rect 324 -727 358 -699
rect 386 -727 420 -699
rect 448 -727 453 -699
rect -453 -732 453 -727
<< via2 >>
rect -448 699 -420 727
rect -386 699 -358 727
rect -324 699 -296 727
rect -262 699 -234 727
rect -200 699 -172 727
rect -138 699 -110 727
rect -76 699 -48 727
rect -14 699 14 727
rect 48 699 76 727
rect 110 699 138 727
rect 172 699 200 727
rect 234 699 262 727
rect 296 699 324 727
rect 358 699 386 727
rect 420 699 448 727
rect -448 637 -420 665
rect -386 637 -358 665
rect -324 637 -296 665
rect -262 637 -234 665
rect -200 637 -172 665
rect -138 637 -110 665
rect -76 637 -48 665
rect -14 637 14 665
rect 48 637 76 665
rect 110 637 138 665
rect 172 637 200 665
rect 234 637 262 665
rect 296 637 324 665
rect 358 637 386 665
rect 420 637 448 665
rect -448 575 -420 603
rect -386 575 -358 603
rect -324 575 -296 603
rect -262 575 -234 603
rect -200 575 -172 603
rect -138 575 -110 603
rect -76 575 -48 603
rect -14 575 14 603
rect 48 575 76 603
rect 110 575 138 603
rect 172 575 200 603
rect 234 575 262 603
rect 296 575 324 603
rect 358 575 386 603
rect 420 575 448 603
rect -448 513 -420 541
rect -386 513 -358 541
rect -324 513 -296 541
rect -262 513 -234 541
rect -200 513 -172 541
rect -138 513 -110 541
rect -76 513 -48 541
rect -14 513 14 541
rect 48 513 76 541
rect 110 513 138 541
rect 172 513 200 541
rect 234 513 262 541
rect 296 513 324 541
rect 358 513 386 541
rect 420 513 448 541
rect -448 451 -420 479
rect -386 451 -358 479
rect -324 451 -296 479
rect -262 451 -234 479
rect -200 451 -172 479
rect -138 451 -110 479
rect -76 451 -48 479
rect -14 451 14 479
rect 48 451 76 479
rect 110 451 138 479
rect 172 451 200 479
rect 234 451 262 479
rect 296 451 324 479
rect 358 451 386 479
rect 420 451 448 479
rect -448 389 -420 417
rect -386 389 -358 417
rect -324 389 -296 417
rect -262 389 -234 417
rect -200 389 -172 417
rect -138 389 -110 417
rect -76 389 -48 417
rect -14 389 14 417
rect 48 389 76 417
rect 110 389 138 417
rect 172 389 200 417
rect 234 389 262 417
rect 296 389 324 417
rect 358 389 386 417
rect 420 389 448 417
rect -448 327 -420 355
rect -386 327 -358 355
rect -324 327 -296 355
rect -262 327 -234 355
rect -200 327 -172 355
rect -138 327 -110 355
rect -76 327 -48 355
rect -14 327 14 355
rect 48 327 76 355
rect 110 327 138 355
rect 172 327 200 355
rect 234 327 262 355
rect 296 327 324 355
rect 358 327 386 355
rect 420 327 448 355
rect -448 265 -420 293
rect -386 265 -358 293
rect -324 265 -296 293
rect -262 265 -234 293
rect -200 265 -172 293
rect -138 265 -110 293
rect -76 265 -48 293
rect -14 265 14 293
rect 48 265 76 293
rect 110 265 138 293
rect 172 265 200 293
rect 234 265 262 293
rect 296 265 324 293
rect 358 265 386 293
rect 420 265 448 293
rect -448 203 -420 231
rect -386 203 -358 231
rect -324 203 -296 231
rect -262 203 -234 231
rect -200 203 -172 231
rect -138 203 -110 231
rect -76 203 -48 231
rect -14 203 14 231
rect 48 203 76 231
rect 110 203 138 231
rect 172 203 200 231
rect 234 203 262 231
rect 296 203 324 231
rect 358 203 386 231
rect 420 203 448 231
rect -448 141 -420 169
rect -386 141 -358 169
rect -324 141 -296 169
rect -262 141 -234 169
rect -200 141 -172 169
rect -138 141 -110 169
rect -76 141 -48 169
rect -14 141 14 169
rect 48 141 76 169
rect 110 141 138 169
rect 172 141 200 169
rect 234 141 262 169
rect 296 141 324 169
rect 358 141 386 169
rect 420 141 448 169
rect -448 79 -420 107
rect -386 79 -358 107
rect -324 79 -296 107
rect -262 79 -234 107
rect -200 79 -172 107
rect -138 79 -110 107
rect -76 79 -48 107
rect -14 79 14 107
rect 48 79 76 107
rect 110 79 138 107
rect 172 79 200 107
rect 234 79 262 107
rect 296 79 324 107
rect 358 79 386 107
rect 420 79 448 107
rect -448 17 -420 45
rect -386 17 -358 45
rect -324 17 -296 45
rect -262 17 -234 45
rect -200 17 -172 45
rect -138 17 -110 45
rect -76 17 -48 45
rect -14 17 14 45
rect 48 17 76 45
rect 110 17 138 45
rect 172 17 200 45
rect 234 17 262 45
rect 296 17 324 45
rect 358 17 386 45
rect 420 17 448 45
rect -448 -45 -420 -17
rect -386 -45 -358 -17
rect -324 -45 -296 -17
rect -262 -45 -234 -17
rect -200 -45 -172 -17
rect -138 -45 -110 -17
rect -76 -45 -48 -17
rect -14 -45 14 -17
rect 48 -45 76 -17
rect 110 -45 138 -17
rect 172 -45 200 -17
rect 234 -45 262 -17
rect 296 -45 324 -17
rect 358 -45 386 -17
rect 420 -45 448 -17
rect -448 -107 -420 -79
rect -386 -107 -358 -79
rect -324 -107 -296 -79
rect -262 -107 -234 -79
rect -200 -107 -172 -79
rect -138 -107 -110 -79
rect -76 -107 -48 -79
rect -14 -107 14 -79
rect 48 -107 76 -79
rect 110 -107 138 -79
rect 172 -107 200 -79
rect 234 -107 262 -79
rect 296 -107 324 -79
rect 358 -107 386 -79
rect 420 -107 448 -79
rect -448 -169 -420 -141
rect -386 -169 -358 -141
rect -324 -169 -296 -141
rect -262 -169 -234 -141
rect -200 -169 -172 -141
rect -138 -169 -110 -141
rect -76 -169 -48 -141
rect -14 -169 14 -141
rect 48 -169 76 -141
rect 110 -169 138 -141
rect 172 -169 200 -141
rect 234 -169 262 -141
rect 296 -169 324 -141
rect 358 -169 386 -141
rect 420 -169 448 -141
rect -448 -231 -420 -203
rect -386 -231 -358 -203
rect -324 -231 -296 -203
rect -262 -231 -234 -203
rect -200 -231 -172 -203
rect -138 -231 -110 -203
rect -76 -231 -48 -203
rect -14 -231 14 -203
rect 48 -231 76 -203
rect 110 -231 138 -203
rect 172 -231 200 -203
rect 234 -231 262 -203
rect 296 -231 324 -203
rect 358 -231 386 -203
rect 420 -231 448 -203
rect -448 -293 -420 -265
rect -386 -293 -358 -265
rect -324 -293 -296 -265
rect -262 -293 -234 -265
rect -200 -293 -172 -265
rect -138 -293 -110 -265
rect -76 -293 -48 -265
rect -14 -293 14 -265
rect 48 -293 76 -265
rect 110 -293 138 -265
rect 172 -293 200 -265
rect 234 -293 262 -265
rect 296 -293 324 -265
rect 358 -293 386 -265
rect 420 -293 448 -265
rect -448 -355 -420 -327
rect -386 -355 -358 -327
rect -324 -355 -296 -327
rect -262 -355 -234 -327
rect -200 -355 -172 -327
rect -138 -355 -110 -327
rect -76 -355 -48 -327
rect -14 -355 14 -327
rect 48 -355 76 -327
rect 110 -355 138 -327
rect 172 -355 200 -327
rect 234 -355 262 -327
rect 296 -355 324 -327
rect 358 -355 386 -327
rect 420 -355 448 -327
rect -448 -417 -420 -389
rect -386 -417 -358 -389
rect -324 -417 -296 -389
rect -262 -417 -234 -389
rect -200 -417 -172 -389
rect -138 -417 -110 -389
rect -76 -417 -48 -389
rect -14 -417 14 -389
rect 48 -417 76 -389
rect 110 -417 138 -389
rect 172 -417 200 -389
rect 234 -417 262 -389
rect 296 -417 324 -389
rect 358 -417 386 -389
rect 420 -417 448 -389
rect -448 -479 -420 -451
rect -386 -479 -358 -451
rect -324 -479 -296 -451
rect -262 -479 -234 -451
rect -200 -479 -172 -451
rect -138 -479 -110 -451
rect -76 -479 -48 -451
rect -14 -479 14 -451
rect 48 -479 76 -451
rect 110 -479 138 -451
rect 172 -479 200 -451
rect 234 -479 262 -451
rect 296 -479 324 -451
rect 358 -479 386 -451
rect 420 -479 448 -451
rect -448 -541 -420 -513
rect -386 -541 -358 -513
rect -324 -541 -296 -513
rect -262 -541 -234 -513
rect -200 -541 -172 -513
rect -138 -541 -110 -513
rect -76 -541 -48 -513
rect -14 -541 14 -513
rect 48 -541 76 -513
rect 110 -541 138 -513
rect 172 -541 200 -513
rect 234 -541 262 -513
rect 296 -541 324 -513
rect 358 -541 386 -513
rect 420 -541 448 -513
rect -448 -603 -420 -575
rect -386 -603 -358 -575
rect -324 -603 -296 -575
rect -262 -603 -234 -575
rect -200 -603 -172 -575
rect -138 -603 -110 -575
rect -76 -603 -48 -575
rect -14 -603 14 -575
rect 48 -603 76 -575
rect 110 -603 138 -575
rect 172 -603 200 -575
rect 234 -603 262 -575
rect 296 -603 324 -575
rect 358 -603 386 -575
rect 420 -603 448 -575
rect -448 -665 -420 -637
rect -386 -665 -358 -637
rect -324 -665 -296 -637
rect -262 -665 -234 -637
rect -200 -665 -172 -637
rect -138 -665 -110 -637
rect -76 -665 -48 -637
rect -14 -665 14 -637
rect 48 -665 76 -637
rect 110 -665 138 -637
rect 172 -665 200 -637
rect 234 -665 262 -637
rect 296 -665 324 -637
rect 358 -665 386 -637
rect 420 -665 448 -637
rect -448 -727 -420 -699
rect -386 -727 -358 -699
rect -324 -727 -296 -699
rect -262 -727 -234 -699
rect -200 -727 -172 -699
rect -138 -727 -110 -699
rect -76 -727 -48 -699
rect -14 -727 14 -699
rect 48 -727 76 -699
rect 110 -727 138 -699
rect 172 -727 200 -699
rect 234 -727 262 -699
rect 296 -727 324 -699
rect 358 -727 386 -699
rect 420 -727 448 -699
<< metal3 >>
rect -453 727 453 732
rect -453 699 -448 727
rect -420 699 -386 727
rect -358 699 -324 727
rect -296 699 -262 727
rect -234 699 -200 727
rect -172 699 -138 727
rect -110 699 -76 727
rect -48 699 -14 727
rect 14 699 48 727
rect 76 699 110 727
rect 138 699 172 727
rect 200 699 234 727
rect 262 699 296 727
rect 324 699 358 727
rect 386 699 420 727
rect 448 699 453 727
rect -453 665 453 699
rect -453 637 -448 665
rect -420 637 -386 665
rect -358 637 -324 665
rect -296 637 -262 665
rect -234 637 -200 665
rect -172 637 -138 665
rect -110 637 -76 665
rect -48 637 -14 665
rect 14 637 48 665
rect 76 637 110 665
rect 138 637 172 665
rect 200 637 234 665
rect 262 637 296 665
rect 324 637 358 665
rect 386 637 420 665
rect 448 637 453 665
rect -453 603 453 637
rect -453 575 -448 603
rect -420 575 -386 603
rect -358 575 -324 603
rect -296 575 -262 603
rect -234 575 -200 603
rect -172 575 -138 603
rect -110 575 -76 603
rect -48 575 -14 603
rect 14 575 48 603
rect 76 575 110 603
rect 138 575 172 603
rect 200 575 234 603
rect 262 575 296 603
rect 324 575 358 603
rect 386 575 420 603
rect 448 575 453 603
rect -453 541 453 575
rect -453 513 -448 541
rect -420 513 -386 541
rect -358 513 -324 541
rect -296 513 -262 541
rect -234 513 -200 541
rect -172 513 -138 541
rect -110 513 -76 541
rect -48 513 -14 541
rect 14 513 48 541
rect 76 513 110 541
rect 138 513 172 541
rect 200 513 234 541
rect 262 513 296 541
rect 324 513 358 541
rect 386 513 420 541
rect 448 513 453 541
rect -453 479 453 513
rect -453 451 -448 479
rect -420 451 -386 479
rect -358 451 -324 479
rect -296 451 -262 479
rect -234 451 -200 479
rect -172 451 -138 479
rect -110 451 -76 479
rect -48 451 -14 479
rect 14 451 48 479
rect 76 451 110 479
rect 138 451 172 479
rect 200 451 234 479
rect 262 451 296 479
rect 324 451 358 479
rect 386 451 420 479
rect 448 451 453 479
rect -453 417 453 451
rect -453 389 -448 417
rect -420 389 -386 417
rect -358 389 -324 417
rect -296 389 -262 417
rect -234 389 -200 417
rect -172 389 -138 417
rect -110 389 -76 417
rect -48 389 -14 417
rect 14 389 48 417
rect 76 389 110 417
rect 138 389 172 417
rect 200 389 234 417
rect 262 389 296 417
rect 324 389 358 417
rect 386 389 420 417
rect 448 389 453 417
rect -453 355 453 389
rect -453 327 -448 355
rect -420 327 -386 355
rect -358 327 -324 355
rect -296 327 -262 355
rect -234 327 -200 355
rect -172 327 -138 355
rect -110 327 -76 355
rect -48 327 -14 355
rect 14 327 48 355
rect 76 327 110 355
rect 138 327 172 355
rect 200 327 234 355
rect 262 327 296 355
rect 324 327 358 355
rect 386 327 420 355
rect 448 327 453 355
rect -453 293 453 327
rect -453 265 -448 293
rect -420 265 -386 293
rect -358 265 -324 293
rect -296 265 -262 293
rect -234 265 -200 293
rect -172 265 -138 293
rect -110 265 -76 293
rect -48 265 -14 293
rect 14 265 48 293
rect 76 265 110 293
rect 138 265 172 293
rect 200 265 234 293
rect 262 265 296 293
rect 324 265 358 293
rect 386 265 420 293
rect 448 265 453 293
rect -453 231 453 265
rect -453 203 -448 231
rect -420 203 -386 231
rect -358 203 -324 231
rect -296 203 -262 231
rect -234 203 -200 231
rect -172 203 -138 231
rect -110 203 -76 231
rect -48 203 -14 231
rect 14 203 48 231
rect 76 203 110 231
rect 138 203 172 231
rect 200 203 234 231
rect 262 203 296 231
rect 324 203 358 231
rect 386 203 420 231
rect 448 203 453 231
rect -453 169 453 203
rect -453 141 -448 169
rect -420 141 -386 169
rect -358 141 -324 169
rect -296 141 -262 169
rect -234 141 -200 169
rect -172 141 -138 169
rect -110 141 -76 169
rect -48 141 -14 169
rect 14 141 48 169
rect 76 141 110 169
rect 138 141 172 169
rect 200 141 234 169
rect 262 141 296 169
rect 324 141 358 169
rect 386 141 420 169
rect 448 141 453 169
rect -453 107 453 141
rect -453 79 -448 107
rect -420 79 -386 107
rect -358 79 -324 107
rect -296 79 -262 107
rect -234 79 -200 107
rect -172 79 -138 107
rect -110 79 -76 107
rect -48 79 -14 107
rect 14 79 48 107
rect 76 79 110 107
rect 138 79 172 107
rect 200 79 234 107
rect 262 79 296 107
rect 324 79 358 107
rect 386 79 420 107
rect 448 79 453 107
rect -453 45 453 79
rect -453 17 -448 45
rect -420 17 -386 45
rect -358 17 -324 45
rect -296 17 -262 45
rect -234 17 -200 45
rect -172 17 -138 45
rect -110 17 -76 45
rect -48 17 -14 45
rect 14 17 48 45
rect 76 17 110 45
rect 138 17 172 45
rect 200 17 234 45
rect 262 17 296 45
rect 324 17 358 45
rect 386 17 420 45
rect 448 17 453 45
rect -453 -17 453 17
rect -453 -45 -448 -17
rect -420 -45 -386 -17
rect -358 -45 -324 -17
rect -296 -45 -262 -17
rect -234 -45 -200 -17
rect -172 -45 -138 -17
rect -110 -45 -76 -17
rect -48 -45 -14 -17
rect 14 -45 48 -17
rect 76 -45 110 -17
rect 138 -45 172 -17
rect 200 -45 234 -17
rect 262 -45 296 -17
rect 324 -45 358 -17
rect 386 -45 420 -17
rect 448 -45 453 -17
rect -453 -79 453 -45
rect -453 -107 -448 -79
rect -420 -107 -386 -79
rect -358 -107 -324 -79
rect -296 -107 -262 -79
rect -234 -107 -200 -79
rect -172 -107 -138 -79
rect -110 -107 -76 -79
rect -48 -107 -14 -79
rect 14 -107 48 -79
rect 76 -107 110 -79
rect 138 -107 172 -79
rect 200 -107 234 -79
rect 262 -107 296 -79
rect 324 -107 358 -79
rect 386 -107 420 -79
rect 448 -107 453 -79
rect -453 -141 453 -107
rect -453 -169 -448 -141
rect -420 -169 -386 -141
rect -358 -169 -324 -141
rect -296 -169 -262 -141
rect -234 -169 -200 -141
rect -172 -169 -138 -141
rect -110 -169 -76 -141
rect -48 -169 -14 -141
rect 14 -169 48 -141
rect 76 -169 110 -141
rect 138 -169 172 -141
rect 200 -169 234 -141
rect 262 -169 296 -141
rect 324 -169 358 -141
rect 386 -169 420 -141
rect 448 -169 453 -141
rect -453 -203 453 -169
rect -453 -231 -448 -203
rect -420 -231 -386 -203
rect -358 -231 -324 -203
rect -296 -231 -262 -203
rect -234 -231 -200 -203
rect -172 -231 -138 -203
rect -110 -231 -76 -203
rect -48 -231 -14 -203
rect 14 -231 48 -203
rect 76 -231 110 -203
rect 138 -231 172 -203
rect 200 -231 234 -203
rect 262 -231 296 -203
rect 324 -231 358 -203
rect 386 -231 420 -203
rect 448 -231 453 -203
rect -453 -265 453 -231
rect -453 -293 -448 -265
rect -420 -293 -386 -265
rect -358 -293 -324 -265
rect -296 -293 -262 -265
rect -234 -293 -200 -265
rect -172 -293 -138 -265
rect -110 -293 -76 -265
rect -48 -293 -14 -265
rect 14 -293 48 -265
rect 76 -293 110 -265
rect 138 -293 172 -265
rect 200 -293 234 -265
rect 262 -293 296 -265
rect 324 -293 358 -265
rect 386 -293 420 -265
rect 448 -293 453 -265
rect -453 -327 453 -293
rect -453 -355 -448 -327
rect -420 -355 -386 -327
rect -358 -355 -324 -327
rect -296 -355 -262 -327
rect -234 -355 -200 -327
rect -172 -355 -138 -327
rect -110 -355 -76 -327
rect -48 -355 -14 -327
rect 14 -355 48 -327
rect 76 -355 110 -327
rect 138 -355 172 -327
rect 200 -355 234 -327
rect 262 -355 296 -327
rect 324 -355 358 -327
rect 386 -355 420 -327
rect 448 -355 453 -327
rect -453 -389 453 -355
rect -453 -417 -448 -389
rect -420 -417 -386 -389
rect -358 -417 -324 -389
rect -296 -417 -262 -389
rect -234 -417 -200 -389
rect -172 -417 -138 -389
rect -110 -417 -76 -389
rect -48 -417 -14 -389
rect 14 -417 48 -389
rect 76 -417 110 -389
rect 138 -417 172 -389
rect 200 -417 234 -389
rect 262 -417 296 -389
rect 324 -417 358 -389
rect 386 -417 420 -389
rect 448 -417 453 -389
rect -453 -451 453 -417
rect -453 -479 -448 -451
rect -420 -479 -386 -451
rect -358 -479 -324 -451
rect -296 -479 -262 -451
rect -234 -479 -200 -451
rect -172 -479 -138 -451
rect -110 -479 -76 -451
rect -48 -479 -14 -451
rect 14 -479 48 -451
rect 76 -479 110 -451
rect 138 -479 172 -451
rect 200 -479 234 -451
rect 262 -479 296 -451
rect 324 -479 358 -451
rect 386 -479 420 -451
rect 448 -479 453 -451
rect -453 -513 453 -479
rect -453 -541 -448 -513
rect -420 -541 -386 -513
rect -358 -541 -324 -513
rect -296 -541 -262 -513
rect -234 -541 -200 -513
rect -172 -541 -138 -513
rect -110 -541 -76 -513
rect -48 -541 -14 -513
rect 14 -541 48 -513
rect 76 -541 110 -513
rect 138 -541 172 -513
rect 200 -541 234 -513
rect 262 -541 296 -513
rect 324 -541 358 -513
rect 386 -541 420 -513
rect 448 -541 453 -513
rect -453 -575 453 -541
rect -453 -603 -448 -575
rect -420 -603 -386 -575
rect -358 -603 -324 -575
rect -296 -603 -262 -575
rect -234 -603 -200 -575
rect -172 -603 -138 -575
rect -110 -603 -76 -575
rect -48 -603 -14 -575
rect 14 -603 48 -575
rect 76 -603 110 -575
rect 138 -603 172 -575
rect 200 -603 234 -575
rect 262 -603 296 -575
rect 324 -603 358 -575
rect 386 -603 420 -575
rect 448 -603 453 -575
rect -453 -637 453 -603
rect -453 -665 -448 -637
rect -420 -665 -386 -637
rect -358 -665 -324 -637
rect -296 -665 -262 -637
rect -234 -665 -200 -637
rect -172 -665 -138 -637
rect -110 -665 -76 -637
rect -48 -665 -14 -637
rect 14 -665 48 -637
rect 76 -665 110 -637
rect 138 -665 172 -637
rect 200 -665 234 -637
rect 262 -665 296 -637
rect 324 -665 358 -637
rect 386 -665 420 -637
rect 448 -665 453 -637
rect -453 -699 453 -665
rect -453 -727 -448 -699
rect -420 -727 -386 -699
rect -358 -727 -324 -699
rect -296 -727 -262 -699
rect -234 -727 -200 -699
rect -172 -727 -138 -699
rect -110 -727 -76 -699
rect -48 -727 -14 -699
rect 14 -727 48 -699
rect 76 -727 110 -699
rect 138 -727 172 -699
rect 200 -727 234 -699
rect 262 -727 296 -699
rect 324 -727 358 -699
rect 386 -727 420 -699
rect 448 -727 453 -699
rect -453 -732 453 -727
<< end >>
