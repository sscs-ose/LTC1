magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2045 -4677 2045 4677
<< psubdiff >>
rect -45 2655 45 2677
rect -45 -2655 -23 2655
rect 23 -2655 45 2655
rect -45 -2677 45 -2655
<< psubdiffcont >>
rect -23 -2655 23 2655
<< metal1 >>
rect -34 2655 34 2666
rect -34 -2655 -23 2655
rect 23 -2655 34 2655
rect -34 -2666 34 -2655
<< end >>
