magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1253 -1019 1253 1019
<< metal1 >>
rect -253 13 253 19
rect -253 -13 -247 13
rect 247 -13 253 13
rect -253 -19 253 -13
<< via1 >>
rect -247 -13 247 13
<< metal2 >>
rect -253 13 253 19
rect -253 -13 -247 13
rect 247 -13 253 13
rect -253 -19 253 -13
<< end >>
