magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2107 -4959 2107 4959
<< psubdiff >>
rect -107 2937 107 2959
rect -107 2891 -85 2937
rect -39 2891 39 2937
rect 85 2891 107 2937
rect -107 2813 107 2891
rect -107 2767 -85 2813
rect -39 2767 39 2813
rect 85 2767 107 2813
rect -107 2689 107 2767
rect -107 2643 -85 2689
rect -39 2643 39 2689
rect 85 2643 107 2689
rect -107 2565 107 2643
rect -107 2519 -85 2565
rect -39 2519 39 2565
rect 85 2519 107 2565
rect -107 2441 107 2519
rect -107 2395 -85 2441
rect -39 2395 39 2441
rect 85 2395 107 2441
rect -107 2317 107 2395
rect -107 2271 -85 2317
rect -39 2271 39 2317
rect 85 2271 107 2317
rect -107 2193 107 2271
rect -107 2147 -85 2193
rect -39 2147 39 2193
rect 85 2147 107 2193
rect -107 2069 107 2147
rect -107 2023 -85 2069
rect -39 2023 39 2069
rect 85 2023 107 2069
rect -107 1945 107 2023
rect -107 1899 -85 1945
rect -39 1899 39 1945
rect 85 1899 107 1945
rect -107 1821 107 1899
rect -107 1775 -85 1821
rect -39 1775 39 1821
rect 85 1775 107 1821
rect -107 1697 107 1775
rect -107 1651 -85 1697
rect -39 1651 39 1697
rect 85 1651 107 1697
rect -107 1573 107 1651
rect -107 1527 -85 1573
rect -39 1527 39 1573
rect 85 1527 107 1573
rect -107 1449 107 1527
rect -107 1403 -85 1449
rect -39 1403 39 1449
rect 85 1403 107 1449
rect -107 1325 107 1403
rect -107 1279 -85 1325
rect -39 1279 39 1325
rect 85 1279 107 1325
rect -107 1201 107 1279
rect -107 1155 -85 1201
rect -39 1155 39 1201
rect 85 1155 107 1201
rect -107 1077 107 1155
rect -107 1031 -85 1077
rect -39 1031 39 1077
rect 85 1031 107 1077
rect -107 953 107 1031
rect -107 907 -85 953
rect -39 907 39 953
rect 85 907 107 953
rect -107 829 107 907
rect -107 783 -85 829
rect -39 783 39 829
rect 85 783 107 829
rect -107 705 107 783
rect -107 659 -85 705
rect -39 659 39 705
rect 85 659 107 705
rect -107 581 107 659
rect -107 535 -85 581
rect -39 535 39 581
rect 85 535 107 581
rect -107 457 107 535
rect -107 411 -85 457
rect -39 411 39 457
rect 85 411 107 457
rect -107 333 107 411
rect -107 287 -85 333
rect -39 287 39 333
rect 85 287 107 333
rect -107 209 107 287
rect -107 163 -85 209
rect -39 163 39 209
rect 85 163 107 209
rect -107 85 107 163
rect -107 39 -85 85
rect -39 39 39 85
rect 85 39 107 85
rect -107 -39 107 39
rect -107 -85 -85 -39
rect -39 -85 39 -39
rect 85 -85 107 -39
rect -107 -163 107 -85
rect -107 -209 -85 -163
rect -39 -209 39 -163
rect 85 -209 107 -163
rect -107 -287 107 -209
rect -107 -333 -85 -287
rect -39 -333 39 -287
rect 85 -333 107 -287
rect -107 -411 107 -333
rect -107 -457 -85 -411
rect -39 -457 39 -411
rect 85 -457 107 -411
rect -107 -535 107 -457
rect -107 -581 -85 -535
rect -39 -581 39 -535
rect 85 -581 107 -535
rect -107 -659 107 -581
rect -107 -705 -85 -659
rect -39 -705 39 -659
rect 85 -705 107 -659
rect -107 -783 107 -705
rect -107 -829 -85 -783
rect -39 -829 39 -783
rect 85 -829 107 -783
rect -107 -907 107 -829
rect -107 -953 -85 -907
rect -39 -953 39 -907
rect 85 -953 107 -907
rect -107 -1031 107 -953
rect -107 -1077 -85 -1031
rect -39 -1077 39 -1031
rect 85 -1077 107 -1031
rect -107 -1155 107 -1077
rect -107 -1201 -85 -1155
rect -39 -1201 39 -1155
rect 85 -1201 107 -1155
rect -107 -1279 107 -1201
rect -107 -1325 -85 -1279
rect -39 -1325 39 -1279
rect 85 -1325 107 -1279
rect -107 -1403 107 -1325
rect -107 -1449 -85 -1403
rect -39 -1449 39 -1403
rect 85 -1449 107 -1403
rect -107 -1527 107 -1449
rect -107 -1573 -85 -1527
rect -39 -1573 39 -1527
rect 85 -1573 107 -1527
rect -107 -1651 107 -1573
rect -107 -1697 -85 -1651
rect -39 -1697 39 -1651
rect 85 -1697 107 -1651
rect -107 -1775 107 -1697
rect -107 -1821 -85 -1775
rect -39 -1821 39 -1775
rect 85 -1821 107 -1775
rect -107 -1899 107 -1821
rect -107 -1945 -85 -1899
rect -39 -1945 39 -1899
rect 85 -1945 107 -1899
rect -107 -2023 107 -1945
rect -107 -2069 -85 -2023
rect -39 -2069 39 -2023
rect 85 -2069 107 -2023
rect -107 -2147 107 -2069
rect -107 -2193 -85 -2147
rect -39 -2193 39 -2147
rect 85 -2193 107 -2147
rect -107 -2271 107 -2193
rect -107 -2317 -85 -2271
rect -39 -2317 39 -2271
rect 85 -2317 107 -2271
rect -107 -2395 107 -2317
rect -107 -2441 -85 -2395
rect -39 -2441 39 -2395
rect 85 -2441 107 -2395
rect -107 -2519 107 -2441
rect -107 -2565 -85 -2519
rect -39 -2565 39 -2519
rect 85 -2565 107 -2519
rect -107 -2643 107 -2565
rect -107 -2689 -85 -2643
rect -39 -2689 39 -2643
rect 85 -2689 107 -2643
rect -107 -2767 107 -2689
rect -107 -2813 -85 -2767
rect -39 -2813 39 -2767
rect 85 -2813 107 -2767
rect -107 -2891 107 -2813
rect -107 -2937 -85 -2891
rect -39 -2937 39 -2891
rect 85 -2937 107 -2891
rect -107 -2959 107 -2937
<< psubdiffcont >>
rect -85 2891 -39 2937
rect 39 2891 85 2937
rect -85 2767 -39 2813
rect 39 2767 85 2813
rect -85 2643 -39 2689
rect 39 2643 85 2689
rect -85 2519 -39 2565
rect 39 2519 85 2565
rect -85 2395 -39 2441
rect 39 2395 85 2441
rect -85 2271 -39 2317
rect 39 2271 85 2317
rect -85 2147 -39 2193
rect 39 2147 85 2193
rect -85 2023 -39 2069
rect 39 2023 85 2069
rect -85 1899 -39 1945
rect 39 1899 85 1945
rect -85 1775 -39 1821
rect 39 1775 85 1821
rect -85 1651 -39 1697
rect 39 1651 85 1697
rect -85 1527 -39 1573
rect 39 1527 85 1573
rect -85 1403 -39 1449
rect 39 1403 85 1449
rect -85 1279 -39 1325
rect 39 1279 85 1325
rect -85 1155 -39 1201
rect 39 1155 85 1201
rect -85 1031 -39 1077
rect 39 1031 85 1077
rect -85 907 -39 953
rect 39 907 85 953
rect -85 783 -39 829
rect 39 783 85 829
rect -85 659 -39 705
rect 39 659 85 705
rect -85 535 -39 581
rect 39 535 85 581
rect -85 411 -39 457
rect 39 411 85 457
rect -85 287 -39 333
rect 39 287 85 333
rect -85 163 -39 209
rect 39 163 85 209
rect -85 39 -39 85
rect 39 39 85 85
rect -85 -85 -39 -39
rect 39 -85 85 -39
rect -85 -209 -39 -163
rect 39 -209 85 -163
rect -85 -333 -39 -287
rect 39 -333 85 -287
rect -85 -457 -39 -411
rect 39 -457 85 -411
rect -85 -581 -39 -535
rect 39 -581 85 -535
rect -85 -705 -39 -659
rect 39 -705 85 -659
rect -85 -829 -39 -783
rect 39 -829 85 -783
rect -85 -953 -39 -907
rect 39 -953 85 -907
rect -85 -1077 -39 -1031
rect 39 -1077 85 -1031
rect -85 -1201 -39 -1155
rect 39 -1201 85 -1155
rect -85 -1325 -39 -1279
rect 39 -1325 85 -1279
rect -85 -1449 -39 -1403
rect 39 -1449 85 -1403
rect -85 -1573 -39 -1527
rect 39 -1573 85 -1527
rect -85 -1697 -39 -1651
rect 39 -1697 85 -1651
rect -85 -1821 -39 -1775
rect 39 -1821 85 -1775
rect -85 -1945 -39 -1899
rect 39 -1945 85 -1899
rect -85 -2069 -39 -2023
rect 39 -2069 85 -2023
rect -85 -2193 -39 -2147
rect 39 -2193 85 -2147
rect -85 -2317 -39 -2271
rect 39 -2317 85 -2271
rect -85 -2441 -39 -2395
rect 39 -2441 85 -2395
rect -85 -2565 -39 -2519
rect 39 -2565 85 -2519
rect -85 -2689 -39 -2643
rect 39 -2689 85 -2643
rect -85 -2813 -39 -2767
rect 39 -2813 85 -2767
rect -85 -2937 -39 -2891
rect 39 -2937 85 -2891
<< metal1 >>
rect -96 2937 96 2948
rect -96 2891 -85 2937
rect -39 2891 39 2937
rect 85 2891 96 2937
rect -96 2813 96 2891
rect -96 2767 -85 2813
rect -39 2767 39 2813
rect 85 2767 96 2813
rect -96 2689 96 2767
rect -96 2643 -85 2689
rect -39 2643 39 2689
rect 85 2643 96 2689
rect -96 2565 96 2643
rect -96 2519 -85 2565
rect -39 2519 39 2565
rect 85 2519 96 2565
rect -96 2441 96 2519
rect -96 2395 -85 2441
rect -39 2395 39 2441
rect 85 2395 96 2441
rect -96 2317 96 2395
rect -96 2271 -85 2317
rect -39 2271 39 2317
rect 85 2271 96 2317
rect -96 2193 96 2271
rect -96 2147 -85 2193
rect -39 2147 39 2193
rect 85 2147 96 2193
rect -96 2069 96 2147
rect -96 2023 -85 2069
rect -39 2023 39 2069
rect 85 2023 96 2069
rect -96 1945 96 2023
rect -96 1899 -85 1945
rect -39 1899 39 1945
rect 85 1899 96 1945
rect -96 1821 96 1899
rect -96 1775 -85 1821
rect -39 1775 39 1821
rect 85 1775 96 1821
rect -96 1697 96 1775
rect -96 1651 -85 1697
rect -39 1651 39 1697
rect 85 1651 96 1697
rect -96 1573 96 1651
rect -96 1527 -85 1573
rect -39 1527 39 1573
rect 85 1527 96 1573
rect -96 1449 96 1527
rect -96 1403 -85 1449
rect -39 1403 39 1449
rect 85 1403 96 1449
rect -96 1325 96 1403
rect -96 1279 -85 1325
rect -39 1279 39 1325
rect 85 1279 96 1325
rect -96 1201 96 1279
rect -96 1155 -85 1201
rect -39 1155 39 1201
rect 85 1155 96 1201
rect -96 1077 96 1155
rect -96 1031 -85 1077
rect -39 1031 39 1077
rect 85 1031 96 1077
rect -96 953 96 1031
rect -96 907 -85 953
rect -39 907 39 953
rect 85 907 96 953
rect -96 829 96 907
rect -96 783 -85 829
rect -39 783 39 829
rect 85 783 96 829
rect -96 705 96 783
rect -96 659 -85 705
rect -39 659 39 705
rect 85 659 96 705
rect -96 581 96 659
rect -96 535 -85 581
rect -39 535 39 581
rect 85 535 96 581
rect -96 457 96 535
rect -96 411 -85 457
rect -39 411 39 457
rect 85 411 96 457
rect -96 333 96 411
rect -96 287 -85 333
rect -39 287 39 333
rect 85 287 96 333
rect -96 209 96 287
rect -96 163 -85 209
rect -39 163 39 209
rect 85 163 96 209
rect -96 85 96 163
rect -96 39 -85 85
rect -39 39 39 85
rect 85 39 96 85
rect -96 -39 96 39
rect -96 -85 -85 -39
rect -39 -85 39 -39
rect 85 -85 96 -39
rect -96 -163 96 -85
rect -96 -209 -85 -163
rect -39 -209 39 -163
rect 85 -209 96 -163
rect -96 -287 96 -209
rect -96 -333 -85 -287
rect -39 -333 39 -287
rect 85 -333 96 -287
rect -96 -411 96 -333
rect -96 -457 -85 -411
rect -39 -457 39 -411
rect 85 -457 96 -411
rect -96 -535 96 -457
rect -96 -581 -85 -535
rect -39 -581 39 -535
rect 85 -581 96 -535
rect -96 -659 96 -581
rect -96 -705 -85 -659
rect -39 -705 39 -659
rect 85 -705 96 -659
rect -96 -783 96 -705
rect -96 -829 -85 -783
rect -39 -829 39 -783
rect 85 -829 96 -783
rect -96 -907 96 -829
rect -96 -953 -85 -907
rect -39 -953 39 -907
rect 85 -953 96 -907
rect -96 -1031 96 -953
rect -96 -1077 -85 -1031
rect -39 -1077 39 -1031
rect 85 -1077 96 -1031
rect -96 -1155 96 -1077
rect -96 -1201 -85 -1155
rect -39 -1201 39 -1155
rect 85 -1201 96 -1155
rect -96 -1279 96 -1201
rect -96 -1325 -85 -1279
rect -39 -1325 39 -1279
rect 85 -1325 96 -1279
rect -96 -1403 96 -1325
rect -96 -1449 -85 -1403
rect -39 -1449 39 -1403
rect 85 -1449 96 -1403
rect -96 -1527 96 -1449
rect -96 -1573 -85 -1527
rect -39 -1573 39 -1527
rect 85 -1573 96 -1527
rect -96 -1651 96 -1573
rect -96 -1697 -85 -1651
rect -39 -1697 39 -1651
rect 85 -1697 96 -1651
rect -96 -1775 96 -1697
rect -96 -1821 -85 -1775
rect -39 -1821 39 -1775
rect 85 -1821 96 -1775
rect -96 -1899 96 -1821
rect -96 -1945 -85 -1899
rect -39 -1945 39 -1899
rect 85 -1945 96 -1899
rect -96 -2023 96 -1945
rect -96 -2069 -85 -2023
rect -39 -2069 39 -2023
rect 85 -2069 96 -2023
rect -96 -2147 96 -2069
rect -96 -2193 -85 -2147
rect -39 -2193 39 -2147
rect 85 -2193 96 -2147
rect -96 -2271 96 -2193
rect -96 -2317 -85 -2271
rect -39 -2317 39 -2271
rect 85 -2317 96 -2271
rect -96 -2395 96 -2317
rect -96 -2441 -85 -2395
rect -39 -2441 39 -2395
rect 85 -2441 96 -2395
rect -96 -2519 96 -2441
rect -96 -2565 -85 -2519
rect -39 -2565 39 -2519
rect 85 -2565 96 -2519
rect -96 -2643 96 -2565
rect -96 -2689 -85 -2643
rect -39 -2689 39 -2643
rect 85 -2689 96 -2643
rect -96 -2767 96 -2689
rect -96 -2813 -85 -2767
rect -39 -2813 39 -2767
rect 85 -2813 96 -2767
rect -96 -2891 96 -2813
rect -96 -2937 -85 -2891
rect -39 -2937 39 -2891
rect 85 -2937 96 -2891
rect -96 -2948 96 -2937
<< end >>
