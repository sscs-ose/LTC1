magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2038 -3103 2038 3103
<< metal2 >>
rect -38 1093 38 1103
rect -38 1037 -28 1093
rect 28 1037 38 1093
rect -38 951 38 1037
rect -38 895 -28 951
rect 28 895 38 951
rect -38 809 38 895
rect -38 753 -28 809
rect 28 753 38 809
rect -38 667 38 753
rect -38 611 -28 667
rect 28 611 38 667
rect -38 525 38 611
rect -38 469 -28 525
rect 28 469 38 525
rect -38 383 38 469
rect -38 327 -28 383
rect 28 327 38 383
rect -38 241 38 327
rect -38 185 -28 241
rect 28 185 38 241
rect -38 99 38 185
rect -38 43 -28 99
rect 28 43 38 99
rect -38 -43 38 43
rect -38 -99 -28 -43
rect 28 -99 38 -43
rect -38 -185 38 -99
rect -38 -241 -28 -185
rect 28 -241 38 -185
rect -38 -327 38 -241
rect -38 -383 -28 -327
rect 28 -383 38 -327
rect -38 -469 38 -383
rect -38 -525 -28 -469
rect 28 -525 38 -469
rect -38 -611 38 -525
rect -38 -667 -28 -611
rect 28 -667 38 -611
rect -38 -753 38 -667
rect -38 -809 -28 -753
rect 28 -809 38 -753
rect -38 -895 38 -809
rect -38 -951 -28 -895
rect 28 -951 38 -895
rect -38 -1037 38 -951
rect -38 -1093 -28 -1037
rect 28 -1093 38 -1037
rect -38 -1103 38 -1093
<< via2 >>
rect -28 1037 28 1093
rect -28 895 28 951
rect -28 753 28 809
rect -28 611 28 667
rect -28 469 28 525
rect -28 327 28 383
rect -28 185 28 241
rect -28 43 28 99
rect -28 -99 28 -43
rect -28 -241 28 -185
rect -28 -383 28 -327
rect -28 -525 28 -469
rect -28 -667 28 -611
rect -28 -809 28 -753
rect -28 -951 28 -895
rect -28 -1093 28 -1037
<< metal3 >>
rect -38 1093 38 1103
rect -38 1037 -28 1093
rect 28 1037 38 1093
rect -38 951 38 1037
rect -38 895 -28 951
rect 28 895 38 951
rect -38 809 38 895
rect -38 753 -28 809
rect 28 753 38 809
rect -38 667 38 753
rect -38 611 -28 667
rect 28 611 38 667
rect -38 525 38 611
rect -38 469 -28 525
rect 28 469 38 525
rect -38 383 38 469
rect -38 327 -28 383
rect 28 327 38 383
rect -38 241 38 327
rect -38 185 -28 241
rect 28 185 38 241
rect -38 99 38 185
rect -38 43 -28 99
rect 28 43 38 99
rect -38 -43 38 43
rect -38 -99 -28 -43
rect 28 -99 38 -43
rect -38 -185 38 -99
rect -38 -241 -28 -185
rect 28 -241 38 -185
rect -38 -327 38 -241
rect -38 -383 -28 -327
rect 28 -383 38 -327
rect -38 -469 38 -383
rect -38 -525 -28 -469
rect 28 -525 38 -469
rect -38 -611 38 -525
rect -38 -667 -28 -611
rect 28 -667 38 -611
rect -38 -753 38 -667
rect -38 -809 -28 -753
rect 28 -809 38 -753
rect -38 -895 38 -809
rect -38 -951 -28 -895
rect 28 -951 38 -895
rect -38 -1037 38 -951
rect -38 -1093 -28 -1037
rect 28 -1093 38 -1037
rect -38 -1103 38 -1093
<< end >>
