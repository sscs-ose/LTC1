magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1283 1019 1283
<< metal2 >>
rect -19 278 19 283
rect -19 250 -14 278
rect 14 250 19 278
rect -19 212 19 250
rect -19 184 -14 212
rect 14 184 19 212
rect -19 146 19 184
rect -19 118 -14 146
rect 14 118 19 146
rect -19 80 19 118
rect -19 52 -14 80
rect 14 52 19 80
rect -19 14 19 52
rect -19 -14 -14 14
rect 14 -14 19 14
rect -19 -52 19 -14
rect -19 -80 -14 -52
rect 14 -80 19 -52
rect -19 -118 19 -80
rect -19 -146 -14 -118
rect 14 -146 19 -118
rect -19 -184 19 -146
rect -19 -212 -14 -184
rect 14 -212 19 -184
rect -19 -250 19 -212
rect -19 -278 -14 -250
rect 14 -278 19 -250
rect -19 -283 19 -278
<< via2 >>
rect -14 250 14 278
rect -14 184 14 212
rect -14 118 14 146
rect -14 52 14 80
rect -14 -14 14 14
rect -14 -80 14 -52
rect -14 -146 14 -118
rect -14 -212 14 -184
rect -14 -278 14 -250
<< metal3 >>
rect -19 278 19 283
rect -19 250 -14 278
rect 14 250 19 278
rect -19 212 19 250
rect -19 184 -14 212
rect 14 184 19 212
rect -19 146 19 184
rect -19 118 -14 146
rect 14 118 19 146
rect -19 80 19 118
rect -19 52 -14 80
rect 14 52 19 80
rect -19 14 19 52
rect -19 -14 -14 14
rect 14 -14 19 14
rect -19 -52 19 -14
rect -19 -80 -14 -52
rect 14 -80 19 -52
rect -19 -118 19 -80
rect -19 -146 -14 -118
rect 14 -146 19 -118
rect -19 -184 19 -146
rect -19 -212 -14 -184
rect 14 -212 19 -184
rect -19 -250 19 -212
rect -19 -278 -14 -250
rect 14 -278 19 -250
rect -19 -283 19 -278
<< end >>
