* NGSPICE file created from GF_INV16_flat.ext - technology: gf180mcuC

.subckt GF_INV16_flat VDD IN OUT VSS
X0 OUT IN.t0 VDD.t9 VDD.t8 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.35u
X1 VSS IN.t1 OUT.t5 VSS.t7 nfet_03v3 ad=0.364p pd=1.92u as=0.364p ps=1.92u w=1.4u l=0.35u
X2 VDD IN.t2 OUT.t2 VDD.t5 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.35u
X3 VSS IN.t3 OUT.t4 VSS.t4 nfet_03v3 ad=0.616p pd=3.68u as=0.364p ps=1.92u w=1.4u l=0.35u
X4 OUT IN.t4 VSS.t3 VSS.t2 nfet_03v3 ad=0.364p pd=1.92u as=0.616p ps=3.68u w=1.4u l=0.35u
X5 OUT IN.t5 VDD.t4 VDD.t3 pfet_03v3 ad=0.728p pd=3.32u as=1.23p ps=6.48u w=2.8u l=0.35u
X6 OUT IN.t6 VSS.t1 VSS.t0 nfet_03v3 ad=0.364p pd=1.92u as=0.364p ps=1.92u w=1.4u l=0.35u
X7 VDD IN.t7 OUT.t0 VDD.t0 pfet_03v3 ad=1.23p pd=6.48u as=0.728p ps=3.32u w=2.8u l=0.35u
R0 IN.n0 IN.t7 40.8805
R1 IN.n1 IN.t0 40.8805
R2 IN.n2 IN.t2 40.8805
R3 IN.n3 IN.t5 36.0834
R4 IN.n0 IN.t3 25.8634
R5 IN.n1 IN.t6 25.8634
R6 IN.n2 IN.t1 25.8634
R7 IN.n3 IN.t4 22.1091
R8 IN.n3 IN.n2 17.4409
R9 IN.n1 IN.n0 14.325
R10 IN.n2 IN.n1 14.325
R11 IN IN.n3 8.98512
R12 VDD.n8 VDD.t8 46.3367
R13 VDD.n5 VDD.t0 32.3281
R14 VDD.n19 VDD.t3 16.8707
R15 VDD.n15 VDD.t5 16.1643
R16 VDD.n4 VDD.n2 3.94592
R17 VDD.n18 VDD.t4 3.92746
R18 VDD.n14 VDD.n1 3.27746
R19 VDD.n4 VDD.n3 3.1505
R20 VDD.n7 VDD.n6 3.1505
R21 VDD.n6 VDD.n5 3.1505
R22 VDD.n10 VDD.n9 3.1505
R23 VDD.n9 VDD.n8 3.1505
R24 VDD.n13 VDD.n12 3.1505
R25 VDD.n12 VDD.n11 3.1505
R26 VDD.n17 VDD.n16 3.1505
R27 VDD.n16 VDD.n15 3.1505
R28 VDD.n24 VDD.n23 3.1505
R29 VDD.n23 VDD.n22 3.1505
R30 VDD.n21 VDD.n20 3.1505
R31 VDD.n1 VDD.t9 0.6505
R32 VDD.n1 VDD.n0 0.6505
R33 VDD.n20 VDD.n19 0.209419
R34 VDD.n7 VDD.n4 0.117038
R35 VDD.n10 VDD.n7 0.117038
R36 VDD.n13 VDD.n10 0.117038
R37 VDD.n24 VDD.n21 0.117038
R38 VDD.n21 VDD.n18 0.0858846
R39 VDD.n17 VDD.n14 0.0835769
R40 VDD VDD.n17 0.0708846
R41 VDD VDD.n24 0.0466538
R42 VDD.n14 VDD.n13 0.0339615
R43 OUT.n9 OUT.n3 3.58485
R44 OUT.n8 OUT.n7 3.58485
R45 OUT.n9 OUT.n1 3.32833
R46 OUT.n8 OUT.n5 3.32833
R47 OUT.n3 OUT.t4 1.1705
R48 OUT.n3 OUT.n2 1.1705
R49 OUT.n7 OUT.t5 1.1705
R50 OUT.n7 OUT.n6 1.1705
R51 OUT.n9 OUT.n8 0.68137
R52 OUT.n1 OUT.t0 0.6505
R53 OUT.n1 OUT.n0 0.6505
R54 OUT.n5 OUT.t2 0.6505
R55 OUT.n5 OUT.n4 0.6505
R56 OUT OUT.n9 0.297891
R57 VSS.n16 VSS.n15 440.101
R58 VSS.n78 VSS.n77 310.293
R59 VSS.n121 VSS.t2 286.442
R60 VSS.n61 VSS.t0 253.391
R61 VSS.n55 VSS.t4 165.255
R62 VSS.n45 VSS.n44 126.695
R63 VSS.n99 VSS.n98 57.6928
R64 VSS.n124 VSS.t7 16.5259
R65 VSS.n54 VSS.n2 4.79593
R66 VSS.n117 VSS.t3 4.79593
R67 VSS VSS.n1 3.60246
R68 VSS.n79 VSS.n78 2.60204
R69 VSS.n20 VSS.n19 2.6005
R70 VSS.n19 VSS.n18 2.6005
R71 VSS.n48 VSS.n47 2.6005
R72 VSS.n43 VSS.n42 2.6005
R73 VSS.n41 VSS.n40 2.6005
R74 VSS.n38 VSS.n37 2.6005
R75 VSS.n37 VSS.n36 2.6005
R76 VSS.n35 VSS.n34 2.6005
R77 VSS.n34 VSS.n33 2.6005
R78 VSS.n32 VSS.n31 2.6005
R79 VSS.n31 VSS.n30 2.6005
R80 VSS.n29 VSS.n28 2.6005
R81 VSS.n28 VSS.n27 2.6005
R82 VSS.n26 VSS.n25 2.6005
R83 VSS.n25 VSS.n24 2.6005
R84 VSS.n23 VSS.n22 2.6005
R85 VSS.n22 VSS.n21 2.6005
R86 VSS.n17 VSS.n16 2.6005
R87 VSS.n14 VSS.n13 2.6005
R88 VSS.n13 VSS.n12 2.6005
R89 VSS.n11 VSS.n10 2.6005
R90 VSS.n10 VSS.n9 2.6005
R91 VSS.n8 VSS.n7 2.6005
R92 VSS.n7 VSS.n6 2.6005
R93 VSS.n5 VSS.n4 2.6005
R94 VSS.n4 VSS.n3 2.6005
R95 VSS.n66 VSS.n65 2.6005
R96 VSS.n65 VSS.n64 2.6005
R97 VSS.n69 VSS.n68 2.6005
R98 VSS.n68 VSS.n67 2.6005
R99 VSS.n72 VSS.n71 2.6005
R100 VSS.n71 VSS.n70 2.6005
R101 VSS.n75 VSS.n74 2.6005
R102 VSS.n74 VSS.n73 2.6005
R103 VSS.n85 VSS.n84 2.6005
R104 VSS.n84 VSS.n83 2.6005
R105 VSS.n88 VSS.n87 2.6005
R106 VSS.n87 VSS.n86 2.6005
R107 VSS.n91 VSS.n90 2.6005
R108 VSS.n90 VSS.n89 2.6005
R109 VSS.n94 VSS.n93 2.6005
R110 VSS.n93 VSS.n92 2.6005
R111 VSS.n97 VSS.n96 2.6005
R112 VSS.n96 VSS.n95 2.6005
R113 VSS.n101 VSS.n100 2.6005
R114 VSS.n100 VSS.n99 2.6005
R115 VSS.n104 VSS.n103 2.6005
R116 VSS.n106 VSS.n105 2.6005
R117 VSS.n110 VSS.n109 2.6005
R118 VSS.n82 VSS.n81 2.6005
R119 VSS.n81 VSS.n80 2.6005
R120 VSS.n50 VSS.n49 2.6005
R121 VSS.n53 VSS.n52 2.6005
R122 VSS.n52 VSS.n51 2.6005
R123 VSS.n57 VSS.n56 2.6005
R124 VSS.n56 VSS.n55 2.6005
R125 VSS.n60 VSS.n59 2.6005
R126 VSS.n59 VSS.n58 2.6005
R127 VSS.n63 VSS.n62 2.6005
R128 VSS.n62 VSS.n61 2.6005
R129 VSS.n126 VSS.n125 2.6005
R130 VSS.n125 VSS.n124 2.6005
R131 VSS.n123 VSS.n122 2.6005
R132 VSS.n122 VSS.n121 2.6005
R133 VSS.n120 VSS.n119 2.6005
R134 VSS.n119 VSS.n118 2.6005
R135 VSS.n116 VSS.n115 2.6005
R136 VSS.n115 VSS.n114 2.6005
R137 VSS.n113 VSS.n112 2.6005
R138 VSS.n112 VSS.n111 2.6005
R139 VSS.n40 VSS.n39 1.36979
R140 VSS.n103 VSS.n102 1.36965
R141 VSS.n109 VSS.n108 1.36965
R142 VSS.n47 VSS.n46 1.36965
R143 VSS.n1 VSS.t1 1.1705
R144 VSS.n1 VSS.n0 1.1705
R145 VSS.n46 VSS.n45 0.8219
R146 VSS.n108 VSS.n107 0.8219
R147 VSS.n82 VSS.n79 0.127656
R148 VSS.n20 VSS.n17 0.122589
R149 VSS.n78 VSS.n76 0.120158
R150 VSS.n53 VSS.n50 0.119731
R151 VSS.n79 VSS.n75 0.118962
R152 VSS.n23 VSS.n20 0.111968
R153 VSS.n26 VSS.n23 0.111968
R154 VSS.n29 VSS.n26 0.111968
R155 VSS.n32 VSS.n29 0.111968
R156 VSS.n35 VSS.n32 0.111968
R157 VSS.n38 VSS.n35 0.111968
R158 VSS.n41 VSS.n38 0.111968
R159 VSS.n43 VSS.n41 0.111968
R160 VSS.n48 VSS.n43 0.111968
R161 VSS.n85 VSS.n82 0.111968
R162 VSS.n88 VSS.n85 0.111968
R163 VSS.n91 VSS.n88 0.111968
R164 VSS.n94 VSS.n91 0.111968
R165 VSS.n97 VSS.n94 0.111968
R166 VSS.n101 VSS.n97 0.111968
R167 VSS.n104 VSS.n101 0.111968
R168 VSS.n106 VSS.n104 0.111968
R169 VSS.n110 VSS.n106 0.111968
R170 VSS.n17 VSS.n14 0.0966538
R171 VSS.n14 VSS.n11 0.0966538
R172 VSS.n11 VSS.n8 0.0966538
R173 VSS.n8 VSS.n5 0.0966538
R174 VSS.n69 VSS.n66 0.0966538
R175 VSS.n72 VSS.n69 0.0966538
R176 VSS.n75 VSS.n72 0.0966538
R177 VSS.n60 VSS.n57 0.0966538
R178 VSS.n63 VSS.n60 0.0966538
R179 VSS.n126 VSS.n123 0.0966538
R180 VSS.n123 VSS.n120 0.0966538
R181 VSS.n116 VSS.n113 0.0966538
R182 VSS.n117 VSS.n116 0.0858846
R183 VSS.n50 VSS.n48 0.0657294
R184 VSS.n127 VSS.n126 0.0651154
R185 VSS.n113 VSS.n110 0.0598931
R186 VSS.n54 VSS.n53 0.0528077
R187 VSS.n57 VSS.n54 0.0443462
R188 VSS.n127 VSS.n63 0.0320385
R189 VSS VSS.n127 0.0239783
R190 VSS.n120 VSS.n117 0.0112692
C0 VDD IN 0.62f
C1 OUT IN 0.23f
C2 VDD OUT 0.952f
.ends

