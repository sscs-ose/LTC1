magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2045 -9095 2045 9095
<< psubdiff >>
rect -45 7073 45 7095
rect -45 -7073 -23 7073
rect 23 -7073 45 7073
rect -45 -7095 45 -7073
<< psubdiffcont >>
rect -23 -7073 23 7073
<< metal1 >>
rect -34 7073 34 7084
rect -34 -7073 -23 7073
rect 23 -7073 34 7073
rect -34 -7084 34 -7073
<< end >>
