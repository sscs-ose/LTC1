magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -2632 -2180 2632 2180
<< nwell >>
rect -632 -180 632 180
<< pmos >>
rect -458 -50 -358 50
rect -254 -50 -154 50
rect -50 -50 50 50
rect 154 -50 254 50
rect 358 -50 458 50
<< pdiff >>
rect -546 23 -458 50
rect -546 -23 -533 23
rect -487 -23 -458 23
rect -546 -50 -458 -23
rect -358 23 -254 50
rect -358 -23 -329 23
rect -283 -23 -254 23
rect -358 -50 -254 -23
rect -154 23 -50 50
rect -154 -23 -125 23
rect -79 -23 -50 23
rect -154 -50 -50 -23
rect 50 23 154 50
rect 50 -23 79 23
rect 125 -23 154 23
rect 50 -50 154 -23
rect 254 23 358 50
rect 254 -23 283 23
rect 329 -23 358 23
rect 254 -50 358 -23
rect 458 23 546 50
rect 458 -23 487 23
rect 533 -23 546 23
rect 458 -50 546 -23
<< pdiffc >>
rect -533 -23 -487 23
rect -329 -23 -283 23
rect -125 -23 -79 23
rect 79 -23 125 23
rect 283 -23 329 23
rect 487 -23 533 23
<< polysilicon >>
rect -458 50 -358 94
rect -254 50 -154 94
rect -50 50 50 94
rect 154 50 254 94
rect 358 50 458 94
rect -458 -94 -358 -50
rect -254 -94 -154 -50
rect -50 -94 50 -50
rect 154 -94 254 -50
rect 358 -94 458 -50
<< metal1 >>
rect -533 23 -487 48
rect -533 -48 -487 -23
rect -329 23 -283 48
rect -329 -48 -283 -23
rect -125 23 -79 48
rect -125 -48 -79 -23
rect 79 23 125 48
rect 79 -48 125 -23
rect 283 23 329 48
rect 283 -48 329 -23
rect 487 23 533 48
rect 487 -48 533 -23
<< end >>
