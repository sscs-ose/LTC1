magic
tech gf180mcuD
magscale 1 10
timestamp 1713971361
<< checkpaint >>
rect -2090 -2027 25932 9176
<< pwell >>
rect 6991 4685 7927 4953
<< metal1 >>
rect 7054 6973 8052 7077
rect 5860 5758 6162 5843
rect 19018 4885 19138 4925
rect 19018 4833 19051 4885
rect 19103 4833 19138 4885
rect 19018 4795 19138 4833
rect 19224 4882 19344 4922
rect 19224 4830 19257 4882
rect 19309 4830 19344 4882
rect 19224 4792 19344 4830
rect 19416 4869 19536 4909
rect 19416 4817 19449 4869
rect 19501 4817 19536 4869
rect 19416 4779 19536 4817
rect 19604 4863 19724 4903
rect 19604 4811 19637 4863
rect 19689 4811 19724 4863
rect 19604 4773 19724 4811
rect 19831 4874 19951 4914
rect 19831 4822 19864 4874
rect 19916 4822 19951 4874
rect 19831 4784 19951 4822
rect 16154 4134 16971 4346
rect 17810 4016 17915 4427
rect 20697 4055 20802 4419
rect 21896 3994 22039 4446
rect 22540 4053 22654 4416
rect 22731 4022 23135 4118
rect 23481 3927 23860 3946
rect 23481 3912 23932 3927
rect 17167 3866 17300 3911
rect 17167 3814 17209 3866
rect 17261 3814 17300 3866
rect 23481 3860 23504 3912
rect 23556 3860 23646 3912
rect 23698 3860 23785 3912
rect 23837 3860 23932 3912
rect 23481 3845 23932 3860
rect 23481 3825 23860 3845
rect 17167 3694 17300 3814
rect 22811 3699 23024 3741
rect 17167 3654 17490 3694
rect 17167 3602 17224 3654
rect 17276 3602 17398 3654
rect 17450 3602 17490 3654
rect 22811 3647 22823 3699
rect 22875 3647 22943 3699
rect 22995 3647 23024 3699
rect 22811 3608 23024 3647
rect 17167 3578 17490 3602
rect 16145 3288 16962 3500
rect 22874 2837 22982 2860
rect 23311 2847 23695 2858
rect 22874 2785 22899 2837
rect 22951 2785 22982 2837
rect 22874 2695 22982 2785
rect 23310 2837 23768 2847
rect 23310 2785 23354 2837
rect 23406 2785 23479 2837
rect 23531 2785 23625 2837
rect 23677 2785 23768 2837
rect 23310 2775 23768 2785
rect 23311 2764 23695 2775
rect 22874 2643 22899 2695
rect 22951 2643 22982 2695
rect 16150 2324 16967 2536
rect 22874 2523 22982 2643
rect 22874 2471 22899 2523
rect 22951 2471 22982 2523
rect 22874 2454 22982 2471
rect 22889 2188 22961 2454
rect 15168 1473 15807 1476
rect 15168 1413 15822 1473
rect 16154 1430 16971 1642
rect 15168 1411 15728 1413
rect 15168 1359 15206 1411
rect 15258 1409 15728 1411
rect 15258 1359 15466 1409
rect 15168 1357 15466 1359
rect 15518 1361 15728 1409
rect 15780 1361 15822 1413
rect 15518 1357 15822 1361
rect 15168 1200 15822 1357
rect 15183 1197 15822 1200
rect 15185 1122 15547 1197
rect 15231 1115 15547 1122
rect 15231 706 15439 1115
rect 15696 1111 15813 1197
rect 16150 592 16967 804
rect 19733 690 19996 755
rect 19733 687 19925 690
rect 19733 635 19750 687
rect 19802 638 19925 687
rect 19977 638 19996 690
rect 19802 635 19996 638
rect 19733 618 19996 635
rect 20589 224 20684 565
rect 20889 224 20984 565
<< via1 >>
rect 19051 4833 19103 4885
rect 19257 4830 19309 4882
rect 19449 4817 19501 4869
rect 19637 4811 19689 4863
rect 19864 4822 19916 4874
rect 17209 3814 17261 3866
rect 23504 3860 23556 3912
rect 23646 3860 23698 3912
rect 23785 3860 23837 3912
rect 17224 3602 17276 3654
rect 17398 3602 17450 3654
rect 22823 3647 22875 3699
rect 22943 3647 22995 3699
rect 22899 2785 22951 2837
rect 23354 2785 23406 2837
rect 23479 2785 23531 2837
rect 23625 2785 23677 2837
rect 22899 2643 22951 2695
rect 22899 2471 22951 2523
rect 15206 1359 15258 1411
rect 15466 1357 15518 1409
rect 15728 1361 15780 1413
rect 19750 635 19802 687
rect 19925 638 19977 690
<< metal2 >>
rect 17169 5029 23406 5161
rect 17169 3911 17301 5029
rect 19003 4889 20046 4936
rect 19003 4833 19048 4889
rect 19104 4886 20046 4889
rect 19104 4833 19254 4886
rect 19003 4830 19254 4833
rect 19310 4878 20046 4886
rect 19310 4873 19861 4878
rect 19310 4830 19446 4873
rect 19003 4817 19446 4830
rect 19502 4867 19861 4873
rect 19502 4817 19634 4867
rect 19003 4811 19634 4817
rect 19690 4822 19861 4867
rect 19917 4822 20046 4878
rect 19690 4811 20046 4822
rect 19003 4549 20046 4811
rect 19910 4170 20035 4549
rect 19936 4147 20008 4170
rect 17167 3866 17301 3911
rect 17167 3814 17209 3866
rect 17261 3847 17301 3866
rect 23274 3927 23406 5029
rect 23481 3927 23860 3946
rect 23274 3912 23861 3927
rect 23274 3860 23504 3912
rect 23556 3860 23646 3912
rect 23698 3860 23785 3912
rect 23837 3860 23861 3912
rect 17261 3814 17300 3847
rect 17167 3694 17300 3814
rect 23274 3845 23861 3860
rect 22811 3739 23024 3741
rect 23274 3739 23406 3845
rect 23481 3825 23860 3845
rect 22811 3699 23406 3739
rect 17167 3654 17490 3694
rect 17167 3602 17224 3654
rect 17276 3602 17398 3654
rect 17450 3602 17490 3654
rect 22811 3647 22823 3699
rect 22875 3647 22943 3699
rect 22995 3647 23406 3699
rect 22811 3608 23406 3647
rect 22821 3607 23406 3608
rect 17167 3578 17490 3602
rect 22874 2847 22982 2860
rect 23311 2847 23695 2858
rect 22874 2837 23696 2847
rect 22874 2785 22899 2837
rect 22951 2785 23354 2837
rect 23406 2785 23479 2837
rect 23531 2785 23625 2837
rect 23677 2785 23696 2837
rect 22874 2775 23696 2785
rect 22874 2695 22982 2775
rect 23311 2764 23695 2775
rect 22874 2643 22899 2695
rect 22951 2643 22982 2695
rect 22874 2523 22982 2643
rect 22874 2471 22899 2523
rect 22951 2471 22982 2523
rect 22874 2454 22982 2471
rect 15659 1476 15849 1687
rect 15168 1413 15849 1476
rect 15168 1411 15728 1413
rect 15168 1359 15206 1411
rect 15258 1409 15728 1411
rect 15258 1359 15466 1409
rect 15168 1357 15466 1359
rect 15518 1361 15728 1409
rect 15780 1361 15849 1413
rect 15518 1357 15849 1361
rect 15168 1200 15849 1357
rect 15183 1197 15849 1200
rect 15659 163 15849 1197
rect 19733 699 19996 755
rect 20097 699 20192 712
rect 19733 690 20192 699
rect 19733 687 19925 690
rect 19733 635 19750 687
rect 19802 638 19925 687
rect 19977 638 20192 690
rect 19802 635 20192 638
rect 19733 630 20192 635
rect 19733 618 19996 630
rect 20097 163 20192 630
rect 15659 -27 20239 163
<< via2 >>
rect 19048 4885 19104 4889
rect 19048 4833 19051 4885
rect 19051 4833 19103 4885
rect 19103 4833 19104 4885
rect 19254 4882 19310 4886
rect 19254 4830 19257 4882
rect 19257 4830 19309 4882
rect 19309 4830 19310 4882
rect 19861 4874 19917 4878
rect 19446 4869 19502 4873
rect 19446 4817 19449 4869
rect 19449 4817 19501 4869
rect 19501 4817 19502 4869
rect 19634 4863 19690 4867
rect 19634 4811 19637 4863
rect 19637 4811 19689 4863
rect 19689 4811 19690 4863
rect 19861 4822 19864 4874
rect 19864 4822 19916 4874
rect 19916 4822 19917 4874
<< metal3 >>
rect 19008 4889 20046 4933
rect 19008 4833 19048 4889
rect 19104 4886 20046 4889
rect 19104 4833 19254 4886
rect 19008 4830 19254 4833
rect 19310 4878 20046 4886
rect 19310 4873 19861 4878
rect 19310 4830 19446 4873
rect 19008 4817 19446 4830
rect 19502 4867 19861 4873
rect 19502 4817 19634 4867
rect 19008 4811 19634 4817
rect 19690 4822 19861 4867
rect 19917 4822 20046 4878
rect 19690 4811 20046 4822
rect 19008 4726 20046 4811
rect 16603 4546 20046 4726
rect 6472 480 6581 654
rect 6436 357 6616 480
rect 16603 357 16783 4546
rect 6436 177 16783 357
use DFF_3_mag  DFF_3_mag_0
timestamp 1713185578
transform 1 0 21146 0 1 418
box -4189 -222 2082 4087
use VCO_C  VCO_C_0
timestamp 1713971361
transform 1 0 1330 0 1 36
box -1420 -36 14830 7134
<< labels >>
flabel metal1 s 23729 2805 23729 2805 0 FreeSans 2500 0 0 0 OUT
port 1 nsew
flabel metal1 s 23891 3883 23891 3883 0 FreeSans 2500 0 0 0 OUTB
port 2 nsew
flabel metal1 s 16348 4249 16348 4249 0 FreeSans 2500 0 0 0 VSS
port 3 nsew
flabel metal1 s 15330 802 15330 802 0 FreeSans 2500 0 0 0 VDD
port 4 nsew
flabel metal1 s 7087 7018 7087 7018 0 FreeSans 2500 0 0 0 VCTRL2
port 5 nsew
flabel metal1 s 6120 5786 6120 5786 0 FreeSans 2500 0 0 0 VCTRL
port 6 nsew
<< end >>
