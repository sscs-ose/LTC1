magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2845 -2095 2845 2095
<< psubdiff >>
rect -845 70 845 95
rect -845 -70 -822 70
rect 822 -70 845 70
rect -845 -95 845 -70
<< psubdiffcont >>
rect -822 -70 822 70
<< metal1 >>
rect -834 70 834 84
rect -834 -70 -822 70
rect 822 -70 834 70
rect -834 -84 834 -70
<< end >>
