* NGSPICE file created from nor_3_mag_flat.ext - technology: gf180mcuC

.subckt nor_3_mag_flat IN3 IN2 IN1 OUT VDD VSS
X0 a_720_997# IN2.t0 a_560_997# VDD.t0 pfet_03v3 ad=0.624p pd=2.92u as=0.624p ps=2.92u w=2.4u l=0.28u
X1 OUT IN3.t0 VSS.t6 VSS.t5 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X2 OUT IN1.t0 a_720_997# VDD.t1 pfet_03v3 ad=1.06p pd=5.68u as=0.624p ps=2.92u w=2.4u l=0.28u
X3 OUT IN1.t1 VSS.t1 VSS.t0 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X4 a_560_997# IN3.t1 VDD.t3 VDD.t2 pfet_03v3 ad=0.624p pd=2.92u as=1.06p ps=5.68u w=2.4u l=0.28u
X5 VSS IN2.t1 OUT.t1 VSS.t2 nfet_03v3 ad=86.8f pd=0.92u as=86.8f ps=0.92u w=0.22u l=0.28u
R0 IN2.n0 IN2.t0 40.7733
R1 IN2.n0 IN2.t1 27.7883
R2 IN2 IN2.n0 4.05105
R3 VDD.t0 VDD.t1 175.631
R4 VDD.n1 VDD.t2 153.678
R5 VDD.n1 VDD.t0 21.9544
R6 VDD VDD.t3 4.11425
R7 VDD VDD.n2 3.15126
R8 VDD.n2 VDD.n1 3.1505
R9 VDD.n2 VDD.n0 0.0401226
R10 IN3.n0 IN3.t1 40.7733
R11 IN3.n0 IN3.t0 25.1594
R12 IN3 IN3.n0 4.04735
R13 VSS.t2 VSS.t0 1278.69
R14 VSS.n2 VSS.t2 745.903
R15 VSS.n2 VSS.t5 532.788
R16 VSS VSS.t6 9.49031
R17 VSS.n1 VSS.n0 6.01414
R18 VSS.n1 VSS.t1 6.01414
R19 VSS.n5 VSS.n1 3.50163
R20 VSS.n5 VSS.n4 2.6005
R21 VSS.n4 VSS.n2 2.6005
R22 VSS.n4 VSS.n3 0.301575
R23 VSS VSS.n5 0.00352521
R24 OUT.n4 OUT.n3 9.28675
R25 OUT.n2 OUT.n1 6.01414
R26 OUT.n2 OUT.t1 6.01414
R27 OUT.n5 OUT.n0 3.87666
R28 OUT.n4 OUT.n2 3.74699
R29 OUT.n5 OUT.n4 0.0409348
R30 OUT OUT.n5 0.0239783
R31 IN1.n0 IN1.t0 40.4409
R32 IN1.n0 IN1.t1 29.9982
R33 IN1 IN1.n0 4.05968
C0 OUT a_720_997# 0.198f
C1 VDD a_560_997# 0.234f
C2 IN1 a_720_997# 0.0168f
C3 IN2 a_720_997# 8.64e-19
C4 OUT VDD 0.0708f
C5 IN1 VDD 0.125f
C6 IN2 VDD 0.115f
C7 IN3 VDD 0.146f
C8 VDD a_720_997# 0.0407f
C9 OUT a_560_997# 0.0132f
C10 IN2 a_560_997# 0.00365f
C11 IN3 a_560_997# 8.64e-19
C12 OUT IN1 0.201f
C13 OUT IN2 0.109f
C14 OUT IN3 0.00868f
C15 IN2 IN1 0.0964f
C16 IN2 IN3 0.0829f
C17 a_560_997# a_720_997# 0.186f
.ends

