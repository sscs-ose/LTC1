magic
tech gf180mcuC
magscale 1 10
timestamp 1693229188
<< psubdiff >>
rect 645 1399 4765 1415
rect 645 1259 679 1399
rect 889 1259 1029 1399
rect 1239 1259 1379 1399
rect 1589 1259 1729 1399
rect 1939 1259 2079 1399
rect 2289 1259 2429 1399
rect 2639 1259 2779 1399
rect 2989 1259 3129 1399
rect 3339 1259 3479 1399
rect 3689 1259 3829 1399
rect 4039 1259 4179 1399
rect 4389 1259 4529 1399
rect 4739 1259 4765 1399
rect 645 1205 4765 1259
rect 37 140 4717 181
rect 37 0 130 140
rect 340 0 480 140
rect 690 0 830 140
rect 1040 0 1180 140
rect 1390 0 1530 140
rect 1740 0 1880 140
rect 2090 0 2230 140
rect 2440 0 2580 140
rect 2790 0 2930 140
rect 3140 0 3280 140
rect 3490 0 3630 140
rect 3840 0 3980 140
rect 4190 0 4330 140
rect 4540 0 4717 140
rect 37 -60 4717 0
<< psubdiffcont >>
rect 679 1259 889 1399
rect 1029 1259 1239 1399
rect 1379 1259 1589 1399
rect 1729 1259 1939 1399
rect 2079 1259 2289 1399
rect 2429 1259 2639 1399
rect 2779 1259 2989 1399
rect 3129 1259 3339 1399
rect 3479 1259 3689 1399
rect 3829 1259 4039 1399
rect 4179 1259 4389 1399
rect 4529 1259 4739 1399
rect 130 0 340 140
rect 480 0 690 140
rect 830 0 1040 140
rect 1180 0 1390 140
rect 1530 0 1740 140
rect 1880 0 2090 140
rect 2230 0 2440 140
rect 2580 0 2790 140
rect 2930 0 3140 140
rect 3280 0 3490 140
rect 3630 0 3840 140
rect 3980 0 4190 140
rect 4330 0 4540 140
<< polysilicon >>
rect 112 1166 4872 1180
rect 112 1087 180 1166
rect 259 1087 4872 1166
rect 112 1073 4872 1087
rect 112 976 312 1073
rect 1024 976 1224 1073
rect 1328 976 1528 1073
rect 2240 976 2440 1073
rect 2544 976 2744 1073
rect 3456 976 3656 1073
rect 3760 976 3960 1073
rect 4672 976 4872 1073
rect -112 709 -25 729
rect -112 661 -92 709
rect -43 703 -25 709
rect 416 703 616 768
rect 720 703 920 768
rect 1632 703 1832 768
rect 1936 703 2136 768
rect 2848 703 3048 768
rect 3152 703 3352 768
rect 4064 703 4264 768
rect 4368 703 4568 768
rect -43 666 4872 703
rect -43 661 -25 666
rect -112 642 -25 661
rect 112 594 312 666
rect 1024 594 1224 666
rect 1328 594 1528 666
rect 2240 594 2440 666
rect 2544 594 2744 666
rect 3456 594 3656 666
rect 3760 594 3960 666
rect 4672 594 4872 666
rect 507 386 616 430
rect 147 324 265 327
rect 147 312 290 324
rect 147 247 188 312
rect 253 263 290 312
rect 416 263 616 386
rect 720 263 920 386
rect 1632 263 1832 386
rect 1936 263 2136 386
rect 2848 263 3048 386
rect 3152 263 3352 386
rect 4064 263 4264 386
rect 4368 263 4568 386
rect 253 247 4568 263
rect 147 230 4568 247
rect 182 226 4568 230
<< polycontact >>
rect 180 1087 259 1166
rect -92 661 -43 709
rect 188 247 253 312
<< metal1 >>
rect 4751 1415 4999 1437
rect 645 1409 5009 1415
rect 645 1408 4916 1409
rect 645 1399 4772 1408
rect 645 1259 679 1399
rect 889 1259 1029 1399
rect 1239 1259 1379 1399
rect 1589 1259 1729 1399
rect 1939 1259 2079 1399
rect 2289 1259 2429 1399
rect 2639 1259 2779 1399
rect 2989 1259 3129 1399
rect 3339 1259 3479 1399
rect 3689 1259 3829 1399
rect 4039 1259 4179 1399
rect 4389 1259 4529 1399
rect 4739 1348 4772 1399
rect 4832 1348 4916 1408
rect 4739 1347 4916 1348
rect 4978 1347 5009 1409
rect 4739 1295 5009 1347
rect 4739 1259 4765 1295
rect 645 1233 4765 1259
rect 4827 1294 5009 1295
rect 4827 1234 4917 1294
rect 4977 1234 5009 1294
rect 4827 1233 5009 1234
rect 645 1205 5009 1233
rect 171 1166 268 1175
rect 171 1087 180 1166
rect 259 1087 268 1166
rect 171 1078 268 1087
rect 645 921 691 1205
rect 1861 928 1907 1205
rect 3077 930 3123 1205
rect 4293 930 4339 1205
rect 325 906 403 917
rect 325 838 333 906
rect 393 838 403 906
rect 325 829 403 838
rect 939 910 1017 922
rect 939 844 949 910
rect 1006 844 1017 910
rect 939 834 1017 844
rect 1538 906 1616 918
rect 1538 840 1548 906
rect 1605 840 1616 906
rect 1538 830 1616 840
rect 2145 908 2223 920
rect 2145 842 2155 908
rect 2212 842 2223 908
rect 2145 832 2223 842
rect 2755 908 2833 920
rect 2755 842 2765 908
rect 2822 842 2833 908
rect 2755 832 2833 842
rect 3361 906 3439 918
rect 3361 840 3371 906
rect 3428 840 3439 906
rect 3361 830 3439 840
rect 3969 906 4047 918
rect 3969 840 3979 906
rect 4036 840 4047 906
rect 3969 830 4047 840
rect 4580 910 4658 922
rect 4580 844 4590 910
rect 4647 844 4658 910
rect 4580 834 4658 844
rect 37 755 83 815
rect 1253 755 1299 814
rect 2469 755 2515 814
rect 3685 755 3731 814
rect 4901 755 4947 814
rect -112 709 -25 729
rect -112 661 -92 709
rect -43 661 -25 709
rect 37 675 5231 755
rect -112 642 -25 661
rect 645 548 691 675
rect 1861 548 1907 675
rect 3077 548 3123 675
rect 4293 548 4339 675
rect 316 526 394 538
rect 316 460 326 526
rect 383 460 394 526
rect 316 450 394 460
rect 933 529 1011 541
rect 933 463 943 529
rect 1000 463 1011 529
rect 933 453 1011 463
rect 1537 528 1615 540
rect 1537 462 1547 528
rect 1604 462 1615 528
rect 1537 452 1615 462
rect 2146 525 2224 537
rect 2146 459 2156 525
rect 2213 459 2224 525
rect 2146 449 2224 459
rect 2755 521 2833 533
rect 2755 455 2765 521
rect 2822 455 2833 521
rect 2755 445 2833 455
rect 3368 521 3446 533
rect 3368 455 3378 521
rect 3435 455 3446 521
rect 3368 445 3446 455
rect 3969 527 4047 539
rect 3969 461 3979 527
rect 4036 461 4047 527
rect 4582 537 4660 549
rect 4582 471 4592 537
rect 4649 471 4660 537
rect 4582 461 4660 471
rect 3969 451 4047 461
rect 37 181 83 432
rect 147 312 265 327
rect 147 247 188 312
rect 253 247 265 312
rect 147 230 265 247
rect 1253 181 1299 432
rect 2469 181 2515 432
rect 3685 181 3731 432
rect 4901 181 4947 432
rect 37 170 4947 181
rect 37 166 4847 170
rect 37 140 4718 166
rect 37 0 130 140
rect 340 0 480 140
rect 690 0 830 140
rect 1040 0 1180 140
rect 1390 0 1530 140
rect 1740 0 1880 140
rect 2090 0 2230 140
rect 2440 0 2580 140
rect 2790 0 2930 140
rect 3140 0 3280 140
rect 3490 0 3630 140
rect 3840 0 3980 140
rect 4190 0 4330 140
rect 4540 106 4718 140
rect 4778 108 4847 166
rect 4909 108 4947 170
rect 4778 106 4947 108
rect 4540 56 4947 106
rect 4540 49 4848 56
rect 4540 0 4717 49
rect 37 -13 4717 0
rect 4779 -4 4848 49
rect 4908 -4 4947 56
rect 4779 -13 4947 -4
rect 37 -60 4947 -13
<< via1 >>
rect 4772 1348 4832 1408
rect 4916 1347 4978 1409
rect 4765 1233 4827 1295
rect 4917 1234 4977 1294
rect 190 1098 246 1154
rect 333 838 393 906
rect 949 844 1006 910
rect 1548 840 1605 906
rect 2155 842 2212 908
rect 2765 842 2822 908
rect 3371 840 3428 906
rect 3979 840 4036 906
rect 4590 844 4647 910
rect 326 460 383 526
rect 943 463 1000 529
rect 1547 462 1604 528
rect 2156 459 2213 525
rect 2765 455 2822 521
rect 3378 455 3435 521
rect 3979 461 4036 527
rect 4592 471 4649 537
rect 191 249 245 303
rect 4718 106 4778 166
rect 4847 108 4909 170
rect 4717 -13 4779 49
rect 4848 -4 4908 56
<< metal2 >>
rect 4751 1409 4999 1437
rect 4751 1408 4916 1409
rect 4751 1348 4772 1408
rect 4832 1348 4916 1408
rect 4751 1347 4916 1348
rect 4978 1347 4999 1409
rect 4751 1295 4999 1347
rect 4751 1233 4765 1295
rect 4827 1294 4999 1295
rect 4827 1234 4917 1294
rect 4977 1234 4999 1294
rect 4827 1233 4999 1234
rect 4751 1216 4999 1233
rect 165 1167 279 1181
rect 152 1154 279 1167
rect 152 1098 190 1154
rect 246 1098 279 1154
rect 152 1070 279 1098
rect 152 327 246 1070
rect 325 906 403 917
rect 325 838 333 906
rect 393 838 403 906
rect 325 829 403 838
rect 939 910 1017 922
rect 939 844 949 910
rect 1006 844 1017 910
rect 939 834 1017 844
rect 1538 906 1616 918
rect 1538 840 1548 906
rect 1605 840 1616 906
rect 331 674 393 829
rect 944 674 1006 834
rect 1538 830 1616 840
rect 2145 908 2223 920
rect 2145 842 2155 908
rect 2212 842 2223 908
rect 2145 832 2223 842
rect 2755 908 2833 920
rect 2755 842 2765 908
rect 2822 842 2833 908
rect 2755 832 2833 842
rect 3361 906 3439 918
rect 3361 840 3371 906
rect 3428 840 3439 906
rect 1546 674 1608 830
rect 2157 674 2219 832
rect 2762 674 2824 832
rect 3361 830 3439 840
rect 3969 906 4047 918
rect 3969 840 3979 906
rect 4036 840 4047 906
rect 3969 830 4047 840
rect 4580 910 4658 922
rect 4580 844 4590 910
rect 4647 844 4658 910
rect 4580 834 4658 844
rect 3374 674 3436 830
rect 3980 674 4042 830
rect 4588 674 4650 834
rect 331 612 4650 674
rect 331 538 393 612
rect 944 541 1006 612
rect 316 526 394 538
rect 316 460 326 526
rect 383 460 394 526
rect 316 450 394 460
rect 933 529 1011 541
rect 1546 540 1608 612
rect 933 463 943 529
rect 1000 463 1011 529
rect 933 453 1011 463
rect 1537 528 1615 540
rect 2157 537 2219 612
rect 1537 462 1547 528
rect 1604 462 1615 528
rect 1537 452 1615 462
rect 2146 525 2224 537
rect 2762 533 2824 612
rect 3374 533 3436 612
rect 3980 539 4042 612
rect 4588 549 4650 612
rect 2146 459 2156 525
rect 2213 459 2224 525
rect 2146 449 2224 459
rect 2755 521 2833 533
rect 2755 455 2765 521
rect 2822 455 2833 521
rect 2755 445 2833 455
rect 3368 521 3446 533
rect 3368 455 3378 521
rect 3435 455 3446 521
rect 3368 445 3446 455
rect 3969 527 4047 539
rect 3969 461 3979 527
rect 4036 461 4047 527
rect 4582 537 4660 549
rect 4582 471 4592 537
rect 4649 471 4660 537
rect 4582 461 4660 471
rect 3969 451 4047 461
rect 147 303 265 327
rect 147 249 191 303
rect 245 249 265 303
rect 147 230 265 249
rect 4765 179 4909 1216
rect 4698 170 4937 179
rect 4698 166 4847 170
rect 4698 106 4718 166
rect 4778 108 4847 166
rect 4909 108 4937 170
rect 4778 106 4937 108
rect 4698 56 4937 106
rect 4698 49 4848 56
rect 4698 -13 4717 49
rect 4779 -4 4848 49
rect 4908 -4 4937 56
rect 4779 -13 4937 -4
rect 4698 -48 4937 -13
use nmos_3p3_GJ7FB7  nmos_3p3_GJ7FB7_0
timestamp 1693226830
transform 1 0 2492 0 1 872
box -2492 -128 2492 128
use nmos_3p3_GJ7FB7  nmos_3p3_GJ7FB7_1
timestamp 1693226830
transform 1 0 2492 0 1 490
box -2492 -128 2492 128
<< labels >>
flabel psubdiffcont 2534 1326 2534 1326 0 FreeSans 640 0 0 0 VSS
port 0 nsew
flabel metal1 5166 721 5166 721 0 FreeSans 640 0 0 0 OUT
port 1 nsew
flabel polycontact -72 694 -72 694 0 FreeSans 640 0 0 0 IM
port 2 nsew
flabel via1 214 1126 214 1126 0 FreeSans 640 0 0 0 IM_T
port 3 nsew
<< end >>
