** sch_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/TB_TOP_MUX_F6_sch.sch
**.subckt TB_TOP_MUX_F6_sch
V1 VSS GND 0
.save i(v1)
V3 VCTRL2 VSS 3.3
.save i(v3)
V4 VCTRL_IN VSS 0.6
.save i(v4)
V6 F_IN VSS pulse(0 3.3 200n 100p 100p 50n 100n)
.save i(v6)
I4 VDD ITAIL 100u
V8 S1 VSS 0
.save i(v8)
V9 S2 VSS 0
.save i(v9)
V10 S3 VSS 0
.save i(v10)
V11 S4 VSS 0
.save i(v11)
V12 S6 VSS 0
.save i(v12)
V13 DN_INPUT VSS pulse(0 3.3 10n 100p 100p 500n 1000n)
.save i(v13)
V14 UP_INPUT VSS pulse(0 3.3 0 100p 100p 500n 1000n)
.save i(v14)
V15 VDD_TEST VSS 3.3
.save i(v15)
C1 LF_OFFCHIP VSS 11.27p m=1
R1 LF_OFFCHIP net1 74k m=1
C2 net1 VSS 239p m=1
V16 S5 VSS 0
.save i(v16)
V17 D0 VSS 0
.save i(v17)
V18 D1 VSS 3.3
.save i(v18)
V19 D2 VSS 0
.save i(v19)
V20 D3 VSS 0
.save i(v20)
V21 D4 VSS 0
.save i(v21)
V22 D5 VSS 3.3
.save i(v22)
V23 D6 VSS 3.3
.save i(v23)
V29 D12 VSS 0
.save i(v29)
V30 D13 VSS 0
.save i(v30)
V31 D14 VSS 0
.save i(v31)
V32 D15 VSS 3.3
.save i(v32)
V33 D16 VSS 0
.save i(v33)
V2 S7 VSS 0
.save i(v2)
V5 VDD VSS pwl(0 0 0.05US 0 0.050001US 3.3)
.save i(v5)
V7 D7 VSS 0
.save i(v7)
V34 D8 VSS 0
.save i(v34)
V35 D9 VSS 0
.save i(v35)
V36 D10 VSS 3.3
.save i(v36)
V37 D11 VSS 0
.save i(v37)
V24 DIV_OUT2 VSS pulse(0 3.3 700n 100p 100p 500n 1000n)
.save i(v24)
V25 D26G GND 0
.save i(v25)
V26 D27G GND 0
.save i(v26)
V27 D17G GND 0
.save i(v27)
x1 VDD_TEST D12 D0 UP_INPUT D13 D1 DN_INPUT VSS D14 D2 PRE_SCALAR UP_OUT D15 D3 F_IN DN_OUT D16 D4
+ ITAIL DIV_OUT D5 S1 S6 D6 VCTRL_IN D7 VCTRL2 S2 D8 S3 OUT D9 OUTB S4 LF_OFFCHIP D10 S5 S7 D11 OUT1
+ DIV_OUT2 D27G D26G D17G D16G VDD PLL_TOP5
V28 D16G GND 0
.save i(v28)
**** begin user architecture code


.include pex_A_MUX.spice
.include pex_VCO_DFF_C.spice
.include Tappered-Buffer_1_pex.spice
.include pex_PFD_T2.spice
.include pex_CP.spice
.include Res_74k_pex.spice
.include pex_cap_11p.spice
.include pex_cap_240p.spice
.include pex_PLL_TOP_MUX_6.spice
.include pex_7b_divider_magic.spice
*.include pex_PLL_TOP_MUX_2.spice
*.include Tappered-Buffer_1_pex.spice
*.option RSHUNT=1e18
**.option ABSTOL=1e-12
**.option VNTOL=1e-12
**.option CHGTOL=1e-14
**.option RELTOL=1e-5
.option gmin=1e-15
**.option trtol=1
**.OPTION ITL4=500
.control
save x1.vco_dff_c_0.vctrl.t19  x1.pre_scalar.n0  pre_scalar  x1.vss.t6260  x1.vdd.n7823
+  x1.vctrl_in.t6  x1.vctrl2.t62  x1.vco_dff_c_0.vco_c_0.outb.t53  x1.vco_dff_c_0.vco_c_0.inv_2_5.in.n34
+  x1.vco_dff_c_0.vco_c_0.inv_2_3.out.n2  x1.vco_dff_c_0.vco_c_0.inv_2_2.in.n30  x1.vco_dff_c_0.vco_c_0.inv_2_0.in.n51
+  x1.vco_dff_c_0.outb.t31  x1.vco_dff_c_0.out.t10  x1.up_out.t60  x1.up_input.n12  x1.up1.n10  x1.up.n28  x1.dn
+  x1.a_mux_6.in1.n194  x1.a_mux_5.in1.t163  x1.a_mux_2.out.n14  x1.a_mux_1.out  x1.a_mux_6.out
+  x1.7b_divider_magic_2.p2_gen_magic_0.dff_magic_0.tg_magic_3.out  x1.7b_divider_magic_2.p2_gen_magic_0.dff_magic_0.tg_magic_3.clk
+  x1.7b_divider_magic_2.p2_gen_magic_0.dff_magic_0.tg_magic_2.in.n10  x1.7b_divider_magic_2.p2.t16  x1.7b_divider_magic_2.out1.t8
+  x1.7b_divider_magic_2.divide_by_2_1.tg_magic_3.out  x1.7b_divider_magic_2.divide_by_2_1.tg_magic_3.clk
+  x1.7b_divider_magic_1.p2_gen_magic_0.dff_magic_0.tg_magic_1.in.n19  x1.7b_divider_magic_1.ld  x1.7b_divider_magic_1.divide_by_2_1.tg_magic_2.in.n14
+  x1.7b_divider_magic_1.divide_by_2_0.tg_magic_3.out  x1.7b_divider_magic_1.divide_by_2_0.tg_magic_3.in  x1.7b_divider_magic_0.out1
+  x1.7b_divider_magic_0.ld.n38  x1.vctrl_obv  x1.a_mux_6.out.n27  out1  out  outb  net1  lf_offchip  itail1  itail  f_in  dn_out
+  up_out  dn_input  div_out
*set ngbehavior=hsa
*set ng_nomodcheck
tran 500n 20u
set appendwrite
write TB_TOP_MUX_F6_sch.raw
.endc



.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice res_typical
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice cap_mim
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice moscap_typical
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice mimcap_typical

**** end user architecture code
**.ends

* expanding   symbol:  PLL_TOP5.sym # of pins=46
** sym_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/PLL_TOP5.sym
** sch_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/PLL_TOP5.sch
.subckt PLL_TOP5 VDD_TEST D12 D0 UP_INPUT D13 D1 DN_INPUT VSS D14 D2 PRE_SCALAR UP_OUT D15 D3 F_IN
+ DN_OUT D16 D4 ITAIL DIV_OUT D5 S1 S6 D6 VCTRL_IN D7 VCTRL2 S2 D8 S3 OUT D9 OUTB S4 LF_OFFCHIP D10 S5 S7
+ D11 OUT1 DIV_OUT2 D27G D26G D17G D16G VDD
*.ipin UP_INPUT
*.ipin DN_INPUT
*.opin UP_OUT
*.opin DN_OUT
*.ipin ITAIL
*.ipin VCTRL2
*.opin OUT
*.iopin OUTB
*.iopin VDD
*.iopin VSS
*.opin PRE_SCALAR
*.ipin F_IN
*.opin DIV_OUT
*.ipin S1
*.ipin S6
*.ipin S2
*.ipin S3
*.ipin VCTRL_IN
*.ipin S4
*.ipin S5
*.ipin LF_OFFCHIP
*.ipin D0
*.ipin D1
*.ipin D2
*.ipin D3
*.ipin D4
*.ipin D5
*.ipin D6
*.ipin D7
*.ipin D8
*.ipin D9
*.ipin D10
*.ipin D11
*.ipin D12
*.ipin D13
*.ipin D14
*.ipin D15
*.ipin D16
*.opin OUT1
*.ipin S7
*.iopin VDD_TEST
*.ipin DIV_OUT2
*.ipin D27G
*.ipin D26G
*.ipin D17G
*.ipin D16G
x17 VDD LD1 D17G Q11 D16G Q12 D16 D15 Q13 Q14 D14 D13 Q15 D12 Q16 Q17 OUT_D VSS OUT11 P12 7b_divider
x18 VDD LD2 D27G Q21 D26G Q22 D11 D10 Q23 Q24 D9 D8 Q25 D7 Q26 Q27 F_IN VSS net5 P22
+ pex_7b_divider_magic
x13 VSS VDD_TEST PRE_SCALAR net5 Tappered-Buffer_1_pex
x2 VDD VSS net5 F_IN S1 net8 A_MUX_pex
x3 VDD VSS OUT01 DIV_OUT2 S6 net9 A_MUX_pex
x4 VDD VSS net2 UP_INPUT S2 UP A_MUX_pex
x5 VDD VSS net3 DN_INPUT S3 DN A_MUX_pex
x6 VDD VSS net7 VCTRL_IN S4 VCTRL_OBV A_MUX_pex
x12 VDD VSS net6 LF_OFFCHIP S5 net7 A_MUX_pex
x14 VSS VDD_TEST UP_OUT UP Tappered-Buffer_1_pex
x15 VSS VDD_TEST OUT net1 Tappered-Buffer_1_pex
x19 VSS VDD_TEST OUTB net10 Tappered-Buffer_1_pex
x20 VSS VDD_TEST OUT_D net1 Tappered-Buffer_1_pex
x21 VSS VDD_TEST DIV_OUT OUT01 Tappered-Buffer_1_pex
x22 VSS VDD_TEST OUT1 OUT11 Tappered-Buffer_1_pex
x23 VSS VDD_TEST DN_OUT DN Tappered-Buffer_1_pex
x16 VDD LD0 D6 Q01 D5 Q02 D4 D3 Q03 Q04 D2 D1 Q05 D0 Q06 Q07 IN_DIV VSS OUT01 P02
+ pex_7b_divider_magic
x1 net2 VDD VSS net8 net9 net3 PFD_ver_2_pex
x24 VDD VSS OUT_D F_IN S7 IN_DIV A_MUX_pex
x9 net6 VDD net4 Res_74k_pex
x10 net6 VSS cap_11p_pex
x11 net4 VSS cap_240p_pex
x8 VDD ITAIL_SINK ITAIL_SRC net7 DN UP VSS loop_filter_V1_pex
x7 VDD VSS VCTRL_OBV VCTRL2 net1 net10 pex_VCO_DFF_C
x25 VDD ITAIL ITAIL_SRC ITAIL_SINK VSS Current_Mirror_Top_s
.ends


* expanding   symbol:  7b_divider.sym # of pins=20
** sym_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/7b_divider.sym
** sch_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/7b_divider.sch
.subckt 7b_divider VDD LD D2_7 Q1 D2_6 Q2 D2_5 D2_4 Q3 Q4 D2_3 D2_2 Q5 D2_1 Q6 Q7 CLK VSS OUT1 P2
*.iopin VDD
*.iopin VSS
*.ipin D2_1
*.ipin CLK
*.ipin D2_2
*.ipin D2_3
*.ipin D2_4
*.ipin D2_5
*.ipin D2_6
*.ipin D2_7
*.opin LD
*.opin Q1
*.opin Q2
*.opin Q3
*.opin Q4
*.opin Q5
*.opin Q6
*.opin Q7
*.opin P2
*.opin OUT1
x4 VDD Q2 b D2_3 VSS XNOR
x5 VDD Q1 a D2_2 VSS XNOR
x6 VDD Q3 c D2_4 VSS XNOR
x7 VDD net1 a b c VSS 3_inp_AND
x2 VDD Q4 d D2_5 VSS XNOR
x3 VDD Q5 e D2_6 VSS XNOR
x9 VDD Q6 f D2_7 VSS XNOR
x10 VDD Q7 g D2_1 VSS XNOR
x15 VDD net4 net1 net2 net3 VSS 3_inp_AND
x16 VDD P0 P2 net5 VSS OR
x17 net5 VDD OUT3 VSS div_by_2
x1 LD VDD Q6 Q4 Q2 Q5 Q1 Q3 Q7 D2_7 D2_6 D2_3 D2_5 D2_2 D2_4 D2_1 CLK VSS 7b_counter_new
x11 VDD net2 d e VSS AND
x12 VDD net3 f g VSS AND
x8 CLK VDD LD P0 VSS DFF
x14 VDD Q2 j2 D2_3 VSS XNOR
x18 VDD Q1 j1 D2_2 VSS XNOR
x19 VDD Q3 j3 D2_4 VSS XNOR
x20 VDD Q4 j4 D2_5 VSS XNOR
x21 VDD Q5 j5 D2_6 VSS XNOR
x22 VDD Q6 j6 D2_7 VSS XNOR
x23 VDD Q7 j7 D2_1B VSS XNOR
x24 VDD D2_1 D2_1B VSS inverter
x25 VDD net6 j1 j2 j3 VSS 3_inp_AND
x26 VDD net9 net6 net7 net8 VSS 3_inp_AND
x27 VDD net7 j4 j5 VSS AND
x28 VDD net8 j6 j7 VSS AND
x29 CLK VDD net9 P3 VSS ned_DFF
x30 VDD P0 P3 net10 VSS OR
x31 net10 VDD OUT2 VSS div_by_2
x32 VDD D2_1 OUT3 OUT1 VSS OUT2 MUX
x13 CLK VDD net4 P2 VSS DFF
.ends


* expanding   symbol:  Current_Mirror_Top_s.sym # of pins=5
** sym_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/Current_Mirror_Top_s.sym
** sch_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/Current_Mirror_Top_s.sch
.subckt Current_Mirror_Top_s VDD ITAIL ITAIL_SRC ITAIL_SINK VSS
*.ipin ITAIL
*.iopin VDD
*.iopin VSS
*.opin ITAIL_SRC
*.opin ITAIL_SINK
XM1 net2 ITAIL net1 VSS nfet_03v3 L=0.5u W=20u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 net1 net5 VSS VSS nfet_03v3 L=0.5u W=20u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM7 net2 net2 net3 VDD pfet_03v3 L=0.5u W=20u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM8 net3 net3 VDD VDD pfet_03v3 L=0.5u W=20u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM9 G_sink_up net2 net4 VDD pfet_03v3 L=0.5u W=4u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM10 net4 net3 VDD VDD pfet_03v3 L=0.5u W=4u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM11 G_sink_up G_sink_up G_sink_dn VSS nfet_03v3 L=0.5u W=4.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u'
+ as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)'
+ nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM12 G_sink_dn G_sink_dn VSS VSS nfet_03v3 L=0.5u W=4.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 ITAIL ITAIL net5 VSS nfet_03v3 L=0.5u W=20u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 net5 net5 VSS VSS nfet_03v3 L=0.5u W=20u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM5 G_source_dn G_sink_up net6 VSS nfet_03v3 L=0.5u W=4.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM6 net6 G_sink_dn VSS VSS nfet_03v3 L=0.5u W=4.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM13 G_source_dn G_source_dn G_source_up VDD pfet_03v3 L=0.5u W=4.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u'
+ as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)'
+ nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM14 G_source_up G_source_up VDD VDD pfet_03v3 L=0.5u W=4.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM15 ITAIL_SINK G_sink_up net7 VSS nfet_03v3 L=0.5u W=4.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM16 net7 G_sink_dn VSS VSS nfet_03v3 L=0.5u W=4.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM17 ITAIL_SRC G_source_dn net8 VDD pfet_03v3 L=0.5u W=4.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM18 net8 G_source_up VDD VDD pfet_03v3 L=0.5u W=4.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  XNOR.sym # of pins=5
** sym_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/XNOR.sym
** sch_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/XNOR.sch
.subckt XNOR VDD A OUT B VSS
*.iopin VDD
*.iopin VSS
*.ipin A
*.ipin B
*.opin OUT
XM1 OUT A net3 VSS nfet_03v3 L=0.56u W=1.12u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 net1 A VDD VDD pfet_03v3 L=0.56u W=2.24u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 net2 A_bar VDD VDD pfet_03v3 L=0.56u W=2.24u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 OUT B net1 VDD pfet_03v3 L=0.56u W=2.24u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM5 OUT B_bar net2 VDD pfet_03v3 L=0.56u W=2.24u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM6 OUT A_bar net4 VSS nfet_03v3 L=0.56u W=1.12u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM7 net3 B_bar VSS VSS nfet_03v3 L=0.56u W=1.12u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM8 net4 B VSS VSS nfet_03v3 L=0.56u W=1.12u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
x1 VDD A A_bar VSS inverter_1
x2 VDD B B_bar VSS inverter_1
.ends


* expanding   symbol:  3_inp_AND.sym # of pins=6
** sym_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/3_inp_AND.sym
** sch_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/3_inp_AND.sch
.subckt 3_inp_AND VDD VOUT A B C VSS
*.iopin VSS
*.iopin VDD
*.ipin A
*.ipin B
*.ipin C
*.opin VOUT
XM1 net3 A net1 VSS nfet_03v3 L=0.56u W=3.36u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 net3 C VDD VDD pfet_03v3 L=0.56u W=2.24u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 net1 B net2 VSS nfet_03v3 L=0.56u W=3.36u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 net2 C VSS VSS nfet_03v3 L=0.56u W=3.36u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM5 net3 B VDD VDD pfet_03v3 L=0.56u W=2.24u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM6 net3 A VDD VDD pfet_03v3 L=0.56u W=2.24u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM7 VOUT net3 VDD VDD pfet_03v3 L=0.56u W=2.24u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM8 VOUT net3 VSS VSS nfet_03v3 L=0.56u W=1.12u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM9 VOUT VOUT VOUT VDD pfet_03v3 L=0.56u W=1.12u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM10 VDD VDD VDD VDD pfet_03v3 L=0.56u W=1.12u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  OR.sym # of pins=5
** sym_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/OR.sym
** sch_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/OR.sch
.subckt OR VDD A B VOUT VSS
*.iopin VSS
*.iopin VDD
*.ipin A
*.ipin B
*.opin VOUT
XM1 net1 A VSS VSS nfet_03v3 L=0.56u W=1.12u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 net1 B net2 VDD pfet_03v3 L=0.56u W=4.48u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 net1 B VSS VSS nfet_03v3 L=0.56u W=1.12u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM6 net2 A VDD VDD pfet_03v3 L=0.56u W=4.48u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 VOUT net1 VDD VDD pfet_03v3 L=0.56u W=2.24u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM5 VOUT net1 VSS VSS nfet_03v3 L=0.56u W=1.12u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  div_by_2.sym # of pins=4
** sym_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/div_by_2.sym
** sch_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/div_by_2.sch
.subckt div_by_2 CLK VDD Q VSS
*.iopin VDD
*.iopin VSS
*.opin Q
*.ipin CLK
x1 VDD CLKB VSS net2 net1 tg
x3 VDD CLK VSS net2 net5 tg
x4 VDD CLK VSS net1 net3 tg
x5 VDD CLKB VSS net1 net4 tg
x2 VDD net2 net3 VSS inverter
x6 VDD net1 Q VSS inverter
x7 VDD Q net4 VSS inverter
x8 VDD net3 net5 VSS inverter
x9 VDD CLK CLKB VSS inverter
.ends


* expanding   symbol:  7b_counter_new.sym # of pins=18
** sym_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/7b_counter_new.sym
** sch_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/7b_counter_new.sch
.subckt 7b_counter_new LD VDD Q6 Q4 Q2 Q5 Q1 Q3 Q7 D2_7 D2_6 D2_3 D2_5 D2_2 D2_4 D2_1 G-CLK VSS
*.iopin VDD
*.iopin VSS
*.opin Q3
*.opin Q1
*.ipin D2_1
*.ipin D2_2
*.ipin D2_3
*.ipin G-CLK
*.opin Q2
*.opin LD
*.ipin D2_4
*.opin Q4
*.ipin D2_5
*.opin Q5
*.opin Q6
*.ipin D2_6
*.opin Q7
*.ipin D2_7
x6 VDD net3 net2 net1 VSS NAND
x9 VDD Q1 Q2 Q3 net9 VSS 3_inp_NOR
x7 G-CLK VDD net3 net2 VSS DFF
x8 VDD net2 LD VSS inverter
x1 VDD LD3 D2_1 Q1 a a VSS G-CLK G-CLK MOD_DFF_latest
x3 VDD LD3 D2_2 Q2 b b VSS Q1 G-CLK MOD_DFF_latest
x4 VDD LD1 D2_3 Q3 c c VSS Q2 G-CLK MOD_DFF_latest
x2 VDD LD1 D2_4 Q4 d d VSS Q3 G-CLK MOD_DFF_latest
x10 VDD LD2 D2_5 Q5 e e VSS Q4 G-CLK MOD_DFF_latest
x11 VDD LD1 D2_6 Q6 f f VSS Q5 G-CLK MOD_DFF_latest
x12 VDD LD2 D2_7 Q7 g g VSS Q6 G-CLK MOD_DFF_latest
x5 VDD net1 net5 net4 net9 VSS 3_inp_AND
x13 VDD Q4 Q5 net5 VSS NOR
x14 VDD Q6 Q7 net4 VSS NOR
XM4 net6 LD VDD VDD pfet_03v3 L=0.56u W=6.72u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM5 net6 LD VSS VSS nfet_03v3 L=0.56u W=3.36u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM1 LD1 net6 VSS VSS nfet_03v3 L=0.56u W=3.36u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 LD1 net6 VDD VDD pfet_03v3 L=0.56u W=6.72u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 net7 LD VSS VSS nfet_03v3 L=0.56u W=3.36u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM6 net7 LD VDD VDD pfet_03v3 L=0.56u W=6.72u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM7 LD2 net7 VDD VDD pfet_03v3 L=0.56u W=6.72u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM8 net8 LD VDD VDD pfet_03v3 L=0.56u W=6.72u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM9 LD3 net8 VDD VDD pfet_03v3 L=0.56u W=6.72u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM10 LD2 net7 VSS VSS nfet_03v3 L=0.56u W=3.36u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM11 net8 LD VSS VSS nfet_03v3 L=0.56u W=3.36u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM12 LD3 net8 VSS VSS nfet_03v3 L=0.56u W=3.36u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  AND.sym # of pins=5
** sym_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/AND.sym
** sch_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/AND.sch
.subckt AND VDD VOUT A B VSS
*.iopin VDD
*.iopin VSS
*.ipin A
*.ipin B
*.opin VOUT
XM1 net1 A net2 VSS nfet_03v3 L=0.56u W=2.24u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 net1 A VDD VDD pfet_03v3 L=0.56u W=2.24u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 net1 B VDD VDD pfet_03v3 L=0.56u W=2.24u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 net2 B VSS VSS nfet_03v3 L=0.56u W=2.24u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM5 VOUT net1 VDD VDD pfet_03v3 L=0.56u W=2.24u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM6 VOUT net1 VSS VSS nfet_03v3 L=0.56u W=1.12u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  DFF.sym # of pins=5
** sym_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/DFF.sym
** sch_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/DFF.sch
.subckt DFF CLK VDD D Q VSS
*.ipin D
*.iopin VDD
*.iopin VSS
*.opin Q
*.ipin CLK
x2 VDD net1 net2 VSS inverter
x6 VDD net3 Q VSS inverter
x7 VDD Q net4 VSS inverter
x8 VDD net2 net5 VSS inverter
x9 VDD CLK CLKB VSS inverter
x1 VDD CLKB VSS net1 D tg
x3 VDD CLK VSS net3 net2 tg
x4 VDD CLK VSS net1 net5 tg
x5 VDD CLKB VSS net3 net4 tg
.ends


* expanding   symbol:  inverter.sym # of pins=4
** sym_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/inverter.sym
** sch_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/inverter.sch
.subckt inverter VDD VIN VOUT VSS
*.iopin VDD
*.ipin VIN
*.opin VOUT
*.iopin VSS
XM4 VOUT VIN VDD VDD pfet_03v3 L=0.56u W=4.48u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM5 VOUT VIN VSS VSS nfet_03v3 L=0.56u W=2.24u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  ned_DFF.sym # of pins=5
** sym_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/ned_DFF.sym
** sch_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/ned_DFF.sch
.subckt ned_DFF CLK VDD D Q VSS
*.ipin D
*.iopin VDD
*.iopin VSS
*.opin Q
*.ipin CLK
x1 VDD CLK VSS net1 D tg
x3 VDD CLKB VSS net3 net2 tg
x4 VDD CLKB VSS net1 net5 tg
x5 VDD CLK VSS net3 net4 tg
x2 VDD CLK CLKB VSS inverter
x6 VDD net1 net2 VSS inverter
x7 VDD net2 net5 VSS inverter
x8 VDD Q net4 VSS inverter
x9 VDD net3 Q VSS inverter
.ends


* expanding   symbol:  MUX.sym # of pins=6
** sym_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/MUX.sym
** sch_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/MUX.sch
.subckt MUX VDD SEL IN1 VOUT VSS IN2
*.ipin SEL
*.ipin IN1
*.ipin IN2
*.opin VOUT
*.iopin VDD
*.iopin VSS
x2 VDD net3 net1 IN1 VSS AND
x3 VDD net2 SEL IN2 VSS AND
XM4 net1 SEL VDD VDD pfet_03v3 L=0.56u W=6.72u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM5 net1 SEL VSS VSS nfet_03v3 L=0.56u W=3.36u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
x1 VDD net3 net2 VOUT VSS OR
.ends


* expanding   symbol:  inverter_1.sym # of pins=4
** sym_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/inverter_1.sym
** sch_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/inverter_1.sch
.subckt inverter_1 VDD VIN VOUT VSS
*.iopin VDD
*.ipin VIN
*.opin VOUT
*.iopin VSS
XM4 VOUT VIN VDD VDD pfet_03v3 L=0.56u W=4.48u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM5 VOUT VIN VSS VSS nfet_03v3 L=0.56u W=2.24u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  tg.sym # of pins=5
** sym_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/tg.sym
** sch_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/tg.sch
.subckt tg VDD CLK VSS OUT IN
*.iopin VDD
*.iopin VSS
*.ipin CLK
*.ipin IN
*.opin OUT
x1 VDD CLK net1 VSS inverter
XM1 OUT net1 IN VDD pfet_03v3 L=0.56u W=3.36u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 OUT CLK IN VSS nfet_03v3 L=0.56u W=3.36u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  NAND.sym # of pins=5
** sym_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/NAND.sym
** sch_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/NAND.sch
.subckt NAND VDD VOUT A B VSS
*.iopin VDD
*.iopin VSS
*.ipin A
*.ipin B
*.opin VOUT
XM1 VOUT A net1 VSS nfet_03v3 L=0.56u W=2.24u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 VOUT A VDD VDD pfet_03v3 L=0.56u W=2.24u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 VOUT B VDD VDD pfet_03v3 L=0.56u W=2.24u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 net1 B VSS VSS nfet_03v3 L=0.56u W=2.24u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  3_inp_NOR.sym # of pins=6
** sym_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/3_inp_NOR.sym
** sch_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/3_inp_NOR.sch
.subckt 3_inp_NOR VDD A B C VOUT VSS
*.iopin VSS
*.iopin VDD
*.ipin A
*.ipin B
*.ipin C
*.opin VOUT
XM1 VOUT A VSS VSS nfet_03v3 L=0.56u W=1.12u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 net1 B net2 VDD pfet_03v3 L=0.56u W=6.72u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 VOUT B VSS VSS nfet_03v3 L=0.56u W=1.12u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 VOUT C VSS VSS nfet_03v3 L=0.56u W=1.12u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM5 VOUT C net1 VDD pfet_03v3 L=0.56u W=6.72u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM6 net2 A VDD VDD pfet_03v3 L=0.56u W=6.72u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  MOD_DFF_latest.sym # of pins=9
** sym_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/MOD_DFF_latest.sym
** sch_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/MOD_DFF_latest.sch
.subckt MOD_DFF_latest VDD LD DATA Q QB D1 VSS CLK G-CLK
*.iopin VDD
*.ipin LD
*.iopin VSS
*.ipin D1
*.ipin CLK
*.ipin G-CLK
*.opin Q
*.opin QB
*.ipin DATA
x1 VDD QB net1 ab net2 VSS tspc_FF
x2 VDD LD D1 net2 VSS DATA MUX
x3 VDD LD net1 Q VSS DATA MUX
x4 VDD LD CLK ab VSS G-CLK MUX
.ends


* expanding   symbol:  NOR.sym # of pins=5
** sym_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/NOR.sym
** sch_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/NOR.sch
.subckt NOR VDD A B VOUT VSS
*.iopin VSS
*.iopin VDD
*.ipin A
*.ipin B
*.opin VOUT
XM1 VOUT A VSS VSS nfet_03v3 L=0.56u W=1.12u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 VOUT B net1 VDD pfet_03v3 L=0.56u W=4.48u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 VOUT B VSS VSS nfet_03v3 L=0.56u W=1.12u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM6 net1 A VDD VDD pfet_03v3 L=0.56u W=4.48u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  tspc_FF.sym # of pins=6
** sym_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/tspc_FF.sym
** sch_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/tspc_FF.sch
.subckt tspc_FF VDD QB Q CLK D VSS
*.ipin D
*.ipin CLK
*.iopin VDD
*.iopin VSS
*.opin QB
*.opin Q
XM1 net1 D VSS VSS nfet_03v3 L=0.56u W=1.12u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 net1 CLK net2 VDD pfet_03v3 L=0.56u W=4.48u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 net2 D VDD VDD pfet_03v3 L=0.56u W=4.48u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 net3 CLK VDD VDD pfet_03v3 L=0.56u W=2.24u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM5 net3 net1 net4 VSS nfet_03v3 L=0.56u W=2.24u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM6 net4 CLK VSS VSS nfet_03v3 L=0.56u W=2.24u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM7 QB net3 VDD VDD pfet_03v3 L=0.56u W=2.24u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM8 QB CLK net5 VSS nfet_03v3 L=0.56u W=2.24u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM9 net5 net3 VSS VSS nfet_03v3 L=0.56u W=2.24u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM10 Q QB VDD VDD pfet_03v3 L=0.56u W=2.24u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM11 Q QB VSS VSS nfet_03v3 L=0.56u W=1.12u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends

.GLOBAL GND
.end
