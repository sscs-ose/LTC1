magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1112 -1856 1112 1856
<< metal1 >>
rect -112 850 112 856
rect -112 824 -106 850
rect -80 824 -44 850
rect -18 824 18 850
rect 44 824 80 850
rect 106 824 112 850
rect -112 788 112 824
rect -112 762 -106 788
rect -80 762 -44 788
rect -18 762 18 788
rect 44 762 80 788
rect 106 762 112 788
rect -112 726 112 762
rect -112 700 -106 726
rect -80 700 -44 726
rect -18 700 18 726
rect 44 700 80 726
rect 106 700 112 726
rect -112 664 112 700
rect -112 638 -106 664
rect -80 638 -44 664
rect -18 638 18 664
rect 44 638 80 664
rect 106 638 112 664
rect -112 602 112 638
rect -112 576 -106 602
rect -80 576 -44 602
rect -18 576 18 602
rect 44 576 80 602
rect 106 576 112 602
rect -112 540 112 576
rect -112 514 -106 540
rect -80 514 -44 540
rect -18 514 18 540
rect 44 514 80 540
rect 106 514 112 540
rect -112 478 112 514
rect -112 452 -106 478
rect -80 452 -44 478
rect -18 452 18 478
rect 44 452 80 478
rect 106 452 112 478
rect -112 416 112 452
rect -112 390 -106 416
rect -80 390 -44 416
rect -18 390 18 416
rect 44 390 80 416
rect 106 390 112 416
rect -112 354 112 390
rect -112 328 -106 354
rect -80 328 -44 354
rect -18 328 18 354
rect 44 328 80 354
rect 106 328 112 354
rect -112 292 112 328
rect -112 266 -106 292
rect -80 266 -44 292
rect -18 266 18 292
rect 44 266 80 292
rect 106 266 112 292
rect -112 230 112 266
rect -112 204 -106 230
rect -80 204 -44 230
rect -18 204 18 230
rect 44 204 80 230
rect 106 204 112 230
rect -112 168 112 204
rect -112 142 -106 168
rect -80 142 -44 168
rect -18 142 18 168
rect 44 142 80 168
rect 106 142 112 168
rect -112 106 112 142
rect -112 80 -106 106
rect -80 80 -44 106
rect -18 80 18 106
rect 44 80 80 106
rect 106 80 112 106
rect -112 44 112 80
rect -112 18 -106 44
rect -80 18 -44 44
rect -18 18 18 44
rect 44 18 80 44
rect 106 18 112 44
rect -112 -18 112 18
rect -112 -44 -106 -18
rect -80 -44 -44 -18
rect -18 -44 18 -18
rect 44 -44 80 -18
rect 106 -44 112 -18
rect -112 -80 112 -44
rect -112 -106 -106 -80
rect -80 -106 -44 -80
rect -18 -106 18 -80
rect 44 -106 80 -80
rect 106 -106 112 -80
rect -112 -142 112 -106
rect -112 -168 -106 -142
rect -80 -168 -44 -142
rect -18 -168 18 -142
rect 44 -168 80 -142
rect 106 -168 112 -142
rect -112 -204 112 -168
rect -112 -230 -106 -204
rect -80 -230 -44 -204
rect -18 -230 18 -204
rect 44 -230 80 -204
rect 106 -230 112 -204
rect -112 -266 112 -230
rect -112 -292 -106 -266
rect -80 -292 -44 -266
rect -18 -292 18 -266
rect 44 -292 80 -266
rect 106 -292 112 -266
rect -112 -328 112 -292
rect -112 -354 -106 -328
rect -80 -354 -44 -328
rect -18 -354 18 -328
rect 44 -354 80 -328
rect 106 -354 112 -328
rect -112 -390 112 -354
rect -112 -416 -106 -390
rect -80 -416 -44 -390
rect -18 -416 18 -390
rect 44 -416 80 -390
rect 106 -416 112 -390
rect -112 -452 112 -416
rect -112 -478 -106 -452
rect -80 -478 -44 -452
rect -18 -478 18 -452
rect 44 -478 80 -452
rect 106 -478 112 -452
rect -112 -514 112 -478
rect -112 -540 -106 -514
rect -80 -540 -44 -514
rect -18 -540 18 -514
rect 44 -540 80 -514
rect 106 -540 112 -514
rect -112 -576 112 -540
rect -112 -602 -106 -576
rect -80 -602 -44 -576
rect -18 -602 18 -576
rect 44 -602 80 -576
rect 106 -602 112 -576
rect -112 -638 112 -602
rect -112 -664 -106 -638
rect -80 -664 -44 -638
rect -18 -664 18 -638
rect 44 -664 80 -638
rect 106 -664 112 -638
rect -112 -700 112 -664
rect -112 -726 -106 -700
rect -80 -726 -44 -700
rect -18 -726 18 -700
rect 44 -726 80 -700
rect 106 -726 112 -700
rect -112 -762 112 -726
rect -112 -788 -106 -762
rect -80 -788 -44 -762
rect -18 -788 18 -762
rect 44 -788 80 -762
rect 106 -788 112 -762
rect -112 -824 112 -788
rect -112 -850 -106 -824
rect -80 -850 -44 -824
rect -18 -850 18 -824
rect 44 -850 80 -824
rect 106 -850 112 -824
rect -112 -856 112 -850
<< via1 >>
rect -106 824 -80 850
rect -44 824 -18 850
rect 18 824 44 850
rect 80 824 106 850
rect -106 762 -80 788
rect -44 762 -18 788
rect 18 762 44 788
rect 80 762 106 788
rect -106 700 -80 726
rect -44 700 -18 726
rect 18 700 44 726
rect 80 700 106 726
rect -106 638 -80 664
rect -44 638 -18 664
rect 18 638 44 664
rect 80 638 106 664
rect -106 576 -80 602
rect -44 576 -18 602
rect 18 576 44 602
rect 80 576 106 602
rect -106 514 -80 540
rect -44 514 -18 540
rect 18 514 44 540
rect 80 514 106 540
rect -106 452 -80 478
rect -44 452 -18 478
rect 18 452 44 478
rect 80 452 106 478
rect -106 390 -80 416
rect -44 390 -18 416
rect 18 390 44 416
rect 80 390 106 416
rect -106 328 -80 354
rect -44 328 -18 354
rect 18 328 44 354
rect 80 328 106 354
rect -106 266 -80 292
rect -44 266 -18 292
rect 18 266 44 292
rect 80 266 106 292
rect -106 204 -80 230
rect -44 204 -18 230
rect 18 204 44 230
rect 80 204 106 230
rect -106 142 -80 168
rect -44 142 -18 168
rect 18 142 44 168
rect 80 142 106 168
rect -106 80 -80 106
rect -44 80 -18 106
rect 18 80 44 106
rect 80 80 106 106
rect -106 18 -80 44
rect -44 18 -18 44
rect 18 18 44 44
rect 80 18 106 44
rect -106 -44 -80 -18
rect -44 -44 -18 -18
rect 18 -44 44 -18
rect 80 -44 106 -18
rect -106 -106 -80 -80
rect -44 -106 -18 -80
rect 18 -106 44 -80
rect 80 -106 106 -80
rect -106 -168 -80 -142
rect -44 -168 -18 -142
rect 18 -168 44 -142
rect 80 -168 106 -142
rect -106 -230 -80 -204
rect -44 -230 -18 -204
rect 18 -230 44 -204
rect 80 -230 106 -204
rect -106 -292 -80 -266
rect -44 -292 -18 -266
rect 18 -292 44 -266
rect 80 -292 106 -266
rect -106 -354 -80 -328
rect -44 -354 -18 -328
rect 18 -354 44 -328
rect 80 -354 106 -328
rect -106 -416 -80 -390
rect -44 -416 -18 -390
rect 18 -416 44 -390
rect 80 -416 106 -390
rect -106 -478 -80 -452
rect -44 -478 -18 -452
rect 18 -478 44 -452
rect 80 -478 106 -452
rect -106 -540 -80 -514
rect -44 -540 -18 -514
rect 18 -540 44 -514
rect 80 -540 106 -514
rect -106 -602 -80 -576
rect -44 -602 -18 -576
rect 18 -602 44 -576
rect 80 -602 106 -576
rect -106 -664 -80 -638
rect -44 -664 -18 -638
rect 18 -664 44 -638
rect 80 -664 106 -638
rect -106 -726 -80 -700
rect -44 -726 -18 -700
rect 18 -726 44 -700
rect 80 -726 106 -700
rect -106 -788 -80 -762
rect -44 -788 -18 -762
rect 18 -788 44 -762
rect 80 -788 106 -762
rect -106 -850 -80 -824
rect -44 -850 -18 -824
rect 18 -850 44 -824
rect 80 -850 106 -824
<< metal2 >>
rect -112 850 112 856
rect -112 824 -106 850
rect -80 824 -44 850
rect -18 824 18 850
rect 44 824 80 850
rect 106 824 112 850
rect -112 788 112 824
rect -112 762 -106 788
rect -80 762 -44 788
rect -18 762 18 788
rect 44 762 80 788
rect 106 762 112 788
rect -112 726 112 762
rect -112 700 -106 726
rect -80 700 -44 726
rect -18 700 18 726
rect 44 700 80 726
rect 106 700 112 726
rect -112 664 112 700
rect -112 638 -106 664
rect -80 638 -44 664
rect -18 638 18 664
rect 44 638 80 664
rect 106 638 112 664
rect -112 602 112 638
rect -112 576 -106 602
rect -80 576 -44 602
rect -18 576 18 602
rect 44 576 80 602
rect 106 576 112 602
rect -112 540 112 576
rect -112 514 -106 540
rect -80 514 -44 540
rect -18 514 18 540
rect 44 514 80 540
rect 106 514 112 540
rect -112 478 112 514
rect -112 452 -106 478
rect -80 452 -44 478
rect -18 452 18 478
rect 44 452 80 478
rect 106 452 112 478
rect -112 416 112 452
rect -112 390 -106 416
rect -80 390 -44 416
rect -18 390 18 416
rect 44 390 80 416
rect 106 390 112 416
rect -112 354 112 390
rect -112 328 -106 354
rect -80 328 -44 354
rect -18 328 18 354
rect 44 328 80 354
rect 106 328 112 354
rect -112 292 112 328
rect -112 266 -106 292
rect -80 266 -44 292
rect -18 266 18 292
rect 44 266 80 292
rect 106 266 112 292
rect -112 230 112 266
rect -112 204 -106 230
rect -80 204 -44 230
rect -18 204 18 230
rect 44 204 80 230
rect 106 204 112 230
rect -112 168 112 204
rect -112 142 -106 168
rect -80 142 -44 168
rect -18 142 18 168
rect 44 142 80 168
rect 106 142 112 168
rect -112 106 112 142
rect -112 80 -106 106
rect -80 80 -44 106
rect -18 80 18 106
rect 44 80 80 106
rect 106 80 112 106
rect -112 44 112 80
rect -112 18 -106 44
rect -80 18 -44 44
rect -18 18 18 44
rect 44 18 80 44
rect 106 18 112 44
rect -112 -18 112 18
rect -112 -44 -106 -18
rect -80 -44 -44 -18
rect -18 -44 18 -18
rect 44 -44 80 -18
rect 106 -44 112 -18
rect -112 -80 112 -44
rect -112 -106 -106 -80
rect -80 -106 -44 -80
rect -18 -106 18 -80
rect 44 -106 80 -80
rect 106 -106 112 -80
rect -112 -142 112 -106
rect -112 -168 -106 -142
rect -80 -168 -44 -142
rect -18 -168 18 -142
rect 44 -168 80 -142
rect 106 -168 112 -142
rect -112 -204 112 -168
rect -112 -230 -106 -204
rect -80 -230 -44 -204
rect -18 -230 18 -204
rect 44 -230 80 -204
rect 106 -230 112 -204
rect -112 -266 112 -230
rect -112 -292 -106 -266
rect -80 -292 -44 -266
rect -18 -292 18 -266
rect 44 -292 80 -266
rect 106 -292 112 -266
rect -112 -328 112 -292
rect -112 -354 -106 -328
rect -80 -354 -44 -328
rect -18 -354 18 -328
rect 44 -354 80 -328
rect 106 -354 112 -328
rect -112 -390 112 -354
rect -112 -416 -106 -390
rect -80 -416 -44 -390
rect -18 -416 18 -390
rect 44 -416 80 -390
rect 106 -416 112 -390
rect -112 -452 112 -416
rect -112 -478 -106 -452
rect -80 -478 -44 -452
rect -18 -478 18 -452
rect 44 -478 80 -452
rect 106 -478 112 -452
rect -112 -514 112 -478
rect -112 -540 -106 -514
rect -80 -540 -44 -514
rect -18 -540 18 -514
rect 44 -540 80 -514
rect 106 -540 112 -514
rect -112 -576 112 -540
rect -112 -602 -106 -576
rect -80 -602 -44 -576
rect -18 -602 18 -576
rect 44 -602 80 -576
rect 106 -602 112 -576
rect -112 -638 112 -602
rect -112 -664 -106 -638
rect -80 -664 -44 -638
rect -18 -664 18 -638
rect 44 -664 80 -638
rect 106 -664 112 -638
rect -112 -700 112 -664
rect -112 -726 -106 -700
rect -80 -726 -44 -700
rect -18 -726 18 -700
rect 44 -726 80 -700
rect 106 -726 112 -700
rect -112 -762 112 -726
rect -112 -788 -106 -762
rect -80 -788 -44 -762
rect -18 -788 18 -762
rect 44 -788 80 -762
rect 106 -788 112 -762
rect -112 -824 112 -788
rect -112 -850 -106 -824
rect -80 -850 -44 -824
rect -18 -850 18 -824
rect 44 -850 80 -824
rect 106 -850 112 -824
rect -112 -856 112 -850
<< end >>
