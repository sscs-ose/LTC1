magic
tech gf180mcuC
magscale 1 10
timestamp 1691568605
<< nwell >>
rect -209 -330 209 330
<< pmos >>
rect -35 -200 35 200
<< pdiff >>
rect -123 187 -35 200
rect -123 -187 -110 187
rect -64 -187 -35 187
rect -123 -200 -35 -187
rect 35 187 123 200
rect 35 -187 64 187
rect 110 -187 123 187
rect 35 -200 123 -187
<< pdiffc >>
rect -110 -187 -64 187
rect 64 -187 110 187
<< polysilicon >>
rect -35 200 35 244
rect -35 -244 35 -200
<< metal1 >>
rect -110 187 -64 198
rect -110 -198 -64 -187
rect 64 187 110 198
rect 64 -198 110 -187
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 2 l 0.35 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
