* NGSPICE file created from Local_Enc_v2.ext - technology: gf180mcuC

.subckt pmos_3p3_M8RWPS a_n28_n94# w_n202_n180# a_n116_n50# a_28_n50#
X0 a_28_n50# a_n28_n94# a_n116_n50# w_n202_n180# pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
.ends

.subckt nmos_3p3_HZS5UA a_n28_n94# a_n116_n50# a_28_n50# VSUBS
X0 a_28_n50# a_n28_n94# a_n116_n50# VSUBS nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
.ends

.subckt NAND VDD VSS B A OUT
Xpmos_3p3_M8RWPS_0 A VDD VDD OUT pmos_3p3_M8RWPS
Xpmos_3p3_M8RWPS_1 B VDD VDD OUT pmos_3p3_M8RWPS
Xnmos_3p3_HZS5UA_0 A m1_184_67# OUT VSS nmos_3p3_HZS5UA
Xnmos_3p3_HZS5UA_1 B VSS m1_184_67# VSS nmos_3p3_HZS5UA
.ends

.subckt Local_Enc_v2 QB Q Ri-1 Ri Ci
XNAND_0 NAND_9/VDD VSUBS Ci Ci NAND_12/B NAND
XNAND_1 NAND_9/VDD VSUBS NAND_1/B NAND_1/B NAND_13/B NAND
XNAND_2 NAND_9/VDD VSUBS NAND_9/B NAND_9/B NAND_3/B NAND
XNAND_3 NAND_9/VDD VSUBS NAND_3/B Q QB NAND
XNAND_9 NAND_9/VDD VSUBS NAND_9/B QB Q NAND
XNAND_11 NAND_9/VDD VSUBS Ri Ri NAND_12/A NAND
XNAND_12 NAND_9/VDD VSUBS NAND_12/B NAND_12/A NAND_13/A NAND
XNAND_13 NAND_9/VDD VSUBS NAND_13/B NAND_13/A NAND_9/B NAND
XNAND_14 NAND_9/VDD VSUBS Ri-1 Ri-1 NAND_1/B NAND
.ends

