magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1247 -1551 1247 1551
<< metal2 >>
rect -247 546 247 551
rect -247 518 -242 546
rect -214 518 -166 546
rect -138 518 -90 546
rect -62 518 -14 546
rect 14 518 62 546
rect 90 518 138 546
rect 166 518 214 546
rect 242 518 247 546
rect -247 470 247 518
rect -247 442 -242 470
rect -214 442 -166 470
rect -138 442 -90 470
rect -62 442 -14 470
rect 14 442 62 470
rect 90 442 138 470
rect 166 442 214 470
rect 242 442 247 470
rect -247 394 247 442
rect -247 366 -242 394
rect -214 366 -166 394
rect -138 366 -90 394
rect -62 366 -14 394
rect 14 366 62 394
rect 90 366 138 394
rect 166 366 214 394
rect 242 366 247 394
rect -247 318 247 366
rect -247 290 -242 318
rect -214 290 -166 318
rect -138 290 -90 318
rect -62 290 -14 318
rect 14 290 62 318
rect 90 290 138 318
rect 166 290 214 318
rect 242 290 247 318
rect -247 242 247 290
rect -247 214 -242 242
rect -214 214 -166 242
rect -138 214 -90 242
rect -62 214 -14 242
rect 14 214 62 242
rect 90 214 138 242
rect 166 214 214 242
rect 242 214 247 242
rect -247 166 247 214
rect -247 138 -242 166
rect -214 138 -166 166
rect -138 138 -90 166
rect -62 138 -14 166
rect 14 138 62 166
rect 90 138 138 166
rect 166 138 214 166
rect 242 138 247 166
rect -247 90 247 138
rect -247 62 -242 90
rect -214 62 -166 90
rect -138 62 -90 90
rect -62 62 -14 90
rect 14 62 62 90
rect 90 62 138 90
rect 166 62 214 90
rect 242 62 247 90
rect -247 14 247 62
rect -247 -14 -242 14
rect -214 -14 -166 14
rect -138 -14 -90 14
rect -62 -14 -14 14
rect 14 -14 62 14
rect 90 -14 138 14
rect 166 -14 214 14
rect 242 -14 247 14
rect -247 -62 247 -14
rect -247 -90 -242 -62
rect -214 -90 -166 -62
rect -138 -90 -90 -62
rect -62 -90 -14 -62
rect 14 -90 62 -62
rect 90 -90 138 -62
rect 166 -90 214 -62
rect 242 -90 247 -62
rect -247 -138 247 -90
rect -247 -166 -242 -138
rect -214 -166 -166 -138
rect -138 -166 -90 -138
rect -62 -166 -14 -138
rect 14 -166 62 -138
rect 90 -166 138 -138
rect 166 -166 214 -138
rect 242 -166 247 -138
rect -247 -214 247 -166
rect -247 -242 -242 -214
rect -214 -242 -166 -214
rect -138 -242 -90 -214
rect -62 -242 -14 -214
rect 14 -242 62 -214
rect 90 -242 138 -214
rect 166 -242 214 -214
rect 242 -242 247 -214
rect -247 -290 247 -242
rect -247 -318 -242 -290
rect -214 -318 -166 -290
rect -138 -318 -90 -290
rect -62 -318 -14 -290
rect 14 -318 62 -290
rect 90 -318 138 -290
rect 166 -318 214 -290
rect 242 -318 247 -290
rect -247 -366 247 -318
rect -247 -394 -242 -366
rect -214 -394 -166 -366
rect -138 -394 -90 -366
rect -62 -394 -14 -366
rect 14 -394 62 -366
rect 90 -394 138 -366
rect 166 -394 214 -366
rect 242 -394 247 -366
rect -247 -442 247 -394
rect -247 -470 -242 -442
rect -214 -470 -166 -442
rect -138 -470 -90 -442
rect -62 -470 -14 -442
rect 14 -470 62 -442
rect 90 -470 138 -442
rect 166 -470 214 -442
rect 242 -470 247 -442
rect -247 -518 247 -470
rect -247 -546 -242 -518
rect -214 -546 -166 -518
rect -138 -546 -90 -518
rect -62 -546 -14 -518
rect 14 -546 62 -518
rect 90 -546 138 -518
rect 166 -546 214 -518
rect 242 -546 247 -518
rect -247 -551 247 -546
<< via2 >>
rect -242 518 -214 546
rect -166 518 -138 546
rect -90 518 -62 546
rect -14 518 14 546
rect 62 518 90 546
rect 138 518 166 546
rect 214 518 242 546
rect -242 442 -214 470
rect -166 442 -138 470
rect -90 442 -62 470
rect -14 442 14 470
rect 62 442 90 470
rect 138 442 166 470
rect 214 442 242 470
rect -242 366 -214 394
rect -166 366 -138 394
rect -90 366 -62 394
rect -14 366 14 394
rect 62 366 90 394
rect 138 366 166 394
rect 214 366 242 394
rect -242 290 -214 318
rect -166 290 -138 318
rect -90 290 -62 318
rect -14 290 14 318
rect 62 290 90 318
rect 138 290 166 318
rect 214 290 242 318
rect -242 214 -214 242
rect -166 214 -138 242
rect -90 214 -62 242
rect -14 214 14 242
rect 62 214 90 242
rect 138 214 166 242
rect 214 214 242 242
rect -242 138 -214 166
rect -166 138 -138 166
rect -90 138 -62 166
rect -14 138 14 166
rect 62 138 90 166
rect 138 138 166 166
rect 214 138 242 166
rect -242 62 -214 90
rect -166 62 -138 90
rect -90 62 -62 90
rect -14 62 14 90
rect 62 62 90 90
rect 138 62 166 90
rect 214 62 242 90
rect -242 -14 -214 14
rect -166 -14 -138 14
rect -90 -14 -62 14
rect -14 -14 14 14
rect 62 -14 90 14
rect 138 -14 166 14
rect 214 -14 242 14
rect -242 -90 -214 -62
rect -166 -90 -138 -62
rect -90 -90 -62 -62
rect -14 -90 14 -62
rect 62 -90 90 -62
rect 138 -90 166 -62
rect 214 -90 242 -62
rect -242 -166 -214 -138
rect -166 -166 -138 -138
rect -90 -166 -62 -138
rect -14 -166 14 -138
rect 62 -166 90 -138
rect 138 -166 166 -138
rect 214 -166 242 -138
rect -242 -242 -214 -214
rect -166 -242 -138 -214
rect -90 -242 -62 -214
rect -14 -242 14 -214
rect 62 -242 90 -214
rect 138 -242 166 -214
rect 214 -242 242 -214
rect -242 -318 -214 -290
rect -166 -318 -138 -290
rect -90 -318 -62 -290
rect -14 -318 14 -290
rect 62 -318 90 -290
rect 138 -318 166 -290
rect 214 -318 242 -290
rect -242 -394 -214 -366
rect -166 -394 -138 -366
rect -90 -394 -62 -366
rect -14 -394 14 -366
rect 62 -394 90 -366
rect 138 -394 166 -366
rect 214 -394 242 -366
rect -242 -470 -214 -442
rect -166 -470 -138 -442
rect -90 -470 -62 -442
rect -14 -470 14 -442
rect 62 -470 90 -442
rect 138 -470 166 -442
rect 214 -470 242 -442
rect -242 -546 -214 -518
rect -166 -546 -138 -518
rect -90 -546 -62 -518
rect -14 -546 14 -518
rect 62 -546 90 -518
rect 138 -546 166 -518
rect 214 -546 242 -518
<< metal3 >>
rect -247 546 247 551
rect -247 518 -242 546
rect -214 518 -166 546
rect -138 518 -90 546
rect -62 518 -14 546
rect 14 518 62 546
rect 90 518 138 546
rect 166 518 214 546
rect 242 518 247 546
rect -247 470 247 518
rect -247 442 -242 470
rect -214 442 -166 470
rect -138 442 -90 470
rect -62 442 -14 470
rect 14 442 62 470
rect 90 442 138 470
rect 166 442 214 470
rect 242 442 247 470
rect -247 394 247 442
rect -247 366 -242 394
rect -214 366 -166 394
rect -138 366 -90 394
rect -62 366 -14 394
rect 14 366 62 394
rect 90 366 138 394
rect 166 366 214 394
rect 242 366 247 394
rect -247 318 247 366
rect -247 290 -242 318
rect -214 290 -166 318
rect -138 290 -90 318
rect -62 290 -14 318
rect 14 290 62 318
rect 90 290 138 318
rect 166 290 214 318
rect 242 290 247 318
rect -247 242 247 290
rect -247 214 -242 242
rect -214 214 -166 242
rect -138 214 -90 242
rect -62 214 -14 242
rect 14 214 62 242
rect 90 214 138 242
rect 166 214 214 242
rect 242 214 247 242
rect -247 166 247 214
rect -247 138 -242 166
rect -214 138 -166 166
rect -138 138 -90 166
rect -62 138 -14 166
rect 14 138 62 166
rect 90 138 138 166
rect 166 138 214 166
rect 242 138 247 166
rect -247 90 247 138
rect -247 62 -242 90
rect -214 62 -166 90
rect -138 62 -90 90
rect -62 62 -14 90
rect 14 62 62 90
rect 90 62 138 90
rect 166 62 214 90
rect 242 62 247 90
rect -247 14 247 62
rect -247 -14 -242 14
rect -214 -14 -166 14
rect -138 -14 -90 14
rect -62 -14 -14 14
rect 14 -14 62 14
rect 90 -14 138 14
rect 166 -14 214 14
rect 242 -14 247 14
rect -247 -62 247 -14
rect -247 -90 -242 -62
rect -214 -90 -166 -62
rect -138 -90 -90 -62
rect -62 -90 -14 -62
rect 14 -90 62 -62
rect 90 -90 138 -62
rect 166 -90 214 -62
rect 242 -90 247 -62
rect -247 -138 247 -90
rect -247 -166 -242 -138
rect -214 -166 -166 -138
rect -138 -166 -90 -138
rect -62 -166 -14 -138
rect 14 -166 62 -138
rect 90 -166 138 -138
rect 166 -166 214 -138
rect 242 -166 247 -138
rect -247 -214 247 -166
rect -247 -242 -242 -214
rect -214 -242 -166 -214
rect -138 -242 -90 -214
rect -62 -242 -14 -214
rect 14 -242 62 -214
rect 90 -242 138 -214
rect 166 -242 214 -214
rect 242 -242 247 -214
rect -247 -290 247 -242
rect -247 -318 -242 -290
rect -214 -318 -166 -290
rect -138 -318 -90 -290
rect -62 -318 -14 -290
rect 14 -318 62 -290
rect 90 -318 138 -290
rect 166 -318 214 -290
rect 242 -318 247 -290
rect -247 -366 247 -318
rect -247 -394 -242 -366
rect -214 -394 -166 -366
rect -138 -394 -90 -366
rect -62 -394 -14 -366
rect 14 -394 62 -366
rect 90 -394 138 -366
rect 166 -394 214 -366
rect 242 -394 247 -366
rect -247 -442 247 -394
rect -247 -470 -242 -442
rect -214 -470 -166 -442
rect -138 -470 -90 -442
rect -62 -470 -14 -442
rect 14 -470 62 -442
rect 90 -470 138 -442
rect 166 -470 214 -442
rect 242 -470 247 -442
rect -247 -518 247 -470
rect -247 -546 -242 -518
rect -214 -546 -166 -518
rect -138 -546 -90 -518
rect -62 -546 -14 -518
rect 14 -546 62 -518
rect 90 -546 138 -518
rect 166 -546 214 -518
rect 242 -546 247 -518
rect -247 -551 247 -546
<< end >>
