magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1931 -1019 1931 1019
<< metal1 >>
rect -931 13 931 19
rect -931 -13 -925 13
rect -899 -13 -849 13
rect -823 -13 -773 13
rect -747 -13 -697 13
rect -671 -13 -621 13
rect -595 -13 -545 13
rect -519 -13 -469 13
rect -443 -13 -393 13
rect -367 -13 -317 13
rect -291 -13 -241 13
rect -215 -13 -165 13
rect -139 -13 -89 13
rect -63 -13 -13 13
rect 13 -13 63 13
rect 89 -13 139 13
rect 165 -13 215 13
rect 241 -13 291 13
rect 317 -13 367 13
rect 393 -13 443 13
rect 469 -13 519 13
rect 545 -13 595 13
rect 621 -13 671 13
rect 697 -13 747 13
rect 773 -13 823 13
rect 849 -13 899 13
rect 925 -13 931 13
rect -931 -19 931 -13
<< via1 >>
rect -925 -13 -899 13
rect -849 -13 -823 13
rect -773 -13 -747 13
rect -697 -13 -671 13
rect -621 -13 -595 13
rect -545 -13 -519 13
rect -469 -13 -443 13
rect -393 -13 -367 13
rect -317 -13 -291 13
rect -241 -13 -215 13
rect -165 -13 -139 13
rect -89 -13 -63 13
rect -13 -13 13 13
rect 63 -13 89 13
rect 139 -13 165 13
rect 215 -13 241 13
rect 291 -13 317 13
rect 367 -13 393 13
rect 443 -13 469 13
rect 519 -13 545 13
rect 595 -13 621 13
rect 671 -13 697 13
rect 747 -13 773 13
rect 823 -13 849 13
rect 899 -13 925 13
<< metal2 >>
rect -931 13 931 19
rect -931 -13 -925 13
rect -899 -13 -849 13
rect -823 -13 -773 13
rect -747 -13 -697 13
rect -671 -13 -621 13
rect -595 -13 -545 13
rect -519 -13 -469 13
rect -443 -13 -393 13
rect -367 -13 -317 13
rect -291 -13 -241 13
rect -215 -13 -165 13
rect -139 -13 -89 13
rect -63 -13 -13 13
rect 13 -13 63 13
rect 89 -13 139 13
rect 165 -13 215 13
rect 241 -13 291 13
rect 317 -13 367 13
rect 393 -13 443 13
rect 469 -13 519 13
rect 545 -13 595 13
rect 621 -13 671 13
rect 697 -13 747 13
rect 773 -13 823 13
rect 849 -13 899 13
rect 925 -13 931 13
rect -931 -19 931 -13
<< end >>
