magic
tech gf180mcuC
magscale 1 10
timestamp 1695121232
<< nwell >>
rect -40 -1170 3230 490
<< psubdiff >>
rect -231 642 3409 681
rect -231 628 41 642
rect -231 571 -187 628
rect -130 585 41 628
rect 98 585 246 642
rect 303 585 451 642
rect 508 585 656 642
rect 713 585 861 642
rect 918 585 1066 642
rect 1123 585 1271 642
rect 1328 585 1476 642
rect 1533 585 1681 642
rect 1738 585 1886 642
rect 1943 585 2091 642
rect 2148 585 2296 642
rect 2353 585 2501 642
rect 2558 585 2706 642
rect 2763 585 2911 642
rect 2968 585 3116 642
rect 3173 585 3321 642
rect 3378 585 3409 642
rect -130 571 3409 585
rect -231 541 3409 571
rect -231 423 -91 541
rect -231 366 -187 423
rect -130 366 -91 423
rect -231 218 -91 366
rect -231 161 -187 218
rect -130 161 -91 218
rect -231 13 -91 161
rect -231 -44 -187 13
rect -130 -44 -91 13
rect -231 -192 -91 -44
rect -231 -249 -187 -192
rect -130 -249 -91 -192
rect -231 -397 -91 -249
rect -231 -454 -187 -397
rect -130 -454 -91 -397
rect -231 -602 -91 -454
rect -231 -659 -187 -602
rect -130 -659 -91 -602
rect -231 -807 -91 -659
rect -231 -864 -187 -807
rect -130 -864 -91 -807
rect -231 -1012 -91 -864
rect -231 -1069 -187 -1012
rect -130 -1069 -91 -1012
rect -231 -1199 -91 -1069
rect 3269 423 3409 541
rect 3269 366 3313 423
rect 3370 366 3409 423
rect 3269 218 3409 366
rect 3269 161 3313 218
rect 3370 161 3409 218
rect 3269 13 3409 161
rect 3269 -44 3313 13
rect 3370 -44 3409 13
rect 3269 -192 3409 -44
rect 3269 -249 3313 -192
rect 3370 -249 3409 -192
rect 3269 -397 3409 -249
rect 3269 -454 3313 -397
rect 3370 -454 3409 -397
rect 3269 -602 3409 -454
rect 3269 -659 3313 -602
rect 3370 -659 3409 -602
rect 3269 -807 3409 -659
rect 3269 -864 3313 -807
rect 3370 -864 3409 -807
rect 3269 -1012 3409 -864
rect 3269 -1069 3313 -1012
rect 3370 -1069 3409 -1012
rect 3269 -1199 3409 -1069
rect -231 -1217 3409 -1199
rect -231 -1274 -187 -1217
rect -130 -1243 3313 -1217
rect -130 -1274 4 -1243
rect -231 -1300 4 -1274
rect 61 -1300 209 -1243
rect 266 -1300 414 -1243
rect 471 -1300 619 -1243
rect 676 -1300 824 -1243
rect 881 -1300 1029 -1243
rect 1086 -1300 1234 -1243
rect 1291 -1300 1439 -1243
rect 1496 -1300 1644 -1243
rect 1701 -1300 1849 -1243
rect 1906 -1300 2054 -1243
rect 2111 -1300 2259 -1243
rect 2316 -1300 2464 -1243
rect 2521 -1300 2669 -1243
rect 2726 -1300 2874 -1243
rect 2931 -1300 3079 -1243
rect 3136 -1274 3313 -1243
rect 3370 -1274 3409 -1217
rect 3136 -1300 3409 -1274
rect -231 -1339 3409 -1300
rect -231 -1422 -91 -1339
rect -231 -1479 -187 -1422
rect -130 -1479 -91 -1422
rect 3269 -1422 3409 -1339
rect -231 -1627 -91 -1479
rect 3269 -1479 3313 -1422
rect 3370 -1479 3409 -1422
rect -231 -1684 -187 -1627
rect -130 -1684 -91 -1627
rect -231 -1832 -91 -1684
rect -231 -1889 -187 -1832
rect -130 -1889 -91 -1832
rect -231 -2037 -91 -1889
rect 3269 -1627 3409 -1479
rect 3269 -1684 3313 -1627
rect 3370 -1684 3409 -1627
rect 3269 -1832 3409 -1684
rect 3269 -1889 3313 -1832
rect 3370 -1889 3409 -1832
rect -231 -2094 -187 -2037
rect -130 -2094 -91 -2037
rect 3269 -2037 3409 -1889
rect -231 -2242 -91 -2094
rect -231 -2299 -187 -2242
rect -130 -2299 -91 -2242
rect -231 -2447 -91 -2299
rect 3269 -2094 3313 -2037
rect 3370 -2094 3409 -2037
rect 3269 -2242 3409 -2094
rect 3269 -2299 3313 -2242
rect 3370 -2299 3409 -2242
rect -231 -2504 -187 -2447
rect -130 -2504 -91 -2447
rect 3269 -2447 3409 -2299
rect -231 -2599 -91 -2504
rect 3269 -2504 3313 -2447
rect 3370 -2504 3409 -2447
rect 3269 -2599 3409 -2504
rect -231 -2643 3409 -2599
rect -231 -2700 -185 -2643
rect -128 -2700 4 -2643
rect 61 -2700 209 -2643
rect 266 -2700 414 -2643
rect 471 -2700 619 -2643
rect 676 -2700 824 -2643
rect 881 -2700 1029 -2643
rect 1086 -2700 1234 -2643
rect 1291 -2700 1439 -2643
rect 1496 -2700 1644 -2643
rect 1701 -2700 1849 -2643
rect 1906 -2700 2054 -2643
rect 2111 -2700 2259 -2643
rect 2316 -2700 2464 -2643
rect 2521 -2700 2669 -2643
rect 2726 -2700 2874 -2643
rect 2931 -2700 3079 -2643
rect 3136 -2700 3316 -2643
rect 3373 -2700 3409 -2643
rect -231 -2739 3409 -2700
<< nsubdiff >>
rect 10 413 3170 440
rect 10 368 245 413
rect 10 320 40 368
rect 88 365 245 368
rect 293 365 450 413
rect 498 365 655 413
rect 703 365 860 413
rect 908 365 1065 413
rect 1113 365 1270 413
rect 1318 365 1475 413
rect 1523 365 1680 413
rect 1728 365 1885 413
rect 1933 365 2090 413
rect 2138 365 2295 413
rect 2343 365 2500 413
rect 2548 365 2705 413
rect 2753 365 2910 413
rect 2958 368 3170 413
rect 2958 365 3090 368
rect 88 340 3090 365
rect 88 320 120 340
rect 10 168 120 320
rect 10 120 40 168
rect 88 120 120 168
rect 10 -32 120 120
rect 10 -80 40 -32
rect 88 -80 120 -32
rect 10 -232 120 -80
rect 3060 320 3090 340
rect 3138 320 3170 368
rect 3060 168 3170 320
rect 3060 120 3090 168
rect 3138 120 3170 168
rect 3060 -32 3170 120
rect 3060 -80 3090 -32
rect 3138 -80 3170 -32
rect 10 -280 40 -232
rect 88 -280 120 -232
rect 10 -432 120 -280
rect 3060 -232 3170 -80
rect 3060 -280 3090 -232
rect 3138 -280 3170 -232
rect 10 -480 40 -432
rect 88 -480 120 -432
rect 10 -632 120 -480
rect 10 -680 40 -632
rect 88 -680 120 -632
rect 10 -832 120 -680
rect 3060 -432 3170 -280
rect 3060 -480 3090 -432
rect 3138 -480 3170 -432
rect 3060 -632 3170 -480
rect 3060 -680 3090 -632
rect 3138 -680 3170 -632
rect 10 -880 40 -832
rect 88 -880 120 -832
rect 3060 -832 3170 -680
rect 10 -1010 120 -880
rect 3060 -880 3090 -832
rect 3138 -880 3170 -832
rect 3060 -1010 3170 -880
rect 10 -1032 3170 -1010
rect 10 -1080 40 -1032
rect 88 -1080 245 -1032
rect 293 -1080 450 -1032
rect 498 -1080 655 -1032
rect 703 -1080 860 -1032
rect 908 -1080 1065 -1032
rect 1113 -1080 1270 -1032
rect 1318 -1080 1475 -1032
rect 1523 -1080 1680 -1032
rect 1728 -1080 1885 -1032
rect 1933 -1080 2090 -1032
rect 2138 -1080 2295 -1032
rect 2343 -1080 2500 -1032
rect 2548 -1080 2705 -1032
rect 2753 -1080 2910 -1032
rect 2958 -1080 3090 -1032
rect 3138 -1080 3170 -1032
rect 10 -1110 3170 -1080
<< psubdiffcont >>
rect -187 571 -130 628
rect 41 585 98 642
rect 246 585 303 642
rect 451 585 508 642
rect 656 585 713 642
rect 861 585 918 642
rect 1066 585 1123 642
rect 1271 585 1328 642
rect 1476 585 1533 642
rect 1681 585 1738 642
rect 1886 585 1943 642
rect 2091 585 2148 642
rect 2296 585 2353 642
rect 2501 585 2558 642
rect 2706 585 2763 642
rect 2911 585 2968 642
rect 3116 585 3173 642
rect 3321 585 3378 642
rect -187 366 -130 423
rect -187 161 -130 218
rect -187 -44 -130 13
rect -187 -249 -130 -192
rect -187 -454 -130 -397
rect -187 -659 -130 -602
rect -187 -864 -130 -807
rect -187 -1069 -130 -1012
rect 3313 366 3370 423
rect 3313 161 3370 218
rect 3313 -44 3370 13
rect 3313 -249 3370 -192
rect 3313 -454 3370 -397
rect 3313 -659 3370 -602
rect 3313 -864 3370 -807
rect 3313 -1069 3370 -1012
rect -187 -1274 -130 -1217
rect 4 -1300 61 -1243
rect 209 -1300 266 -1243
rect 414 -1300 471 -1243
rect 619 -1300 676 -1243
rect 824 -1300 881 -1243
rect 1029 -1300 1086 -1243
rect 1234 -1300 1291 -1243
rect 1439 -1300 1496 -1243
rect 1644 -1300 1701 -1243
rect 1849 -1300 1906 -1243
rect 2054 -1300 2111 -1243
rect 2259 -1300 2316 -1243
rect 2464 -1300 2521 -1243
rect 2669 -1300 2726 -1243
rect 2874 -1300 2931 -1243
rect 3079 -1300 3136 -1243
rect 3313 -1274 3370 -1217
rect -187 -1479 -130 -1422
rect 3313 -1479 3370 -1422
rect -187 -1684 -130 -1627
rect -187 -1889 -130 -1832
rect 3313 -1684 3370 -1627
rect 3313 -1889 3370 -1832
rect -187 -2094 -130 -2037
rect -187 -2299 -130 -2242
rect 3313 -2094 3370 -2037
rect 3313 -2299 3370 -2242
rect -187 -2504 -130 -2447
rect 3313 -2504 3370 -2447
rect -185 -2700 -128 -2643
rect 4 -2700 61 -2643
rect 209 -2700 266 -2643
rect 414 -2700 471 -2643
rect 619 -2700 676 -2643
rect 824 -2700 881 -2643
rect 1029 -2700 1086 -2643
rect 1234 -2700 1291 -2643
rect 1439 -2700 1496 -2643
rect 1644 -2700 1701 -2643
rect 1849 -2700 1906 -2643
rect 2054 -2700 2111 -2643
rect 2259 -2700 2316 -2643
rect 2464 -2700 2521 -2643
rect 2669 -2700 2726 -2643
rect 2874 -2700 2931 -2643
rect 3079 -2700 3136 -2643
rect 3316 -2700 3373 -2643
<< nsubdiffcont >>
rect 40 320 88 368
rect 245 365 293 413
rect 450 365 498 413
rect 655 365 703 413
rect 860 365 908 413
rect 1065 365 1113 413
rect 1270 365 1318 413
rect 1475 365 1523 413
rect 1680 365 1728 413
rect 1885 365 1933 413
rect 2090 365 2138 413
rect 2295 365 2343 413
rect 2500 365 2548 413
rect 2705 365 2753 413
rect 2910 365 2958 413
rect 40 120 88 168
rect 40 -80 88 -32
rect 3090 320 3138 368
rect 3090 120 3138 168
rect 3090 -80 3138 -32
rect 40 -280 88 -232
rect 3090 -280 3138 -232
rect 40 -480 88 -432
rect 40 -680 88 -632
rect 3090 -480 3138 -432
rect 3090 -680 3138 -632
rect 40 -880 88 -832
rect 3090 -880 3138 -832
rect 40 -1080 88 -1032
rect 245 -1080 293 -1032
rect 450 -1080 498 -1032
rect 655 -1080 703 -1032
rect 860 -1080 908 -1032
rect 1065 -1080 1113 -1032
rect 1270 -1080 1318 -1032
rect 1475 -1080 1523 -1032
rect 1680 -1080 1728 -1032
rect 1885 -1080 1933 -1032
rect 2090 -1080 2138 -1032
rect 2295 -1080 2343 -1032
rect 2500 -1080 2548 -1032
rect 2705 -1080 2753 -1032
rect 2910 -1080 2958 -1032
rect 3090 -1080 3138 -1032
<< polysilicon >>
rect 367 -194 1127 -102
rect 367 -244 394 -194
rect 444 -214 1127 -194
rect 1231 -144 1991 -103
rect 1231 -194 1802 -144
rect 1852 -194 1991 -144
rect 444 -244 464 -214
rect 1231 -215 1991 -194
rect 2095 -217 2855 -105
rect 367 -259 464 -244
rect 1015 -348 1127 -330
rect 1015 -398 1047 -348
rect 1097 -398 1127 -348
rect 1015 -424 1127 -398
rect 2743 -428 2855 -217
rect 367 -793 1127 -694
rect 366 -806 1127 -793
rect 1231 -731 1991 -695
rect 1231 -781 1434 -731
rect 1484 -781 1545 -731
rect 1595 -781 1991 -731
rect 366 -856 387 -806
rect 437 -856 463 -806
rect 1231 -807 1991 -781
rect 2095 -734 2855 -696
rect 2095 -784 2173 -734
rect 2223 -735 2855 -734
rect 2223 -784 2278 -735
rect 2095 -785 2278 -784
rect 2328 -785 2855 -735
rect 2095 -808 2855 -785
rect 366 -870 463 -856
rect 562 -1461 1754 -1437
rect 562 -1511 586 -1461
rect 636 -1511 1754 -1461
rect 562 -1549 1754 -1511
rect 1858 -1461 2618 -1438
rect 1858 -1511 2538 -1461
rect 2588 -1511 2618 -1461
rect 1858 -1549 2618 -1511
rect 562 -2001 674 -1978
rect 562 -2051 593 -2001
rect 643 -2051 674 -2001
rect 562 -2079 674 -2051
rect 2506 -2007 2618 -1983
rect 2506 -2057 2537 -2007
rect 2587 -2057 2618 -2007
rect 2506 -2079 2618 -2057
rect 778 -2386 1538 -2349
rect 778 -2436 1456 -2386
rect 1505 -2436 1538 -2386
rect 778 -2460 1538 -2436
rect 1642 -2387 2402 -2350
rect 1642 -2437 2319 -2387
rect 2369 -2437 2402 -2387
rect 1642 -2461 2402 -2437
<< polycontact >>
rect 394 -244 444 -194
rect 1802 -194 1852 -144
rect 1047 -398 1097 -348
rect 1434 -781 1484 -731
rect 1545 -781 1595 -731
rect 387 -856 437 -806
rect 2173 -784 2223 -734
rect 2278 -785 2328 -735
rect 586 -1511 636 -1461
rect 2538 -1511 2588 -1461
rect 593 -2051 643 -2001
rect 2537 -2057 2587 -2007
rect 1456 -2436 1505 -2386
rect 2319 -2437 2369 -2387
<< metal1 >>
rect -231 642 3409 681
rect -231 628 41 642
rect -231 571 -187 628
rect -130 585 41 628
rect 98 585 246 642
rect 303 585 451 642
rect 508 585 656 642
rect 713 585 861 642
rect 918 585 1066 642
rect 1123 585 1271 642
rect 1328 585 1476 642
rect 1533 585 1681 642
rect 1738 585 1886 642
rect 1943 585 2091 642
rect 2148 585 2296 642
rect 2353 585 2501 642
rect 2558 585 2706 642
rect 2763 585 2911 642
rect 2968 585 3116 642
rect 3173 585 3321 642
rect 3378 585 3409 642
rect -130 571 3409 585
rect -231 541 3409 571
rect -231 423 -91 541
rect -231 366 -187 423
rect -130 366 -91 423
rect -231 218 -91 366
rect -231 161 -187 218
rect -130 161 -91 218
rect -231 13 -91 161
rect -231 -44 -187 13
rect -130 -44 -91 13
rect -231 -192 -91 -44
rect -231 -249 -187 -192
rect -130 -249 -91 -192
rect -231 -397 -91 -249
rect -231 -454 -187 -397
rect -130 -454 -91 -397
rect -231 -602 -91 -454
rect -231 -659 -187 -602
rect -130 -659 -91 -602
rect -231 -807 -91 -659
rect -231 -864 -187 -807
rect -130 -864 -91 -807
rect -231 -1012 -91 -864
rect -231 -1069 -187 -1012
rect -130 -1069 -91 -1012
rect -231 -1199 -91 -1069
rect 10 413 3170 440
rect 10 368 245 413
rect 10 320 40 368
rect 88 365 245 368
rect 293 365 450 413
rect 498 365 655 413
rect 703 365 860 413
rect 908 365 1065 413
rect 1113 365 1270 413
rect 1318 365 1475 413
rect 1523 365 1680 413
rect 1728 365 1885 413
rect 1933 365 2090 413
rect 2138 365 2295 413
rect 2343 365 2500 413
rect 2548 365 2705 413
rect 2753 365 2910 413
rect 2958 368 3170 413
rect 2958 365 3090 368
rect 88 340 3090 365
rect 88 320 120 340
rect 10 168 120 320
rect 10 120 40 168
rect 88 120 120 168
rect 10 -32 120 120
rect 3060 320 3090 340
rect 3138 320 3170 368
rect 3060 168 3170 320
rect 3060 120 3090 168
rect 3138 120 3170 168
rect 10 -80 40 -32
rect 88 -80 120 -32
rect 277 100 353 108
rect 277 48 289 100
rect 341 48 353 100
rect 277 -4 353 48
rect 277 -56 289 -4
rect 341 -56 353 -4
rect 277 -67 353 -56
rect 709 100 785 108
rect 709 48 721 100
rect 773 48 785 100
rect 709 -4 785 48
rect 709 -56 721 -4
rect 773 -56 785 -4
rect 1141 100 1217 108
rect 1141 48 1153 100
rect 1205 48 1217 100
rect 1141 -4 1217 48
rect 1141 -56 1153 -4
rect 1205 -56 1217 -4
rect 10 -232 120 -80
rect 508 -178 554 -62
rect 709 -67 785 -56
rect 10 -280 40 -232
rect 88 -280 120 -232
rect 242 -194 554 -178
rect 242 -244 394 -194
rect 444 -195 554 -194
rect 940 -195 986 -56
rect 1141 -67 1217 -56
rect 1573 100 1649 108
rect 1573 48 1585 100
rect 1637 48 1649 100
rect 1573 -4 1649 48
rect 1573 -56 1585 -4
rect 1637 -56 1649 -4
rect 444 -241 986 -195
rect 444 -244 554 -241
rect 242 -259 554 -244
rect 10 -432 120 -280
rect 10 -480 40 -432
rect 88 -480 120 -432
rect 10 -632 120 -480
rect 10 -680 40 -632
rect 88 -680 120 -632
rect 277 -486 353 -478
rect 277 -538 289 -486
rect 341 -538 353 -486
rect 508 -508 554 -259
rect 709 -486 785 -478
rect 277 -590 353 -538
rect 277 -642 289 -590
rect 341 -642 353 -590
rect 277 -653 353 -642
rect 709 -538 721 -486
rect 773 -538 785 -486
rect 709 -590 785 -538
rect 709 -642 721 -590
rect 773 -642 785 -590
rect 709 -653 785 -642
rect 10 -832 120 -680
rect 940 -733 986 -241
rect 1032 -348 1111 -335
rect 1032 -398 1047 -348
rect 1097 -354 1111 -348
rect 1372 -354 1418 -59
rect 1573 -67 1649 -56
rect 2005 100 2081 108
rect 2005 48 2017 100
rect 2069 48 2081 100
rect 2005 -4 2081 48
rect 2005 -56 2017 -4
rect 2069 -56 2081 -4
rect 1804 -131 1850 -62
rect 2005 -67 2081 -56
rect 2437 100 2513 108
rect 2437 48 2449 100
rect 2501 48 2513 100
rect 2437 -4 2513 48
rect 2437 -56 2449 -4
rect 2501 -56 2513 -4
rect 2869 100 2945 108
rect 2869 48 2881 100
rect 2933 48 2945 100
rect 2869 -4 2945 48
rect 1790 -144 1864 -131
rect 1790 -194 1802 -144
rect 1852 -194 1864 -144
rect 1790 -206 1864 -194
rect 1804 -354 1850 -206
rect 2236 -220 2282 -58
rect 2437 -67 2513 -56
rect 2669 -220 2715 -55
rect 2869 -56 2881 -4
rect 2933 -56 2945 -4
rect 2869 -67 2945 -56
rect 3060 -32 3170 120
rect 3060 -80 3090 -32
rect 3138 -80 3170 -32
rect 3060 -220 3170 -80
rect 2236 -232 3170 -220
rect 2236 -266 3090 -232
rect 1097 -398 1850 -354
rect 1032 -400 1850 -398
rect 1032 -413 1111 -400
rect 1141 -486 1217 -478
rect 1372 -486 1418 -400
rect 1573 -486 1649 -478
rect 1141 -538 1153 -486
rect 1205 -538 1217 -486
rect 1141 -590 1217 -538
rect 1141 -642 1153 -590
rect 1205 -642 1217 -590
rect 1141 -653 1217 -642
rect 1573 -538 1585 -486
rect 1637 -538 1649 -486
rect 1573 -590 1649 -538
rect 1573 -642 1585 -590
rect 1637 -642 1649 -590
rect 1573 -653 1649 -642
rect 1423 -731 1607 -720
rect 1423 -733 1434 -731
rect 1484 -732 1545 -731
rect 940 -779 1434 -733
rect 1423 -784 1434 -779
rect 1486 -784 1538 -732
rect 1595 -781 1607 -731
rect 1590 -784 1607 -781
rect 1423 -792 1607 -784
rect 10 -880 40 -832
rect 88 -880 120 -832
rect 230 -806 463 -793
rect 1426 -796 1601 -792
rect 230 -856 387 -806
rect 437 -856 463 -806
rect 1804 -829 1850 -400
rect 2892 -280 3090 -266
rect 3138 -280 3170 -232
rect 2892 -298 3170 -280
rect 2892 -478 2938 -298
rect 3060 -432 3170 -298
rect 2005 -486 2081 -478
rect 2005 -538 2017 -486
rect 2069 -538 2081 -486
rect 2005 -590 2081 -538
rect 2005 -642 2017 -590
rect 2069 -642 2081 -590
rect 2437 -486 2513 -478
rect 2437 -538 2449 -486
rect 2501 -538 2513 -486
rect 2437 -590 2513 -538
rect 2005 -653 2081 -642
rect 2236 -718 2282 -620
rect 2437 -642 2449 -590
rect 2501 -642 2513 -590
rect 2437 -653 2513 -642
rect 2869 -486 2945 -478
rect 2869 -538 2881 -486
rect 2933 -538 2945 -486
rect 2869 -590 2945 -538
rect 2869 -642 2881 -590
rect 2933 -642 2945 -590
rect 2162 -723 2337 -718
rect 2161 -730 2341 -723
rect 2161 -782 2170 -730
rect 2222 -734 2274 -730
rect 2223 -782 2274 -734
rect 2326 -735 2341 -730
rect 2328 -736 2341 -735
rect 2668 -736 2714 -643
rect 2869 -653 2945 -642
rect 3060 -480 3090 -432
rect 3138 -480 3170 -432
rect 3060 -632 3170 -480
rect 2328 -782 2714 -736
rect 3060 -680 3090 -632
rect 3138 -680 3170 -632
rect 2161 -784 2173 -782
rect 2223 -784 2278 -782
rect 2161 -785 2278 -784
rect 2328 -785 2341 -782
rect 2161 -796 2341 -785
rect 230 -870 463 -856
rect 1742 -841 1917 -829
rect 10 -1010 120 -880
rect 1742 -893 1750 -841
rect 1802 -893 1854 -841
rect 1906 -893 1917 -841
rect 1742 -905 1917 -893
rect 3060 -832 3170 -680
rect 3060 -880 3090 -832
rect 3138 -880 3170 -832
rect 3060 -1010 3170 -880
rect 10 -1032 3170 -1010
rect 10 -1080 40 -1032
rect 88 -1080 245 -1032
rect 293 -1080 450 -1032
rect 498 -1080 655 -1032
rect 703 -1080 860 -1032
rect 908 -1080 1065 -1032
rect 1113 -1080 1270 -1032
rect 1318 -1080 1475 -1032
rect 1523 -1080 1680 -1032
rect 1728 -1080 1885 -1032
rect 1933 -1080 2090 -1032
rect 2138 -1080 2295 -1032
rect 2343 -1080 2500 -1032
rect 2548 -1080 2705 -1032
rect 2753 -1080 2910 -1032
rect 2958 -1080 3090 -1032
rect 3138 -1080 3170 -1032
rect 10 -1110 3170 -1080
rect 3269 423 3409 541
rect 3269 366 3313 423
rect 3370 366 3409 423
rect 3269 218 3409 366
rect 3269 161 3313 218
rect 3370 161 3409 218
rect 3269 13 3409 161
rect 3269 -44 3313 13
rect 3370 -44 3409 13
rect 3269 -192 3409 -44
rect 3269 -249 3313 -192
rect 3370 -249 3409 -192
rect 3269 -397 3409 -249
rect 3269 -454 3313 -397
rect 3370 -454 3409 -397
rect 3269 -602 3409 -454
rect 3269 -659 3313 -602
rect 3370 -659 3409 -602
rect 3269 -807 3409 -659
rect 3269 -864 3313 -807
rect 3370 -864 3409 -807
rect 3269 -1012 3409 -864
rect 3269 -1069 3313 -1012
rect 3370 -1069 3409 -1012
rect 3269 -1199 3409 -1069
rect -231 -1217 3409 -1199
rect -231 -1274 -187 -1217
rect -130 -1243 3313 -1217
rect -130 -1274 4 -1243
rect -231 -1300 4 -1274
rect 61 -1300 209 -1243
rect 266 -1300 414 -1243
rect 471 -1300 619 -1243
rect 676 -1300 824 -1243
rect 881 -1300 1029 -1243
rect 1086 -1300 1234 -1243
rect 1291 -1300 1439 -1243
rect 1496 -1300 1644 -1243
rect 1701 -1300 1849 -1243
rect 1906 -1300 2054 -1243
rect 2111 -1300 2259 -1243
rect 2316 -1300 2464 -1243
rect 2521 -1300 2669 -1243
rect 2726 -1300 2874 -1243
rect 2931 -1300 3079 -1243
rect 3136 -1274 3313 -1243
rect 3370 -1274 3409 -1217
rect 3136 -1300 3409 -1274
rect -231 -1339 3409 -1300
rect -231 -1422 -91 -1339
rect -231 -1479 -187 -1422
rect -130 -1479 -91 -1422
rect 3269 -1422 3409 -1339
rect -231 -1627 -91 -1479
rect 476 -1461 648 -1447
rect 476 -1511 586 -1461
rect 636 -1511 648 -1461
rect 2525 -1461 2678 -1446
rect 476 -1524 648 -1511
rect 1136 -1521 1613 -1475
rect 1136 -1591 1182 -1521
rect -231 -1684 -187 -1627
rect -130 -1684 -91 -1627
rect -231 -1832 -91 -1684
rect 687 -1600 763 -1592
rect 687 -1652 699 -1600
rect 751 -1652 763 -1600
rect 687 -1704 763 -1652
rect 687 -1756 699 -1704
rect 751 -1756 763 -1704
rect 687 -1767 763 -1756
rect 1120 -1599 1196 -1591
rect 1567 -1595 1613 -1521
rect 2525 -1511 2538 -1461
rect 2588 -1511 2678 -1461
rect 2525 -1523 2678 -1511
rect 3269 -1479 3313 -1422
rect 3370 -1479 3409 -1422
rect 1120 -1651 1132 -1599
rect 1184 -1651 1196 -1599
rect 1120 -1703 1196 -1651
rect 1120 -1755 1132 -1703
rect 1184 -1755 1196 -1703
rect 1120 -1766 1196 -1755
rect 1981 -1604 2057 -1596
rect 1981 -1656 1993 -1604
rect 2045 -1656 2057 -1604
rect 1981 -1708 2057 -1656
rect 1981 -1760 1993 -1708
rect 2045 -1760 2057 -1708
rect -231 -1889 -187 -1832
rect -130 -1835 -91 -1832
rect 1351 -1835 1397 -1770
rect -130 -1867 1397 -1835
rect 1783 -1867 1829 -1769
rect 1981 -1771 2057 -1760
rect 2417 -1603 2493 -1595
rect 2417 -1655 2429 -1603
rect 2481 -1655 2493 -1603
rect 2417 -1707 2493 -1655
rect 2417 -1759 2429 -1707
rect 2481 -1759 2493 -1707
rect 2215 -1867 2261 -1768
rect 2417 -1770 2493 -1759
rect 3269 -1627 3409 -1479
rect 3269 -1684 3313 -1627
rect 3370 -1684 3409 -1627
rect 2647 -1867 2693 -1771
rect -130 -1889 2693 -1867
rect -231 -1913 2693 -1889
rect 3269 -1832 3409 -1684
rect 3269 -1889 3313 -1832
rect 3370 -1889 3409 -1832
rect -231 -2037 -91 -1913
rect 578 -1999 658 -1986
rect -231 -2094 -187 -2037
rect -130 -2094 -91 -2037
rect -231 -2242 -91 -2094
rect 487 -2001 658 -1999
rect 487 -2051 593 -2001
rect 643 -2051 658 -2001
rect 487 -2067 658 -2051
rect 1289 -1997 1464 -1985
rect 1289 -2049 1297 -1997
rect 1349 -2049 1401 -1997
rect 1453 -2049 1464 -1997
rect 1289 -2061 1464 -2049
rect 1724 -1988 1899 -1976
rect 1724 -2040 1732 -1988
rect 1784 -2040 1836 -1988
rect 1888 -2040 1899 -1988
rect 1724 -2052 1899 -2040
rect 2524 -1999 2601 -1991
rect 2524 -2007 2694 -1999
rect 487 -2134 538 -2067
rect -231 -2299 -187 -2242
rect -130 -2299 -91 -2242
rect -231 -2447 -91 -2299
rect 472 -2142 548 -2134
rect 472 -2194 484 -2142
rect 536 -2194 548 -2142
rect 472 -2246 548 -2194
rect 472 -2298 484 -2246
rect 536 -2298 548 -2246
rect 472 -2309 548 -2298
rect 687 -2141 763 -2133
rect 687 -2193 699 -2141
rect 751 -2193 763 -2141
rect 687 -2245 763 -2193
rect 687 -2297 699 -2245
rect 751 -2297 763 -2245
rect 687 -2308 763 -2297
rect 1119 -2141 1195 -2133
rect 1119 -2193 1131 -2141
rect 1183 -2193 1195 -2141
rect 1119 -2245 1195 -2193
rect 1119 -2297 1131 -2245
rect 1183 -2297 1195 -2245
rect 919 -2395 965 -2299
rect 1119 -2308 1195 -2297
rect 1351 -2395 1397 -2061
rect 1554 -2140 1630 -2132
rect 1554 -2192 1566 -2140
rect 1618 -2192 1630 -2140
rect 1554 -2244 1630 -2192
rect 1554 -2296 1566 -2244
rect 1618 -2296 1630 -2244
rect 1554 -2307 1630 -2296
rect 919 -2441 1397 -2395
rect 1443 -2386 1595 -2371
rect 1443 -2436 1456 -2386
rect 1505 -2436 1595 -2386
rect -231 -2504 -187 -2447
rect -130 -2504 -91 -2447
rect 1443 -2452 1595 -2436
rect 1783 -2402 1829 -2052
rect 2524 -2057 2537 -2007
rect 2587 -2057 2694 -2007
rect 2524 -2072 2694 -2057
rect 1981 -2140 2057 -2132
rect 1981 -2192 1993 -2140
rect 2045 -2192 2057 -2140
rect 1981 -2244 2057 -2192
rect 1981 -2296 1993 -2244
rect 2045 -2296 2057 -2244
rect 2416 -2141 2492 -2133
rect 2646 -2134 2694 -2072
rect 3269 -2037 3409 -1889
rect 3269 -2094 3313 -2037
rect 3370 -2094 3409 -2037
rect 2416 -2193 2428 -2141
rect 2480 -2193 2492 -2141
rect 2416 -2245 2492 -2193
rect 1981 -2307 2057 -2296
rect 2215 -2402 2261 -2291
rect 2416 -2297 2428 -2245
rect 2480 -2297 2492 -2245
rect 2416 -2308 2492 -2297
rect 2632 -2142 2708 -2134
rect 2632 -2194 2644 -2142
rect 2696 -2194 2708 -2142
rect 2632 -2246 2708 -2194
rect 2632 -2298 2644 -2246
rect 2696 -2298 2708 -2246
rect 2632 -2309 2708 -2298
rect 3269 -2242 3409 -2094
rect 3269 -2299 3313 -2242
rect 3370 -2299 3409 -2242
rect 1783 -2448 2261 -2402
rect 2307 -2387 2459 -2373
rect 2307 -2437 2319 -2387
rect 2369 -2437 2459 -2387
rect 2307 -2451 2459 -2437
rect 3269 -2447 3409 -2299
rect -231 -2599 -91 -2504
rect 3269 -2504 3313 -2447
rect 3370 -2504 3409 -2447
rect 3269 -2599 3409 -2504
rect -231 -2643 3409 -2599
rect -231 -2700 -185 -2643
rect -128 -2700 4 -2643
rect 61 -2700 209 -2643
rect 266 -2700 414 -2643
rect 471 -2700 619 -2643
rect 676 -2700 824 -2643
rect 881 -2700 1029 -2643
rect 1086 -2700 1234 -2643
rect 1291 -2700 1439 -2643
rect 1496 -2700 1644 -2643
rect 1701 -2700 1849 -2643
rect 1906 -2700 2054 -2643
rect 2111 -2700 2259 -2643
rect 2316 -2700 2464 -2643
rect 2521 -2700 2669 -2643
rect 2726 -2700 2874 -2643
rect 2931 -2700 3079 -2643
rect 3136 -2700 3316 -2643
rect 3373 -2700 3409 -2643
rect -231 -2739 3409 -2700
<< via1 >>
rect 289 48 341 100
rect 289 -56 341 -4
rect 721 48 773 100
rect 721 -56 773 -4
rect 1153 48 1205 100
rect 1153 -56 1205 -4
rect 1585 48 1637 100
rect 1585 -56 1637 -4
rect 289 -538 341 -486
rect 289 -642 341 -590
rect 721 -538 773 -486
rect 721 -642 773 -590
rect 2017 48 2069 100
rect 2017 -56 2069 -4
rect 2449 48 2501 100
rect 2449 -56 2501 -4
rect 2881 48 2933 100
rect 2881 -56 2933 -4
rect 1153 -538 1205 -486
rect 1153 -642 1205 -590
rect 1585 -538 1637 -486
rect 1585 -642 1637 -590
rect 1434 -781 1484 -732
rect 1484 -781 1486 -732
rect 1434 -784 1486 -781
rect 1538 -781 1545 -732
rect 1545 -781 1590 -732
rect 1538 -784 1590 -781
rect 2017 -538 2069 -486
rect 2017 -642 2069 -590
rect 2449 -538 2501 -486
rect 2449 -642 2501 -590
rect 2881 -538 2933 -486
rect 2881 -642 2933 -590
rect 2170 -734 2222 -730
rect 2170 -782 2173 -734
rect 2173 -782 2222 -734
rect 2274 -735 2326 -730
rect 2274 -782 2278 -735
rect 2278 -782 2326 -735
rect 1750 -893 1802 -841
rect 1854 -893 1906 -841
rect 699 -1652 751 -1600
rect 699 -1756 751 -1704
rect 1132 -1651 1184 -1599
rect 1132 -1755 1184 -1703
rect 1993 -1656 2045 -1604
rect 1993 -1760 2045 -1708
rect 2429 -1655 2481 -1603
rect 2429 -1759 2481 -1707
rect 1297 -2049 1349 -1997
rect 1401 -2049 1453 -1997
rect 1732 -2040 1784 -1988
rect 1836 -2040 1888 -1988
rect 484 -2194 536 -2142
rect 484 -2298 536 -2246
rect 699 -2193 751 -2141
rect 699 -2297 751 -2245
rect 1131 -2193 1183 -2141
rect 1131 -2297 1183 -2245
rect 1566 -2192 1618 -2140
rect 1566 -2296 1618 -2244
rect 1993 -2192 2045 -2140
rect 1993 -2296 2045 -2244
rect 2428 -2193 2480 -2141
rect 2428 -2297 2480 -2245
rect 2644 -2194 2696 -2142
rect 2644 -2298 2696 -2246
<< metal2 >>
rect 277 100 353 108
rect 277 48 289 100
rect 341 51 353 100
rect 709 100 785 108
rect 709 51 721 100
rect 341 48 721 51
rect 773 51 785 100
rect 1141 100 1217 108
rect 1141 51 1153 100
rect 773 48 1153 51
rect 1205 51 1217 100
rect 1573 100 1649 108
rect 1573 51 1585 100
rect 1205 48 1585 51
rect 1637 51 1649 100
rect 2005 100 2081 108
rect 2005 51 2017 100
rect 1637 48 2017 51
rect 2069 51 2081 100
rect 2437 100 2513 108
rect 2437 51 2449 100
rect 2069 48 2449 51
rect 2501 51 2513 100
rect 2869 100 2945 108
rect 2869 51 2881 100
rect 2501 48 2881 51
rect 2933 48 2945 100
rect 277 -4 2945 48
rect 277 -56 289 -4
rect 341 -6 721 -4
rect 341 -56 353 -6
rect 277 -67 353 -56
rect 709 -56 721 -6
rect 773 -6 1153 -4
rect 773 -56 785 -6
rect 709 -67 785 -56
rect 1141 -56 1153 -6
rect 1205 -6 1585 -4
rect 1205 -56 1217 -6
rect 1141 -67 1217 -56
rect 1573 -56 1585 -6
rect 1637 -6 2017 -4
rect 1637 -56 1649 -6
rect 1573 -67 1649 -56
rect 2005 -56 2017 -6
rect 2069 -6 2449 -4
rect 2069 -56 2081 -6
rect 2005 -67 2081 -56
rect 2437 -56 2449 -6
rect 2501 -6 2881 -4
rect 2501 -56 2513 -6
rect 2437 -67 2513 -56
rect 2869 -56 2881 -6
rect 2933 -56 2945 -4
rect 2869 -67 2945 -56
rect 277 -486 353 -478
rect 277 -538 289 -486
rect 341 -535 353 -486
rect 709 -486 785 -478
rect 709 -535 721 -486
rect 341 -538 721 -535
rect 773 -535 785 -486
rect 1141 -486 1217 -478
rect 1141 -535 1153 -486
rect 773 -538 1153 -535
rect 1205 -535 1217 -486
rect 1573 -486 1649 -478
rect 1573 -535 1585 -486
rect 1205 -538 1585 -535
rect 1637 -535 1649 -486
rect 2005 -486 2081 -478
rect 2005 -535 2017 -486
rect 1637 -538 2017 -535
rect 2069 -535 2081 -486
rect 2437 -486 2513 -478
rect 2437 -535 2449 -486
rect 2069 -538 2449 -535
rect 2501 -535 2513 -486
rect 2869 -486 2945 -478
rect 2869 -535 2881 -486
rect 2501 -538 2881 -535
rect 2933 -538 2945 -486
rect 277 -590 2945 -538
rect 277 -642 289 -590
rect 341 -592 721 -590
rect 341 -642 353 -592
rect 277 -653 353 -642
rect 709 -642 721 -592
rect 773 -592 1153 -590
rect 773 -642 785 -592
rect 709 -653 785 -642
rect 1141 -642 1153 -592
rect 1205 -592 1585 -590
rect 1205 -642 1217 -592
rect 1141 -653 1217 -642
rect 1573 -642 1585 -592
rect 1637 -592 2017 -590
rect 1637 -642 1649 -592
rect 1573 -653 1649 -642
rect 2005 -642 2017 -592
rect 2069 -592 2449 -590
rect 2069 -642 2081 -592
rect 2005 -653 2081 -642
rect 2437 -642 2449 -592
rect 2501 -592 2881 -590
rect 2501 -642 2513 -592
rect 2437 -653 2513 -642
rect 2869 -642 2881 -592
rect 2933 -642 2945 -590
rect 2869 -653 2945 -642
rect 1388 -732 1601 -720
rect 1388 -784 1434 -732
rect 1486 -784 1538 -732
rect 1590 -784 1601 -732
rect 1388 -796 1601 -784
rect 2162 -723 2337 -718
rect 2162 -730 2494 -723
rect 2162 -782 2170 -730
rect 2222 -782 2274 -730
rect 2326 -782 2494 -730
rect 2162 -794 2494 -782
rect 687 -1600 763 -1592
rect 687 -1652 699 -1600
rect 751 -1642 763 -1600
rect 1120 -1599 1196 -1591
rect 1120 -1642 1132 -1599
rect 751 -1651 1132 -1642
rect 1184 -1651 1196 -1599
rect 751 -1652 1196 -1651
rect 687 -1703 1196 -1652
rect 687 -1704 1132 -1703
rect 687 -1756 699 -1704
rect 751 -1756 763 -1704
rect 687 -1767 763 -1756
rect 1120 -1755 1132 -1704
rect 1184 -1755 1196 -1703
rect 1120 -1766 1196 -1755
rect 690 -2133 761 -1767
rect 1388 -1985 1464 -796
rect 2291 -801 2494 -794
rect 1742 -841 1917 -829
rect 1742 -893 1750 -841
rect 1802 -893 1854 -841
rect 1906 -893 1917 -841
rect 1742 -905 1917 -893
rect 1823 -1976 1899 -905
rect 1981 -1604 2057 -1596
rect 1981 -1656 1993 -1604
rect 2045 -1649 2057 -1604
rect 2416 -1603 2494 -801
rect 2416 -1649 2429 -1603
rect 2045 -1655 2429 -1649
rect 2481 -1655 2494 -1603
rect 2045 -1656 2494 -1655
rect 1981 -1704 2494 -1656
rect 1981 -1707 2493 -1704
rect 1981 -1708 2429 -1707
rect 1981 -1760 1993 -1708
rect 2045 -1711 2429 -1708
rect 2045 -1760 2057 -1711
rect 1981 -1771 2057 -1760
rect 2417 -1759 2429 -1711
rect 2481 -1759 2493 -1707
rect 2417 -1770 2493 -1759
rect 1289 -1997 1464 -1985
rect 1289 -2049 1297 -1997
rect 1349 -2049 1401 -1997
rect 1453 -2049 1464 -1997
rect 1289 -2061 1464 -2049
rect 1724 -1988 1899 -1976
rect 1724 -2040 1732 -1988
rect 1784 -2040 1836 -1988
rect 1888 -2040 1899 -1988
rect 1724 -2052 1899 -2040
rect 472 -2142 548 -2134
rect 472 -2194 484 -2142
rect 536 -2192 548 -2142
rect 687 -2141 763 -2133
rect 687 -2192 699 -2141
rect 536 -2193 699 -2192
rect 751 -2192 763 -2141
rect 1119 -2141 1195 -2133
rect 1119 -2192 1131 -2141
rect 751 -2193 1131 -2192
rect 1183 -2192 1195 -2141
rect 1554 -2140 1630 -2132
rect 1554 -2192 1566 -2140
rect 1618 -2192 1630 -2140
rect 1981 -2140 2057 -2132
rect 1981 -2192 1993 -2140
rect 2045 -2192 2057 -2140
rect 2416 -2141 2492 -2133
rect 2416 -2192 2428 -2141
rect 1183 -2193 2428 -2192
rect 2480 -2192 2492 -2141
rect 2632 -2142 2708 -2134
rect 2632 -2192 2644 -2142
rect 2480 -2193 2644 -2192
rect 536 -2194 2644 -2193
rect 2696 -2194 2708 -2142
rect 472 -2244 2708 -2194
rect 472 -2245 1566 -2244
rect 472 -2246 699 -2245
rect 472 -2298 484 -2246
rect 536 -2254 699 -2246
rect 536 -2298 548 -2254
rect 472 -2309 548 -2298
rect 687 -2297 699 -2254
rect 751 -2254 1131 -2245
rect 751 -2297 763 -2254
rect 687 -2308 763 -2297
rect 1119 -2297 1131 -2254
rect 1183 -2254 1566 -2245
rect 1183 -2297 1195 -2254
rect 1119 -2308 1195 -2297
rect 1554 -2296 1566 -2254
rect 1618 -2254 1993 -2244
rect 1618 -2296 1630 -2254
rect 1554 -2307 1630 -2296
rect 1981 -2296 1993 -2254
rect 2045 -2245 2708 -2244
rect 2045 -2254 2428 -2245
rect 2045 -2296 2057 -2254
rect 1981 -2307 2057 -2296
rect 2416 -2297 2428 -2254
rect 2480 -2246 2708 -2245
rect 2480 -2254 2644 -2246
rect 2480 -2297 2492 -2254
rect 2416 -2308 2492 -2297
rect 2632 -2298 2644 -2254
rect 2696 -2298 2708 -2246
rect 2632 -2309 2708 -2298
use nmos_3p3_FSHHD6  nmos_3p3_FSHHD6_0
timestamp 1695121232
transform 1 0 1590 0 1 -1681
box -276 -168 276 168
use nmos_3p3_QNHHD6  nmos_3p3_QNHHD6_0
timestamp 1694167386
transform 1 0 618 0 1 -2221
box -168 -168 168 168
use nmos_3p3_QNHHD6  nmos_3p3_QNHHD6_1
timestamp 1694167386
transform 1 0 2562 0 1 -2221
box -168 -168 168 168
use nmos_3p3_VMHHD6  nmos_3p3_VMHHD6_0
timestamp 1694167386
transform 1 0 2238 0 1 -1681
box -492 -168 492 168
use nmos_3p3_VMHHD6  nmos_3p3_VMHHD6_1
timestamp 1694167386
transform 1 0 1158 0 1 -2221
box -492 -168 492 168
use nmos_3p3_VMHHD6  nmos_3p3_VMHHD6_2
timestamp 1694167386
transform 1 0 2022 0 1 -2221
box -492 -168 492 168
use pmos_3p3_ZB3RD7  pmos_3p3_ZB3RD7_0
timestamp 1694080061
transform 1 0 2475 0 1 -568
box -554 -230 554 230
use pmos_3p3_ZB3RD7  pmos_3p3_ZB3RD7_1
timestamp 1694080061
transform 1 0 747 0 1 21
box -554 -230 554 230
use pmos_3p3_ZB3RD7  pmos_3p3_ZB3RD7_2
timestamp 1694080061
transform 1 0 1611 0 1 21
box -554 -230 554 230
use pmos_3p3_ZB3RD7  pmos_3p3_ZB3RD7_3
timestamp 1694080061
transform 1 0 2475 0 1 21
box -554 -230 554 230
use pmos_3p3_ZB3RD7  pmos_3p3_ZB3RD7_4
timestamp 1694080061
transform 1 0 747 0 1 -568
box -554 -230 554 230
use pmos_3p3_ZB3RD7  pmos_3p3_ZB3RD7_5
timestamp 1694080061
transform 1 0 1611 0 1 -568
box -554 -230 554 230
<< labels >>
flabel metal1 275 -223 275 -223 0 FreeSans 800 0 0 0 OUT
port 0 nsew
flabel metal1 272 -834 272 -834 0 FreeSans 800 0 0 0 OUTB
port 1 nsew
flabel metal1 502 -1481 502 -1481 0 FreeSans 800 0 0 0 EN
port 2 nsew
flabel metal1 2658 -1482 2658 -1482 0 FreeSans 800 0 0 0 VCONT
port 3 nsew
flabel metal1 2435 -2414 2435 -2414 0 FreeSans 800 0 0 0 INB
port 4 nsew
flabel metal1 1556 -2415 1556 -2415 0 FreeSans 800 0 0 0 IN
port 5 nsew
flabel metal1 103 -1868 103 -1868 0 FreeSans 800 0 0 0 VSS
port 6 nsew
flabel metal1 2947 -249 2947 -249 0 FreeSans 800 0 0 0 VDD
port 8 nsew
<< end >>
