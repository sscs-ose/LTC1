magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -2161 -5147 7956 2944
<< nwell >>
rect 0 788 5956 944
rect 403 757 3125 788
rect 3295 761 3575 788
rect 3707 760 4844 788
rect 5042 765 5257 788
rect 5524 762 5720 788
<< pwell >>
rect 2920 -2260 2970 -2254
rect 3327 -2260 3381 -2253
rect 3735 -2260 3791 -2252
rect 4144 -2260 4198 -2253
rect 4551 -2260 4605 -2254
rect 4959 -2260 5014 -2254
rect 5368 -2260 5429 -2254
<< psubdiff >>
rect 68 -3067 244 -3051
rect 68 -3113 136 -3067
rect 182 -3113 244 -3067
rect 68 -3130 244 -3113
rect 368 -3067 544 -3051
rect 368 -3113 436 -3067
rect 482 -3113 544 -3067
rect 368 -3130 544 -3113
rect 668 -3067 844 -3051
rect 668 -3113 736 -3067
rect 782 -3113 844 -3067
rect 668 -3130 844 -3113
rect 968 -3067 1144 -3051
rect 968 -3113 1036 -3067
rect 1082 -3113 1144 -3067
rect 968 -3130 1144 -3113
rect 1268 -3067 1444 -3051
rect 1268 -3113 1336 -3067
rect 1382 -3113 1444 -3067
rect 1268 -3130 1444 -3113
rect 1568 -3067 1744 -3051
rect 1568 -3113 1636 -3067
rect 1682 -3113 1744 -3067
rect 1568 -3130 1744 -3113
rect 1868 -3067 2044 -3051
rect 1868 -3113 1936 -3067
rect 1982 -3113 2044 -3067
rect 1868 -3130 2044 -3113
rect 2168 -3067 2344 -3051
rect 2168 -3113 2236 -3067
rect 2282 -3113 2344 -3067
rect 2168 -3130 2344 -3113
rect 2468 -3067 2644 -3051
rect 2468 -3113 2536 -3067
rect 2582 -3113 2644 -3067
rect 2468 -3130 2644 -3113
rect 2768 -3067 2944 -3051
rect 2768 -3113 2836 -3067
rect 2882 -3113 2944 -3067
rect 2768 -3130 2944 -3113
rect 3068 -3067 3244 -3051
rect 3068 -3113 3136 -3067
rect 3182 -3113 3244 -3067
rect 3068 -3130 3244 -3113
rect 3368 -3067 3544 -3051
rect 3368 -3113 3436 -3067
rect 3482 -3113 3544 -3067
rect 3368 -3130 3544 -3113
rect 3668 -3067 3844 -3051
rect 3668 -3113 3736 -3067
rect 3782 -3113 3844 -3067
rect 3668 -3130 3844 -3113
rect 3968 -3067 4144 -3051
rect 3968 -3113 4036 -3067
rect 4082 -3113 4144 -3067
rect 3968 -3130 4144 -3113
rect 4268 -3067 4444 -3051
rect 4268 -3113 4336 -3067
rect 4382 -3113 4444 -3067
rect 4268 -3130 4444 -3113
rect 4568 -3067 4744 -3051
rect 4568 -3113 4636 -3067
rect 4682 -3113 4744 -3067
rect 4568 -3130 4744 -3113
rect 4868 -3067 5044 -3051
rect 4868 -3113 4936 -3067
rect 4982 -3113 5044 -3067
rect 4868 -3130 5044 -3113
rect 5168 -3067 5344 -3051
rect 5168 -3113 5236 -3067
rect 5282 -3113 5344 -3067
rect 5168 -3130 5344 -3113
rect 5468 -3067 5644 -3051
rect 5468 -3113 5536 -3067
rect 5582 -3113 5644 -3067
rect 5468 -3130 5644 -3113
rect 5718 -3067 5894 -3051
rect 5718 -3113 5786 -3067
rect 5832 -3113 5894 -3067
rect 5718 -3130 5894 -3113
<< nsubdiff >>
rect 3315 905 3492 913
rect 3315 896 3493 905
rect 429 871 606 888
rect 429 825 496 871
rect 542 825 606 871
rect 429 809 606 825
rect 673 871 850 888
rect 673 825 740 871
rect 786 825 850 871
rect 673 809 850 825
rect 918 871 1095 888
rect 918 825 985 871
rect 1031 825 1095 871
rect 918 809 1095 825
rect 1162 871 1339 888
rect 1162 825 1229 871
rect 1275 825 1339 871
rect 1162 809 1339 825
rect 1407 871 1584 888
rect 1407 825 1474 871
rect 1520 825 1584 871
rect 1407 809 1584 825
rect 1652 871 1829 888
rect 1652 825 1719 871
rect 1765 825 1829 871
rect 1652 809 1829 825
rect 1896 871 2073 888
rect 1896 825 1963 871
rect 2009 825 2073 871
rect 1896 809 2073 825
rect 2141 871 2318 888
rect 2141 825 2208 871
rect 2254 825 2318 871
rect 2141 809 2318 825
rect 2386 871 2563 888
rect 2386 825 2453 871
rect 2499 825 2563 871
rect 2386 809 2563 825
rect 2630 871 2807 888
rect 2630 825 2697 871
rect 2743 825 2807 871
rect 2630 809 2807 825
rect 2883 881 3060 889
rect 2883 872 3061 881
rect 2883 826 2950 872
rect 2996 826 3061 872
rect 3315 850 3382 896
rect 3428 850 3493 896
rect 3315 839 3493 850
rect 3735 876 3912 884
rect 4157 876 4334 884
rect 4579 876 4756 884
rect 3735 867 3913 876
rect 3315 834 3492 839
rect 2883 815 3061 826
rect 3735 821 3802 867
rect 3848 821 3913 867
rect 2883 810 3060 815
rect 3735 810 3913 821
rect 4157 867 4335 876
rect 4157 821 4224 867
rect 4270 821 4335 867
rect 4157 810 4335 821
rect 4579 867 4757 876
rect 4579 821 4646 867
rect 4692 821 4757 867
rect 4579 810 4757 821
rect 5055 872 5232 880
rect 5055 863 5233 872
rect 5055 817 5122 863
rect 5168 817 5233 863
rect 3735 805 3912 810
rect 4157 805 4334 810
rect 4579 805 4756 810
rect 5055 806 5233 817
rect 5055 801 5232 806
<< psubdiffcont >>
rect 136 -3113 182 -3067
rect 436 -3113 482 -3067
rect 736 -3113 782 -3067
rect 1036 -3113 1082 -3067
rect 1336 -3113 1382 -3067
rect 1636 -3113 1682 -3067
rect 1936 -3113 1982 -3067
rect 2236 -3113 2282 -3067
rect 2536 -3113 2582 -3067
rect 2836 -3113 2882 -3067
rect 3136 -3113 3182 -3067
rect 3436 -3113 3482 -3067
rect 3736 -3113 3782 -3067
rect 4036 -3113 4082 -3067
rect 4336 -3113 4382 -3067
rect 4636 -3113 4682 -3067
rect 4936 -3113 4982 -3067
rect 5236 -3113 5282 -3067
rect 5536 -3113 5582 -3067
rect 5786 -3113 5832 -3067
<< nsubdiffcont >>
rect 496 825 542 871
rect 740 825 786 871
rect 985 825 1031 871
rect 1229 825 1275 871
rect 1474 825 1520 871
rect 1719 825 1765 871
rect 1963 825 2009 871
rect 2208 825 2254 871
rect 2453 825 2499 871
rect 2697 825 2743 871
rect 2950 826 2996 872
rect 3382 850 3428 896
rect 3802 821 3848 867
rect 4224 821 4270 867
rect 4646 821 4692 867
rect 5122 817 5168 863
<< polysilicon >>
rect 175 91 273 120
rect 786 91 878 121
rect 173 89 878 91
rect -158 53 878 89
rect -158 7 -134 53
rect -88 7 878 53
rect -158 -28 878 7
rect 988 58 4150 86
rect 988 12 1011 58
rect 1057 12 4150 58
rect -158 -29 185 -28
rect 988 -30 4150 12
rect 4254 64 5782 88
rect 4254 18 4277 64
rect 4323 18 5782 64
rect 4254 -29 5782 18
rect 5681 -99 5782 -29
rect 174 -728 477 -727
rect 174 -776 5781 -728
rect 2620 -1433 2722 -1404
rect 2620 -1479 2645 -1433
rect 2691 -1479 2722 -1433
rect -161 -1492 -66 -1482
rect -161 -1503 451 -1492
rect -161 -1549 -143 -1503
rect -97 -1549 451 -1503
rect -161 -1563 451 -1549
rect 548 -1501 645 -1487
rect 548 -1547 567 -1501
rect 613 -1511 645 -1501
rect 2620 -1505 2722 -1479
rect 2826 -1490 2926 -1424
rect 3438 -1490 3538 -1424
rect 4050 -1490 4150 -1424
rect 4662 -1490 4762 -1424
rect 5274 -1490 5374 -1424
rect 613 -1547 2076 -1511
rect 548 -1560 2076 -1547
rect 2792 -1560 5748 -1490
rect -161 -1568 -66 -1563
rect 2179 -2203 2279 -2200
rect 2179 -2260 2892 -2203
rect 138 -2895 646 -2887
rect 138 -2897 2279 -2895
rect 138 -2984 2891 -2897
rect 2276 -2985 2891 -2984
rect 2996 -2915 5748 -2890
rect 2996 -2961 3229 -2915
rect 3275 -2961 5748 -2915
rect 2996 -3001 5748 -2961
<< polycontact >>
rect -134 7 -88 53
rect 1011 12 1057 58
rect 4277 18 4323 64
rect 2645 -1479 2691 -1433
rect -143 -1549 -97 -1503
rect 567 -1547 613 -1501
rect 3229 -2961 3275 -2915
<< metal1 >>
rect 0 896 5956 944
rect 0 872 3382 896
rect 0 871 2950 872
rect 0 825 496 871
rect 542 825 740 871
rect 786 825 985 871
rect 1031 825 1229 871
rect 1275 825 1474 871
rect 1520 825 1719 871
rect 1765 825 1963 871
rect 2009 825 2208 871
rect 2254 825 2453 871
rect 2499 825 2697 871
rect 2743 826 2950 871
rect 2996 850 3382 872
rect 3428 867 5956 896
rect 3428 850 3802 867
rect 2996 826 3802 850
rect 2743 825 3802 826
rect 0 821 3802 825
rect 3848 821 4224 867
rect 4270 821 4646 867
rect 4692 863 5956 867
rect 4692 821 5122 863
rect 0 817 5122 821
rect 5168 817 5956 863
rect 0 753 5956 817
rect 99 677 145 753
rect 507 677 553 753
rect 914 675 961 753
rect 1323 677 1369 753
rect 1731 677 1777 753
rect 2139 677 2185 753
rect 2547 677 2593 753
rect 2955 677 3001 753
rect 3363 677 3409 753
rect 3771 676 3817 753
rect 4178 666 4226 753
rect 4587 675 4633 753
rect 4995 677 5041 753
rect 5403 678 5449 753
rect 5811 678 5857 753
rect 300 86 351 136
rect 709 86 758 147
rect -153 53 -76 78
rect 300 73 758 86
rect 1117 82 1166 166
rect 1526 82 1573 155
rect 1934 82 1981 156
rect 2343 82 2390 156
rect 2750 82 2797 154
rect 3158 82 3205 154
rect 3566 82 3613 154
rect 3974 82 4021 155
rect 1117 79 4021 82
rect 4383 80 4430 155
rect 4789 80 4836 155
rect 5198 80 5245 159
rect 5607 80 5654 155
rect 300 58 1070 73
rect 300 54 1011 58
rect -153 28 -134 53
rect -154 7 -134 28
rect -88 7 -76 53
rect -154 -16 -76 7
rect -24 12 1011 54
rect 1057 12 1070 58
rect -24 9 1070 12
rect -24 8 758 9
rect -154 -73 -80 -16
rect -154 -1503 -85 -73
rect -154 -1549 -143 -1503
rect -97 -1549 -85 -1503
rect -154 -1568 -85 -1549
rect -24 -1508 22 8
rect 987 -5 1070 9
rect 1117 64 4336 79
rect 1117 18 4277 64
rect 4323 18 4336 64
rect 1117 3 4336 18
rect 4383 7 5654 80
rect 5606 -164 5654 7
rect 5811 -136 5857 145
rect 68 -327 169 -304
rect 68 -379 94 -327
rect 146 -379 169 -327
rect 68 -401 169 -379
rect 474 -320 575 -294
rect 474 -372 499 -320
rect 551 -372 575 -320
rect 474 -392 575 -372
rect 879 -319 979 -289
rect 879 -371 904 -319
rect 956 -371 979 -319
rect 879 -390 979 -371
rect 1289 -306 1389 -277
rect 1289 -358 1314 -306
rect 1366 -358 1389 -306
rect 1289 -378 1389 -358
rect 1699 -302 1799 -274
rect 1699 -354 1722 -302
rect 1774 -354 1799 -302
rect 1699 -375 1799 -354
rect 2109 -293 2209 -265
rect 2109 -345 2132 -293
rect 2184 -345 2209 -293
rect 2109 -366 2209 -345
rect 2515 -292 2615 -265
rect 2515 -344 2543 -292
rect 2595 -344 2615 -292
rect 2515 -366 2615 -344
rect 2918 -283 3018 -255
rect 2918 -335 2945 -283
rect 2997 -335 3018 -283
rect 2918 -356 3018 -335
rect 3328 -280 3428 -249
rect 3328 -332 3355 -280
rect 3407 -332 3428 -280
rect 3328 -350 3428 -332
rect 3743 -278 3843 -250
rect 3743 -330 3766 -278
rect 3818 -330 3843 -278
rect 3743 -351 3843 -330
rect 4147 -280 4247 -251
rect 4147 -332 4171 -280
rect 4223 -332 4247 -280
rect 4147 -352 4247 -332
rect 4555 -280 4655 -255
rect 4555 -332 4581 -280
rect 4633 -332 4655 -280
rect 4555 -356 4655 -332
rect 4958 -280 5058 -251
rect 4958 -332 4982 -280
rect 5034 -332 5058 -280
rect 4958 -352 5058 -332
rect 5374 -276 5474 -247
rect 5374 -328 5398 -276
rect 5450 -328 5474 -276
rect 5374 -348 5474 -328
rect 5775 -261 5875 -236
rect 5775 -313 5799 -261
rect 5851 -313 5875 -261
rect 5775 -337 5875 -313
rect 302 -728 349 -658
rect 711 -728 757 -658
rect 1119 -728 1165 -651
rect 1526 -728 1572 -651
rect 1934 -728 1980 -651
rect 2342 -728 2388 -651
rect 2751 -728 2797 -653
rect 3158 -728 3204 -651
rect 3566 -728 3612 -652
rect 3975 -728 4021 -660
rect 4382 -728 4428 -662
rect 4791 -728 4837 -658
rect 5198 -728 5244 -657
rect 5606 -728 5653 -662
rect 302 -775 5653 -728
rect 302 -844 349 -775
rect 710 -836 757 -775
rect 1119 -836 1166 -775
rect 1527 -836 1574 -775
rect 1935 -835 1982 -775
rect 2343 -835 2390 -775
rect 2751 -835 2798 -775
rect 3159 -835 3206 -775
rect 3567 -835 3614 -775
rect 3975 -834 4022 -775
rect 4383 -834 4430 -775
rect 4792 -834 4839 -775
rect 5200 -834 5247 -775
rect 5606 -833 5653 -775
rect 5810 -838 5857 -667
rect 68 -1021 183 -988
rect 68 -1073 100 -1021
rect 152 -1073 183 -1021
rect 68 -1097 183 -1073
rect 471 -1015 586 -977
rect 471 -1067 499 -1015
rect 551 -1067 586 -1015
rect 471 -1086 586 -1067
rect 877 -1019 992 -981
rect 877 -1071 907 -1019
rect 959 -1071 992 -1019
rect 877 -1090 992 -1071
rect 1282 -1013 1397 -981
rect 1282 -1065 1312 -1013
rect 1364 -1065 1397 -1013
rect 1282 -1090 1397 -1065
rect 1692 -1030 1807 -995
rect 1692 -1082 1722 -1030
rect 1774 -1082 1807 -1030
rect 1692 -1104 1807 -1082
rect 2100 -1031 2215 -998
rect 2100 -1083 2130 -1031
rect 2182 -1083 2215 -1031
rect 2100 -1107 2215 -1083
rect 2504 -1042 2619 -1008
rect 2504 -1094 2538 -1042
rect 2590 -1094 2619 -1042
rect 2504 -1117 2619 -1094
rect 2918 -1052 3033 -1018
rect 2918 -1104 2950 -1052
rect 3002 -1104 3033 -1052
rect 2918 -1127 3033 -1104
rect 3330 -1038 3445 -1003
rect 3330 -1090 3361 -1038
rect 3413 -1090 3445 -1038
rect 3330 -1112 3445 -1090
rect 3737 -1036 3852 -1006
rect 3737 -1088 3768 -1036
rect 3820 -1088 3852 -1036
rect 3737 -1115 3852 -1088
rect 4139 -1033 4254 -999
rect 4139 -1085 4175 -1033
rect 4227 -1085 4254 -1033
rect 4139 -1108 4254 -1085
rect 4550 -1017 4665 -981
rect 4550 -1069 4580 -1017
rect 4632 -1069 4665 -1017
rect 4550 -1090 4665 -1069
rect 4966 -1005 5081 -972
rect 4966 -1057 4993 -1005
rect 5045 -1057 5081 -1005
rect 4966 -1081 5081 -1057
rect 5372 -999 5487 -964
rect 5372 -1051 5401 -999
rect 5453 -1051 5487 -999
rect 5372 -1073 5487 -1051
rect 5769 -991 5884 -959
rect 5769 -1043 5803 -991
rect 5855 -1043 5884 -991
rect 5769 -1068 5884 -1043
rect 2621 -1430 2718 -1415
rect 2621 -1482 2642 -1430
rect 2694 -1482 2718 -1430
rect 5607 -1438 5654 -1286
rect 258 -1501 628 -1487
rect 2621 -1495 2718 -1482
rect 258 -1508 567 -1501
rect -24 -1547 567 -1508
rect 613 -1547 628 -1501
rect -24 -1554 628 -1547
rect 269 -1617 315 -1554
rect 548 -1560 628 -1554
rect 5572 -1509 5955 -1438
rect 5572 -1615 5619 -1509
rect 654 -1822 743 -1810
rect 654 -1874 673 -1822
rect 725 -1874 743 -1822
rect 654 -1884 743 -1874
rect 1060 -1813 1149 -1798
rect 1060 -1865 1079 -1813
rect 1131 -1865 1149 -1813
rect 1470 -1801 1559 -1785
rect 1470 -1853 1490 -1801
rect 1542 -1853 1559 -1801
rect 1470 -1863 1559 -1853
rect 1875 -1793 1964 -1778
rect 1875 -1845 1894 -1793
rect 1946 -1845 1964 -1793
rect 1875 -1856 1964 -1845
rect 1060 -1876 1149 -1865
rect 2289 -2046 2379 -2029
rect 2289 -2098 2307 -2046
rect 2359 -2098 2379 -2046
rect 2289 -2114 2379 -2098
rect 2692 -2045 2782 -2029
rect 2692 -2097 2711 -2045
rect 2763 -2097 2782 -2045
rect 2692 -2111 2782 -2097
rect 3098 -2041 3192 -2025
rect 3098 -2093 3120 -2041
rect 3172 -2093 3192 -2041
rect 3098 -2105 3192 -2093
rect 3509 -2031 3596 -2016
rect 3509 -2083 3527 -2031
rect 3579 -2083 3596 -2031
rect 3509 -2095 3596 -2083
rect 3916 -2020 4006 -2005
rect 3916 -2072 3936 -2020
rect 3988 -2072 4006 -2020
rect 3916 -2085 4006 -2072
rect 4324 -2023 4415 -2006
rect 4324 -2075 4345 -2023
rect 4397 -2075 4415 -2023
rect 4324 -2089 4415 -2075
rect 4733 -2019 4826 -2005
rect 4733 -2071 4753 -2019
rect 4805 -2071 4826 -2019
rect 4733 -2085 4826 -2071
rect 5142 -2020 5231 -2005
rect 5142 -2072 5160 -2020
rect 5212 -2072 5231 -2020
rect 5142 -2085 5231 -2072
rect 5552 -2022 5640 -2008
rect 5552 -2074 5570 -2022
rect 5622 -2074 5640 -2022
rect 5552 -2086 5640 -2074
rect 64 -2208 111 -2149
rect 472 -2208 519 -2147
rect 881 -2208 928 -2149
rect 1289 -2208 1336 -2148
rect 1696 -2208 1743 -2148
rect 2104 -2208 2151 -2149
rect 2513 -2208 2560 -2147
rect 2920 -2208 2967 -2149
rect 3328 -2208 3375 -2149
rect 3737 -2208 3784 -2149
rect 4145 -2208 4192 -2149
rect 4553 -2208 4600 -2148
rect 4961 -2208 5008 -2148
rect 5369 -2208 5416 -2147
rect 5776 -2208 5823 -2149
rect 64 -2254 5823 -2208
rect 64 -2313 111 -2254
rect 472 -2313 519 -2254
rect 881 -2313 928 -2254
rect 1289 -2312 1336 -2254
rect 1696 -2312 1743 -2254
rect 2104 -2313 2151 -2254
rect 2513 -2311 2560 -2254
rect 2921 -2553 2997 -2254
rect 248 -2605 334 -2589
rect 248 -2657 266 -2605
rect 318 -2657 334 -2605
rect 248 -2671 334 -2657
rect 657 -2600 743 -2583
rect 657 -2652 674 -2600
rect 726 -2652 743 -2600
rect 657 -2666 743 -2652
rect 1063 -2598 1149 -2582
rect 1063 -2650 1081 -2598
rect 1133 -2650 1149 -2598
rect 1063 -2665 1149 -2650
rect 1473 -2598 1560 -2583
rect 1473 -2650 1491 -2598
rect 1543 -2650 1560 -2598
rect 1473 -2665 1560 -2650
rect 1882 -2598 1969 -2582
rect 1882 -2650 1899 -2598
rect 1951 -2650 1969 -2598
rect 1882 -2664 1969 -2650
rect 2287 -2597 2374 -2581
rect 2287 -2649 2304 -2597
rect 2356 -2649 2374 -2597
rect 2287 -2663 2374 -2649
rect 2695 -2596 2782 -2580
rect 2695 -2648 2712 -2596
rect 2764 -2648 2782 -2596
rect 2921 -2645 5822 -2553
rect 2695 -2662 2782 -2648
rect 65 -3024 111 -2858
rect 881 -3024 927 -2858
rect 1691 -3024 1751 -2832
rect 2503 -3024 2563 -2835
rect 3220 -2915 3282 -2645
rect 3220 -2961 3229 -2915
rect 3275 -2961 3282 -2915
rect 3220 -2973 3282 -2961
rect 3724 -3024 3784 -2833
rect 4954 -3024 5014 -2844
rect 0 -3067 5956 -3024
rect 0 -3113 136 -3067
rect 182 -3113 436 -3067
rect 482 -3113 736 -3067
rect 782 -3113 1036 -3067
rect 1082 -3113 1336 -3067
rect 1382 -3113 1636 -3067
rect 1682 -3113 1936 -3067
rect 1982 -3113 2236 -3067
rect 2282 -3113 2536 -3067
rect 2582 -3113 2836 -3067
rect 2882 -3113 3136 -3067
rect 3182 -3113 3436 -3067
rect 3482 -3113 3736 -3067
rect 3782 -3113 4036 -3067
rect 4082 -3113 4336 -3067
rect 4382 -3113 4636 -3067
rect 4682 -3113 4936 -3067
rect 4982 -3113 5236 -3067
rect 5282 -3113 5536 -3067
rect 5582 -3113 5786 -3067
rect 5832 -3113 5956 -3067
rect 0 -3147 5956 -3113
<< via1 >>
rect 94 -379 146 -327
rect 499 -372 551 -320
rect 904 -371 956 -319
rect 1314 -358 1366 -306
rect 1722 -354 1774 -302
rect 2132 -345 2184 -293
rect 2543 -344 2595 -292
rect 2945 -335 2997 -283
rect 3355 -332 3407 -280
rect 3766 -330 3818 -278
rect 4171 -332 4223 -280
rect 4581 -332 4633 -280
rect 4982 -332 5034 -280
rect 5398 -328 5450 -276
rect 5799 -313 5851 -261
rect 100 -1073 152 -1021
rect 499 -1067 551 -1015
rect 907 -1071 959 -1019
rect 1312 -1065 1364 -1013
rect 1722 -1082 1774 -1030
rect 2130 -1083 2182 -1031
rect 2538 -1094 2590 -1042
rect 2950 -1104 3002 -1052
rect 3361 -1090 3413 -1038
rect 3768 -1088 3820 -1036
rect 4175 -1085 4227 -1033
rect 4580 -1069 4632 -1017
rect 4993 -1057 5045 -1005
rect 5401 -1051 5453 -999
rect 5803 -1043 5855 -991
rect 2642 -1433 2694 -1430
rect 2642 -1479 2645 -1433
rect 2645 -1479 2691 -1433
rect 2691 -1479 2694 -1433
rect 2642 -1482 2694 -1479
rect 673 -1874 725 -1822
rect 1079 -1865 1131 -1813
rect 1490 -1853 1542 -1801
rect 1894 -1845 1946 -1793
rect 2307 -2098 2359 -2046
rect 2711 -2097 2763 -2045
rect 3120 -2093 3172 -2041
rect 3527 -2083 3579 -2031
rect 3936 -2072 3988 -2020
rect 4345 -2075 4397 -2023
rect 4753 -2071 4805 -2019
rect 5160 -2072 5212 -2020
rect 5570 -2074 5622 -2022
rect 266 -2657 318 -2605
rect 674 -2652 726 -2600
rect 1081 -2650 1133 -2598
rect 1491 -2650 1543 -2598
rect 1899 -2650 1951 -2598
rect 2304 -2649 2356 -2597
rect 2712 -2648 2764 -2596
<< metal2 >>
rect 66 -261 5875 -234
rect 66 -276 5799 -261
rect 66 -278 5398 -276
rect 66 -280 3766 -278
rect 66 -283 3355 -280
rect 66 -292 2945 -283
rect 66 -293 2543 -292
rect 66 -302 2132 -293
rect 66 -306 1722 -302
rect 66 -319 1314 -306
rect 66 -320 904 -319
rect 66 -327 499 -320
rect 66 -379 94 -327
rect 146 -372 499 -327
rect 551 -371 904 -320
rect 956 -358 1314 -319
rect 1366 -354 1722 -306
rect 1774 -345 2132 -302
rect 2184 -344 2543 -293
rect 2595 -335 2945 -292
rect 2997 -332 3355 -283
rect 3407 -330 3766 -280
rect 3818 -280 5398 -278
rect 3818 -330 4171 -280
rect 3407 -332 4171 -330
rect 4223 -332 4581 -280
rect 4633 -332 4982 -280
rect 5034 -328 5398 -280
rect 5450 -313 5799 -276
rect 5851 -313 5875 -261
rect 5450 -328 5875 -313
rect 5034 -332 5875 -328
rect 2997 -335 5875 -332
rect 2595 -344 5875 -335
rect 2184 -345 5875 -344
rect 1774 -354 5875 -345
rect 1366 -358 5875 -354
rect 956 -371 5875 -358
rect 551 -372 5875 -371
rect 146 -379 5875 -372
rect 66 -400 5875 -379
rect 68 -401 169 -400
rect 61 -991 5885 -949
rect 61 -999 5803 -991
rect 61 -1005 5401 -999
rect 61 -1013 4993 -1005
rect 61 -1015 1312 -1013
rect 61 -1021 499 -1015
rect 61 -1073 100 -1021
rect 152 -1067 499 -1021
rect 551 -1019 1312 -1015
rect 551 -1067 907 -1019
rect 152 -1071 907 -1067
rect 959 -1065 1312 -1019
rect 1364 -1017 4993 -1013
rect 1364 -1030 4580 -1017
rect 1364 -1065 1722 -1030
rect 959 -1071 1722 -1065
rect 152 -1073 1722 -1071
rect 61 -1082 1722 -1073
rect 1774 -1031 4580 -1030
rect 1774 -1082 2130 -1031
rect 61 -1083 2130 -1082
rect 2182 -1033 4580 -1031
rect 2182 -1036 4175 -1033
rect 2182 -1038 3768 -1036
rect 2182 -1042 3361 -1038
rect 2182 -1083 2538 -1042
rect 61 -1094 2538 -1083
rect 2590 -1052 3361 -1042
rect 2590 -1094 2950 -1052
rect 61 -1104 2950 -1094
rect 3002 -1090 3361 -1052
rect 3413 -1088 3768 -1038
rect 3820 -1085 4175 -1036
rect 4227 -1069 4580 -1033
rect 4632 -1057 4993 -1017
rect 5045 -1051 5401 -1005
rect 5453 -1043 5803 -999
rect 5855 -1043 5885 -991
rect 5453 -1051 5885 -1043
rect 5045 -1057 5885 -1051
rect 4632 -1069 5885 -1057
rect 4227 -1085 5885 -1069
rect 3820 -1088 5885 -1085
rect 3413 -1090 5885 -1088
rect 3002 -1104 5885 -1090
rect 61 -1108 5885 -1104
rect 2504 -1117 2619 -1108
rect 2918 -1127 3033 -1108
rect 3330 -1112 3445 -1108
rect 3737 -1115 3852 -1108
rect 2619 -1430 2718 -1413
rect 2619 -1482 2642 -1430
rect 2694 -1482 2718 -1430
rect 2619 -1773 2718 -1482
rect 1883 -1775 2718 -1773
rect 653 -1793 2718 -1775
rect 653 -1801 1894 -1793
rect 653 -1813 1490 -1801
rect 653 -1822 1079 -1813
rect 653 -1874 673 -1822
rect 725 -1865 1079 -1822
rect 1131 -1853 1490 -1813
rect 1542 -1845 1894 -1801
rect 1946 -1845 2718 -1793
rect 1542 -1853 2718 -1845
rect 1131 -1865 2718 -1853
rect 725 -1874 2718 -1865
rect 653 -1884 2718 -1874
rect 2289 -2019 5640 -2003
rect 2289 -2020 4753 -2019
rect 2289 -2031 3936 -2020
rect 2289 -2041 3527 -2031
rect 2289 -2045 3120 -2041
rect 2289 -2046 2711 -2045
rect 2289 -2098 2307 -2046
rect 2359 -2097 2711 -2046
rect 2763 -2093 3120 -2045
rect 3172 -2083 3527 -2041
rect 3579 -2072 3936 -2031
rect 3988 -2023 4753 -2020
rect 3988 -2072 4345 -2023
rect 3579 -2075 4345 -2072
rect 4397 -2071 4753 -2023
rect 4805 -2020 5640 -2019
rect 4805 -2071 5160 -2020
rect 4397 -2072 5160 -2071
rect 5212 -2022 5640 -2020
rect 5212 -2072 5570 -2022
rect 4397 -2074 5570 -2072
rect 5622 -2074 5640 -2022
rect 4397 -2075 5640 -2074
rect 3579 -2083 5640 -2075
rect 3172 -2093 5640 -2083
rect 2763 -2097 5640 -2093
rect 2359 -2098 5640 -2097
rect 2289 -2114 5640 -2098
rect 2398 -2579 2480 -2114
rect 248 -2596 2791 -2579
rect 248 -2597 2712 -2596
rect 248 -2598 2304 -2597
rect 248 -2600 1081 -2598
rect 248 -2605 674 -2600
rect 248 -2657 266 -2605
rect 318 -2652 674 -2605
rect 726 -2650 1081 -2600
rect 1133 -2650 1491 -2598
rect 1543 -2650 1899 -2598
rect 1951 -2649 2304 -2598
rect 2356 -2648 2712 -2597
rect 2764 -2648 2791 -2596
rect 2356 -2649 2791 -2648
rect 1951 -2650 2791 -2649
rect 726 -2652 2791 -2650
rect 318 -2657 2791 -2652
rect 248 -2671 2791 -2657
use nmos_3p3_7NPLVN  nmos_3p3_7NPLVN_0
timestamp 1713185578
transform 1 0 2944 0 1 -2580
box -2916 -348 2916 348
use nmos_3p3_8FEAMQ  nmos_3p3_8FEAMQ_0
timestamp 1713185578
transform 1 0 292 0 1 -1884
box -264 -348 264 348
use nmos_3p3_JEEAMQ  nmos_3p3_JEEAMQ_0
timestamp 1713185578
transform 1 0 1312 0 1 -1884
box -876 -348 876 348
use nmos_3p3_PLQLVN  nmos_3p3_PLQLVN_0
timestamp 1713185578
transform 1 0 3964 0 1 -1884
box -1896 -348 1896 348
use pmos_3p3_MDMPD7  pmos_3p3_MDMPD7_0
timestamp 1713185578
transform 1 0 2978 0 1 -752
box -2978 -758 2978 758
use pmos_3p3_MV44E7  pmos_3p3_MV44E7_0
timestamp 1713185578
transform 1 0 2570 0 1 410
box -1754 -410 1754 410
use pmos_3p3_PPYSL5  pmos_3p3_PPYSL5_0
timestamp 1713185578
transform 1 0 530 0 1 410
box -530 -410 530 410
use pmos_3p3_PPZSL5  pmos_3p3_PPZSL5_0
timestamp 1713185578
transform 1 0 5018 0 1 410
box -938 -410 938 410
<< labels >>
flabel nsubdiffcont 3403 873 3403 873 0 FreeSans 750 0 0 0 VDD
flabel psubdiffcont 2859 -3090 2859 -3090 0 FreeSans 750 0 0 0 VSS
flabel metal1 s -131 -741 -131 -741 0 FreeSans 750 0 0 0 IN
port 1 nsew
flabel metal1 s 5909 -1469 5909 -1469 0 FreeSans 750 0 0 0 OUT
port 2 nsew
<< end >>
