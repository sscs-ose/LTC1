magic
tech gf180mcuC
magscale 1 10
timestamp 1714137641
<< nwell >>
rect -64 682 500 863
<< psubdiff >>
rect 13 -105 402 -91
rect 13 -151 75 -105
rect 333 -151 402 -105
rect 13 -167 402 -151
<< nsubdiff >>
rect 41 814 395 828
rect 41 768 85 814
rect 312 768 395 814
rect 41 755 395 768
<< psubdiffcont >>
rect 75 -151 333 -105
<< nsubdiffcont >>
rect 85 768 312 814
<< polysilicon >>
rect 311 421 391 427
rect 112 334 166 421
rect 63 318 166 334
rect 63 268 81 318
rect 130 268 166 318
rect 63 254 166 268
rect 112 200 166 254
rect 272 414 391 421
rect 272 366 326 414
rect 374 366 391 414
rect 272 360 391 366
rect 272 350 390 360
rect 272 200 327 350
<< polycontact >>
rect 81 268 130 318
rect 326 366 374 414
<< metal1 >>
rect -64 817 500 863
rect -64 814 499 817
rect -64 768 85 814
rect 312 768 499 814
rect -64 708 499 768
rect 32 471 89 708
rect 186 470 253 545
rect 354 473 411 708
rect 63 325 144 334
rect 10 318 144 325
rect 10 278 81 318
rect 63 268 81 278
rect 130 268 144 318
rect 63 254 144 268
rect 191 314 243 470
rect 311 414 465 418
rect 311 366 326 414
rect 374 366 465 414
rect 311 361 465 366
rect 311 360 391 361
rect 191 265 521 314
rect 351 259 521 265
rect 34 -79 88 149
rect 186 70 255 156
rect 351 80 406 259
rect -70 -105 493 -79
rect -70 -151 75 -105
rect 333 -151 493 -105
rect -70 -188 493 -151
use nmos_3p3_5QNVWA  nmos_3p3_5QNVWA_0
timestamp 1714126980
transform 1 0 140 0 1 112
box -140 -112 140 112
use nmos_3p3_5QNVWA  nmos_3p3_5QNVWA_1
timestamp 1714126980
transform 1 0 300 0 1 112
box -140 -112 140 112
use pmos_3p3_M8SWPS  pmos_3p3_M8SWPS_0
timestamp 1714137641
transform 1 0 300 0 1 545
box -202 -210 202 210
use pmos_3p3_M8SWPS  pmos_3p3_M8SWPS_1
timestamp 1714137641
transform 1 0 140 0 1 545
box -202 -210 202 210
<< labels >>
flabel metal1 25 300 25 300 0 FreeSans 320 0 0 0 IN2
port 0 nsew
flabel metal1 495 289 495 289 0 FreeSans 320 0 0 0 OUT
port 1 nsew
flabel metal1 445 398 445 398 0 FreeSans 320 0 0 0 IN1
port 2 nsew
flabel psubdiffcont 210 -130 210 -130 0 FreeSans 320 0 0 0 VSS
port 4 nsew
flabel nsubdiffcont 196 796 196 796 0 FreeSans 480 0 0 0 VDD
port 3 nsew
<< end >>
